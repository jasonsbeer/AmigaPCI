-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 25 2025 18:07:05

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_350_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_376_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_280_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_288_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_325_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_308_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_350_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_355_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_389_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\ : std_logic;
signal \U712_CHIP_RAM.N_348_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \DBRn_c_i_cascade_\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \LATCH_CLK_0_i\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_350\ : std_logic;
signal \U712_CHIP_RAM.N_283\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_403\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_280\ : std_logic;
signal \U712_CHIP_RAM.N_301_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_280_2\ : std_logic;
signal \U712_CHIP_RAM.N_192\ : std_logic;
signal \U712_CHIP_RAM.N_192_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_215\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_345\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_100\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_400_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_266\ : std_logic;
signal \U712_CHIP_RAM.N_304_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_249\ : std_logic;
signal \U712_CHIP_RAM.N_355\ : std_logic;
signal \U712_CHIP_RAM.N_350_0\ : std_logic;
signal \U712_CHIP_RAM.N_291_cascade_\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \N_246\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \LATCH_REG\ : std_logic;
signal \REG_CPU_CYCLE\ : std_logic;
signal \INVU712_REG_SM.REGENnC_net\ : std_logic;
signal \ASn_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \INVU712_REG_SM.ASnC_net\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_399\ : std_logic;
signal \U712_CHIP_RAM.N_399_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_277\ : std_logic;
signal \U712_CHIP_RAM.N_277_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_347_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_353\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_347\ : std_logic;
signal \U712_CHIP_RAM.N_343_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_391\ : std_logic;
signal \U712_CHIP_RAM.N_391_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_387\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\ : std_logic;
signal \U712_CHIP_RAM.N_352\ : std_logic;
signal \U712_CHIP_RAM.N_343\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_234\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0\ : std_logic;
signal \WRITE_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_292\ : std_logic;
signal \U712_CHIP_RAM.N_19\ : std_logic;
signal \U712_BYTE_ENABLE.N_185_i\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_5\ : std_logic;
signal \INVU712_REG_SM.CYCLE_RUNC_net\ : std_logic;
signal \U712_REG_SM.N_229_cascade_\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_0C_net\ : std_logic;
signal \U712_REG_SM.LATCH_REG_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_4\ : std_logic;
signal \U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CPU_CYCLE_e_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_224\ : std_logic;
signal \U712_REG_SM.N_224_cascade_\ : std_logic;
signal \U712_REG_SM.N_209_cascade_\ : std_logic;
signal \U712_REG_SM.LDSn_7_iv_i_0\ : std_logic;
signal \U712_REG_SM.N_297_cascade_\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_295_cascade_\ : std_logic;
signal \U712_REG_SM.N_153\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \INVU712_REG_SM.C3_SYNC_1C_net\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.CYCLE_RUNZ0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \INVU712_REG_SM.C1_SYNC_0C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_136\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_405\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_405_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_303_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_348\ : std_logic;
signal \U712_CHIP_RAM.N_186\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.N_198\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.N_313_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \LATCH_RAM\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_319_cascade_\ : std_logic;
signal \N_58_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_320\ : std_logic;
signal \N_56_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_318\ : std_logic;
signal \U712_BYTE_ENABLE.N_323_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\ : std_logic;
signal \N_54_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLE\ : std_logic;
signal \U712_BYTE_ENABLE.N_315_cascade_\ : std_logic;
signal \N_60_i\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_3\ : std_logic;
signal \REG_WRITE_CYCLE\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_REG_SM.UDSn_7_iv_i_0\ : std_logic;
signal \U712_REG_SM.N_245\ : std_logic;
signal \U712_REG_SM.un15_0_i_0_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_6\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_7\ : std_logic;
signal \U712_REG_SM.N_209\ : std_logic;
signal \U712_REG_SM.N_229\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_1\ : std_logic;
signal \INVU712_REG_SM.REG_TACKC_net\ : std_logic;
signal \N_858_i\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_2\ : std_logic;
signal \U712_REG_SM.REG_TACK_0_sqmuxa\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_1\ : std_logic;
signal \INVU712_REG_SM.DBR_SYNC_0C_net\ : std_logic;
signal \REG_CYCLE\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \N_118_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_BYTE_ENABLE_UUBE_i\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \N_386\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \RASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \CLK40_PLL_g\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.N_8\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \CPU_TACK\ : std_logic;
signal \U712_CYCLE_TERM.N_227_i_0_0_cascade_\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.N_227_i_0_en_cascade_\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CYCLE_TERM.N_227_i_0_en_0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CPU_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4051\,
            RESETB => \N__8704\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11804\,
            DIN => \N__11803\,
            DOUT => \N__11802\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11804\,
            PADOUT => \N__11803\,
            PADIN => \N__11802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11795\,
            DIN => \N__11794\,
            DOUT => \N__11793\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11795\,
            PADOUT => \N__11794\,
            PADIN => \N__11793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11786\,
            DIN => \N__11785\,
            DOUT => \N__11784\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11786\,
            PADOUT => \N__11785\,
            PADIN => \N__11784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9604\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11777\,
            DIN => \N__11776\,
            DOUT => \N__11775\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11777\,
            PADOUT => \N__11776\,
            PADIN => \N__11775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11768\,
            DIN => \N__11767\,
            DOUT => \N__11766\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11768\,
            PADOUT => \N__11767\,
            PADIN => \N__11766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11759\,
            DIN => \N__11758\,
            DOUT => \N__11757\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11759\,
            PADOUT => \N__11758\,
            PADIN => \N__11757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11750\,
            DIN => \N__11749\,
            DOUT => \N__11748\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11750\,
            PADOUT => \N__11749\,
            PADIN => \N__11748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11741\,
            DIN => \N__11740\,
            DOUT => \N__11739\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11741\,
            PADOUT => \N__11740\,
            PADIN => \N__11739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11732\,
            DIN => \N__11731\,
            DOUT => \N__11730\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11732\,
            PADOUT => \N__11731\,
            PADIN => \N__11730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11723\,
            DIN => \N__11722\,
            DOUT => \N__11721\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11723\,
            PADOUT => \N__11722\,
            PADIN => \N__11721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11714\,
            DIN => \N__11713\,
            DOUT => \N__11712\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11714\,
            PADOUT => \N__11713\,
            PADIN => \N__11712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11705\,
            DIN => \N__11704\,
            DOUT => \N__11703\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11705\,
            PADOUT => \N__11704\,
            PADIN => \N__11703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11696\,
            DIN => \N__11695\,
            DOUT => \N__11694\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11696\,
            PADOUT => \N__11695\,
            PADIN => \N__11694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11687\,
            DIN => \N__11686\,
            DOUT => \N__11685\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11687\,
            PADOUT => \N__11686\,
            PADIN => \N__11685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11678\,
            DIN => \N__11677\,
            DOUT => \N__11676\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11678\,
            PADOUT => \N__11677\,
            PADIN => \N__11676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11669\,
            DIN => \N__11668\,
            DOUT => \N__11667\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11669\,
            PADOUT => \N__11668\,
            PADIN => \N__11667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4345\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11660\,
            DIN => \N__11659\,
            DOUT => \N__11658\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11660\,
            PADOUT => \N__11659\,
            PADIN => \N__11658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11651\,
            DIN => \N__11650\,
            DOUT => \N__11649\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11651\,
            PADOUT => \N__11650\,
            PADIN => \N__11649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11642\,
            DIN => \N__11641\,
            DOUT => \N__11640\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11642\,
            PADOUT => \N__11641\,
            PADIN => \N__11640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11633\,
            DIN => \N__11632\,
            DOUT => \N__11631\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11633\,
            PADOUT => \N__11632\,
            PADIN => \N__11631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11624\,
            DIN => \N__11623\,
            DOUT => \N__11622\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11624\,
            PADOUT => \N__11623\,
            PADIN => \N__11622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11615\,
            DIN => \N__11614\,
            DOUT => \N__11613\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11615\,
            PADOUT => \N__11614\,
            PADIN => \N__11613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11606\,
            DIN => \N__11605\,
            DOUT => \N__11604\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11606\,
            PADOUT => \N__11605\,
            PADIN => \N__11604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7903\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11597\,
            DIN => \N__11596\,
            DOUT => \N__11595\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11597\,
            PADOUT => \N__11596\,
            PADIN => \N__11595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11588\,
            DIN => \N__11587\,
            DOUT => \N__11586\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11588\,
            PADOUT => \N__11587\,
            PADIN => \N__11586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11579\,
            DIN => \N__11578\,
            DOUT => \N__11577\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11579\,
            PADOUT => \N__11578\,
            PADIN => \N__11577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11570\,
            DIN => \N__11569\,
            DOUT => \N__11568\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11570\,
            PADOUT => \N__11569\,
            PADIN => \N__11568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11561\,
            DIN => \N__11560\,
            DOUT => \N__11559\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11561\,
            PADOUT => \N__11560\,
            PADIN => \N__11559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11552\,
            DIN => \N__11551\,
            DOUT => \N__11550\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11552\,
            PADOUT => \N__11551\,
            PADIN => \N__11550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11543\,
            DIN => \N__11542\,
            DOUT => \N__11541\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11543\,
            PADOUT => \N__11542\,
            PADIN => \N__11541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11534\,
            DIN => \N__11533\,
            DOUT => \N__11532\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11534\,
            PADOUT => \N__11533\,
            PADIN => \N__11532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11525\,
            DIN => \N__11524\,
            DOUT => \N__11523\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11525\,
            PADOUT => \N__11524\,
            PADIN => \N__11523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11516\,
            DIN => \N__11515\,
            DOUT => \N__11514\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11516\,
            PADOUT => \N__11515\,
            PADIN => \N__11514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11507\,
            DIN => \N__11506\,
            DOUT => \N__11505\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11507\,
            PADOUT => \N__11506\,
            PADIN => \N__11505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11498\,
            DIN => \N__11497\,
            DOUT => \N__11496\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11498\,
            PADOUT => \N__11497\,
            PADIN => \N__11496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8332\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11489\,
            DIN => \N__11488\,
            DOUT => \N__11487\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11489\,
            PADOUT => \N__11488\,
            PADIN => \N__11487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6391\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11480\,
            DIN => \N__11479\,
            DOUT => \N__11478\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11480\,
            PADOUT => \N__11479\,
            PADIN => \N__11478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4389\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11471\,
            DIN => \N__11470\,
            DOUT => \N__11469\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11471\,
            PADOUT => \N__11470\,
            PADIN => \N__11469\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4183\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11462\,
            DIN => \N__11461\,
            DOUT => \N__11460\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11462\,
            PADOUT => \N__11461\,
            PADIN => \N__11460\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11453\,
            DIN => \N__11452\,
            DOUT => \N__11451\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11453\,
            PADOUT => \N__11452\,
            PADIN => \N__11451\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4711\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11444\,
            DIN => \N__11443\,
            DOUT => \N__11442\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11444\,
            PADOUT => \N__11443\,
            PADIN => \N__11442\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11435\,
            DIN => \N__11434\,
            DOUT => \N__11433\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11435\,
            PADOUT => \N__11434\,
            PADIN => \N__11433\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11426\,
            DIN => \N__11425\,
            DOUT => \N__11424\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11426\,
            PADOUT => \N__11425\,
            PADIN => \N__11424\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11417\,
            DIN => \N__11416\,
            DOUT => \N__11415\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11417\,
            PADOUT => \N__11416\,
            PADIN => \N__11415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11408\,
            DIN => \N__11407\,
            DOUT => \N__11406\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11408\,
            PADOUT => \N__11407\,
            PADIN => \N__11406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11399\,
            DIN => \N__11398\,
            DOUT => \N__11397\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11399\,
            PADOUT => \N__11398\,
            PADIN => \N__11397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8725\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11390\,
            DIN => \N__11389\,
            DOUT => \N__11388\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11390\,
            PADOUT => \N__11389\,
            PADIN => \N__11388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11381\,
            DIN => \N__11380\,
            DOUT => \N__11379\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11381\,
            PADOUT => \N__11380\,
            PADIN => \N__11379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4382\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11372\,
            DIN => \N__11371\,
            DOUT => \N__11370\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11372\,
            PADOUT => \N__11371\,
            PADIN => \N__11370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9538\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11363\,
            DIN => \N__11362\,
            DOUT => \N__11361\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11363\,
            PADOUT => \N__11362\,
            PADIN => \N__11361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11354\,
            DIN => \N__11353\,
            DOUT => \N__11352\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11354\,
            PADOUT => \N__11353\,
            PADIN => \N__11352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7078\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11345\,
            DIN => \N__11344\,
            DOUT => \N__11343\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11345\,
            PADOUT => \N__11344\,
            PADIN => \N__11343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8254\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11336\,
            DIN => \N__11335\,
            DOUT => \N__11334\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11336\,
            PADOUT => \N__11335\,
            PADIN => \N__11334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4765\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11327\,
            DIN => \N__11326\,
            DOUT => \N__11325\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11327\,
            PADOUT => \N__11326\,
            PADIN => \N__11325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11318\,
            DIN => \N__11317\,
            DOUT => \N__11316\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11318\,
            PADOUT => \N__11317\,
            PADIN => \N__11316\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11309\,
            DIN => \N__11308\,
            DOUT => \N__11307\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11309\,
            PADOUT => \N__11308\,
            PADIN => \N__11307\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7123\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11300\,
            DIN => \N__11299\,
            DOUT => \N__11298\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11300\,
            PADOUT => \N__11299\,
            PADIN => \N__11298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8314\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11291\,
            DIN => \N__11290\,
            DOUT => \N__11289\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11291\,
            PADOUT => \N__11290\,
            PADIN => \N__11289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11282\,
            DIN => \N__11281\,
            DOUT => \N__11280\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11282\,
            PADOUT => \N__11281\,
            PADIN => \N__11280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11273\,
            DIN => \N__11272\,
            DOUT => \N__11271\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11273\,
            PADOUT => \N__11272\,
            PADIN => \N__11271\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11264\,
            DIN => \N__11263\,
            DOUT => \N__11262\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11264\,
            PADOUT => \N__11263\,
            PADIN => \N__11262\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11255\,
            DIN => \N__11254\,
            DOUT => \N__11253\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11255\,
            PADOUT => \N__11254\,
            PADIN => \N__11253\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11246\,
            DIN => \N__11245\,
            DOUT => \N__11244\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11246\,
            PADOUT => \N__11245\,
            PADIN => \N__11244\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11237\,
            DIN => \N__11236\,
            DOUT => \N__11235\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11237\,
            PADOUT => \N__11236\,
            PADIN => \N__11235\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8179\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11228\,
            DIN => \N__11227\,
            DOUT => \N__11226\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11228\,
            PADOUT => \N__11227\,
            PADIN => \N__11226\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8005\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11219\,
            DIN => \N__11218\,
            DOUT => \N__11217\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11219\,
            PADOUT => \N__11218\,
            PADIN => \N__11217\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11210\,
            DIN => \N__11209\,
            DOUT => \N__11208\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11210\,
            PADOUT => \N__11209\,
            PADIN => \N__11208\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6937\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11201\,
            DIN => \N__11200\,
            DOUT => \N__11199\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11201\,
            PADOUT => \N__11200\,
            PADIN => \N__11199\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7318\,
            DIN0 => OPEN,
            DOUT0 => \N__8413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11192\,
            DIN => \N__11191\,
            DOUT => \N__11190\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11192\,
            PADOUT => \N__11191\,
            PADIN => \N__11190\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9475\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11183\,
            DIN => \N__11182\,
            DOUT => \N__11181\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11183\,
            PADOUT => \N__11182\,
            PADIN => \N__11181\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11174\,
            DIN => \N__11173\,
            DOUT => \N__11172\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11174\,
            PADOUT => \N__11173\,
            PADIN => \N__11172\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11165\,
            DIN => \N__11164\,
            DOUT => \N__11163\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11165\,
            PADOUT => \N__11164\,
            PADIN => \N__11163\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11156\,
            DIN => \N__11155\,
            DOUT => \N__11154\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11156\,
            PADOUT => \N__11155\,
            PADIN => \N__11154\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11147\,
            DIN => \N__11146\,
            DOUT => \N__11145\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11147\,
            PADOUT => \N__11146\,
            PADIN => \N__11145\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11138\,
            DIN => \N__11137\,
            DOUT => \N__11136\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11138\,
            PADOUT => \N__11137\,
            PADIN => \N__11136\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11129\,
            DIN => \N__11128\,
            DOUT => \N__11127\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11129\,
            PADOUT => \N__11128\,
            PADIN => \N__11127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11120\,
            DIN => \N__11119\,
            DOUT => \N__11118\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11120\,
            PADOUT => \N__11119\,
            PADIN => \N__11118\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11111\,
            DIN => \N__11110\,
            DOUT => \N__11109\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11111\,
            PADOUT => \N__11110\,
            PADIN => \N__11109\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11102\,
            DIN => \N__11101\,
            DOUT => \N__11100\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11102\,
            PADOUT => \N__11101\,
            PADIN => \N__11100\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11093\,
            DIN => \N__11092\,
            DOUT => \N__11091\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11093\,
            PADOUT => \N__11092\,
            PADIN => \N__11091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11084\,
            DIN => \N__11083\,
            DOUT => \N__11082\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11084\,
            PADOUT => \N__11083\,
            PADIN => \N__11082\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11075\,
            DIN => \N__11074\,
            DOUT => \N__11073\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11075\,
            PADOUT => \N__11074\,
            PADIN => \N__11073\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11066\,
            DIN => \N__11065\,
            DOUT => \N__11064\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11066\,
            PADOUT => \N__11065\,
            PADIN => \N__11064\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9565\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11057\,
            DIN => \N__11056\,
            DOUT => \N__11055\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11057\,
            PADOUT => \N__11056\,
            PADIN => \N__11055\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11048\,
            DIN => \N__11047\,
            DOUT => \N__11046\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11048\,
            PADOUT => \N__11047\,
            PADIN => \N__11046\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11039\,
            DIN => \N__11038\,
            DOUT => \N__11037\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11039\,
            PADOUT => \N__11038\,
            PADIN => \N__11037\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4408\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11030\,
            DIN => \N__11029\,
            DOUT => \N__11028\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11030\,
            PADOUT => \N__11029\,
            PADIN => \N__11028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11021\,
            DIN => \N__11020\,
            DOUT => \N__11019\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11021\,
            PADOUT => \N__11020\,
            PADIN => \N__11019\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4390\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11012\,
            DIN => \N__11011\,
            DOUT => \N__11010\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11012\,
            PADOUT => \N__11011\,
            PADIN => \N__11010\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__10993\,
            I => \N__10989\
        );

    \I__2673\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10977\
        );

    \I__2672\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10974\
        );

    \I__2671\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10971\
        );

    \I__2670\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10961\
        );

    \I__2669\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10961\
        );

    \I__2668\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10961\
        );

    \I__2667\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10961\
        );

    \I__2666\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10958\
        );

    \I__2665\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10955\
        );

    \I__2664\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10949\
        );

    \I__2663\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10949\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10942\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10942\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10942\
        );

    \I__2659\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10939\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10936\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10931\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10931\
        );

    \I__2655\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10928\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10917\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__10942\,
            I => \N__10914\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10911\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__10936\,
            I => \N__10904\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__10931\,
            I => \N__10904\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10904\
        );

    \I__2648\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10897\
        );

    \I__2647\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10897\
        );

    \I__2646\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10897\
        );

    \I__2645\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10894\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10891\
        );

    \I__2643\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10884\
        );

    \I__2642\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10884\
        );

    \I__2641\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10884\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__10917\,
            I => \N__10881\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__10914\,
            I => \N__10878\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__10911\,
            I => \N__10873\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__10904\,
            I => \N__10873\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10897\,
            I => \N__10866\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__10894\,
            I => \N__10866\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__10891\,
            I => \N__10866\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10863\
        );

    \I__2632\ : Sp12to4
    port map (
            O => \N__10881\,
            I => \N__10858\
        );

    \I__2631\ : Sp12to4
    port map (
            O => \N__10878\,
            I => \N__10858\
        );

    \I__2630\ : Sp12to4
    port map (
            O => \N__10873\,
            I => \N__10855\
        );

    \I__2629\ : Span12Mux_h
    port map (
            O => \N__10866\,
            I => \N__10852\
        );

    \I__2628\ : Span12Mux_v
    port map (
            O => \N__10863\,
            I => \N__10849\
        );

    \I__2627\ : Span12Mux_h
    port map (
            O => \N__10858\,
            I => \N__10846\
        );

    \I__2626\ : Span12Mux_v
    port map (
            O => \N__10855\,
            I => \N__10843\
        );

    \I__2625\ : Span12Mux_v
    port map (
            O => \N__10852\,
            I => \N__10838\
        );

    \I__2624\ : Span12Mux_h
    port map (
            O => \N__10849\,
            I => \N__10838\
        );

    \I__2623\ : Span12Mux_v
    port map (
            O => \N__10846\,
            I => \N__10833\
        );

    \I__2622\ : Span12Mux_h
    port map (
            O => \N__10843\,
            I => \N__10833\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__10838\,
            I => \AGNUS_REV_c\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__10833\,
            I => \AGNUS_REV_c\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10823\
        );

    \I__2618\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10819\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10816\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10813\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10810\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__10819\,
            I => \N__10805\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10816\,
            I => \N__10805\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__10813\,
            I => \N__10800\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10800\
        );

    \I__2610\ : Span4Mux_h
    port map (
            O => \N__10805\,
            I => \N__10797\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__2608\ : Sp12to4
    port map (
            O => \N__10797\,
            I => \N__10791\
        );

    \I__2607\ : Sp12to4
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__2606\ : Span12Mux_v
    port map (
            O => \N__10791\,
            I => \N__10785\
        );

    \I__2605\ : Span12Mux_h
    port map (
            O => \N__10788\,
            I => \N__10782\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__10785\,
            I => \DRA_c_6\
        );

    \I__2603\ : Odrv12
    port map (
            O => \N__10782\,
            I => \DRA_c_6\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10772\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10769\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10766\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10772\,
            I => \N__10762\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10769\,
            I => \N__10759\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10766\,
            I => \N__10756\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__10765\,
            I => \N__10753\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__10762\,
            I => \N__10750\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__10759\,
            I => \N__10745\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__10756\,
            I => \N__10745\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10742\
        );

    \I__2591\ : Sp12to4
    port map (
            O => \N__10750\,
            I => \N__10735\
        );

    \I__2590\ : Sp12to4
    port map (
            O => \N__10745\,
            I => \N__10735\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10735\
        );

    \I__2588\ : Span12Mux_h
    port map (
            O => \N__10735\,
            I => \N__10732\
        );

    \I__2587\ : Odrv12
    port map (
            O => \N__10732\,
            I => \DRA_c_7\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10726\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__10723\,
            I => \N__10720\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__10720\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2582\ : ClkMux
    port map (
            O => \N__10717\,
            I => \N__10702\
        );

    \I__2581\ : ClkMux
    port map (
            O => \N__10716\,
            I => \N__10702\
        );

    \I__2580\ : ClkMux
    port map (
            O => \N__10715\,
            I => \N__10702\
        );

    \I__2579\ : ClkMux
    port map (
            O => \N__10714\,
            I => \N__10702\
        );

    \I__2578\ : ClkMux
    port map (
            O => \N__10713\,
            I => \N__10702\
        );

    \I__2577\ : GlobalMux
    port map (
            O => \N__10702\,
            I => \N__10699\
        );

    \I__2576\ : gio2CtrlBuf
    port map (
            O => \N__10699\,
            I => \C3_c_g\
        );

    \I__2575\ : CEMux
    port map (
            O => \N__10696\,
            I => \N__10669\
        );

    \I__2574\ : CEMux
    port map (
            O => \N__10695\,
            I => \N__10669\
        );

    \I__2573\ : CEMux
    port map (
            O => \N__10694\,
            I => \N__10669\
        );

    \I__2572\ : CEMux
    port map (
            O => \N__10693\,
            I => \N__10669\
        );

    \I__2571\ : CEMux
    port map (
            O => \N__10692\,
            I => \N__10669\
        );

    \I__2570\ : CEMux
    port map (
            O => \N__10691\,
            I => \N__10669\
        );

    \I__2569\ : CEMux
    port map (
            O => \N__10690\,
            I => \N__10669\
        );

    \I__2568\ : CEMux
    port map (
            O => \N__10689\,
            I => \N__10669\
        );

    \I__2567\ : CEMux
    port map (
            O => \N__10688\,
            I => \N__10669\
        );

    \I__2566\ : GlobalMux
    port map (
            O => \N__10669\,
            I => \N__10666\
        );

    \I__2565\ : gio2CtrlBuf
    port map (
            O => \N__10666\,
            I => \DBRn_c_i_0_g\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10657\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10652\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10652\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10649\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10657\,
            I => \N__10636\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10629\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10622\
        );

    \I__2557\ : SRMux
    port map (
            O => \N__10648\,
            I => \N__10516\
        );

    \I__2556\ : SRMux
    port map (
            O => \N__10647\,
            I => \N__10516\
        );

    \I__2555\ : SRMux
    port map (
            O => \N__10646\,
            I => \N__10516\
        );

    \I__2554\ : SRMux
    port map (
            O => \N__10645\,
            I => \N__10516\
        );

    \I__2553\ : SRMux
    port map (
            O => \N__10644\,
            I => \N__10516\
        );

    \I__2552\ : SRMux
    port map (
            O => \N__10643\,
            I => \N__10516\
        );

    \I__2551\ : SRMux
    port map (
            O => \N__10642\,
            I => \N__10516\
        );

    \I__2550\ : SRMux
    port map (
            O => \N__10641\,
            I => \N__10516\
        );

    \I__2549\ : SRMux
    port map (
            O => \N__10640\,
            I => \N__10516\
        );

    \I__2548\ : SRMux
    port map (
            O => \N__10639\,
            I => \N__10516\
        );

    \I__2547\ : Glb2LocalMux
    port map (
            O => \N__10636\,
            I => \N__10516\
        );

    \I__2546\ : SRMux
    port map (
            O => \N__10635\,
            I => \N__10516\
        );

    \I__2545\ : SRMux
    port map (
            O => \N__10634\,
            I => \N__10516\
        );

    \I__2544\ : SRMux
    port map (
            O => \N__10633\,
            I => \N__10516\
        );

    \I__2543\ : SRMux
    port map (
            O => \N__10632\,
            I => \N__10516\
        );

    \I__2542\ : Glb2LocalMux
    port map (
            O => \N__10629\,
            I => \N__10516\
        );

    \I__2541\ : SRMux
    port map (
            O => \N__10628\,
            I => \N__10516\
        );

    \I__2540\ : SRMux
    port map (
            O => \N__10627\,
            I => \N__10516\
        );

    \I__2539\ : SRMux
    port map (
            O => \N__10626\,
            I => \N__10516\
        );

    \I__2538\ : SRMux
    port map (
            O => \N__10625\,
            I => \N__10516\
        );

    \I__2537\ : Glb2LocalMux
    port map (
            O => \N__10622\,
            I => \N__10516\
        );

    \I__2536\ : SRMux
    port map (
            O => \N__10621\,
            I => \N__10516\
        );

    \I__2535\ : SRMux
    port map (
            O => \N__10620\,
            I => \N__10516\
        );

    \I__2534\ : SRMux
    port map (
            O => \N__10619\,
            I => \N__10516\
        );

    \I__2533\ : SRMux
    port map (
            O => \N__10618\,
            I => \N__10516\
        );

    \I__2532\ : SRMux
    port map (
            O => \N__10617\,
            I => \N__10516\
        );

    \I__2531\ : SRMux
    port map (
            O => \N__10616\,
            I => \N__10516\
        );

    \I__2530\ : SRMux
    port map (
            O => \N__10615\,
            I => \N__10516\
        );

    \I__2529\ : SRMux
    port map (
            O => \N__10614\,
            I => \N__10516\
        );

    \I__2528\ : SRMux
    port map (
            O => \N__10613\,
            I => \N__10516\
        );

    \I__2527\ : SRMux
    port map (
            O => \N__10612\,
            I => \N__10516\
        );

    \I__2526\ : SRMux
    port map (
            O => \N__10611\,
            I => \N__10516\
        );

    \I__2525\ : SRMux
    port map (
            O => \N__10610\,
            I => \N__10516\
        );

    \I__2524\ : SRMux
    port map (
            O => \N__10609\,
            I => \N__10516\
        );

    \I__2523\ : SRMux
    port map (
            O => \N__10608\,
            I => \N__10516\
        );

    \I__2522\ : SRMux
    port map (
            O => \N__10607\,
            I => \N__10516\
        );

    \I__2521\ : SRMux
    port map (
            O => \N__10606\,
            I => \N__10516\
        );

    \I__2520\ : SRMux
    port map (
            O => \N__10605\,
            I => \N__10516\
        );

    \I__2519\ : SRMux
    port map (
            O => \N__10604\,
            I => \N__10516\
        );

    \I__2518\ : SRMux
    port map (
            O => \N__10603\,
            I => \N__10516\
        );

    \I__2517\ : SRMux
    port map (
            O => \N__10602\,
            I => \N__10516\
        );

    \I__2516\ : SRMux
    port map (
            O => \N__10601\,
            I => \N__10516\
        );

    \I__2515\ : GlobalMux
    port map (
            O => \N__10516\,
            I => \N__10513\
        );

    \I__2514\ : gio2CtrlBuf
    port map (
            O => \N__10513\,
            I => \RESETn_c_i_g\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10503\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10503\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10499\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10503\,
            I => \N__10496\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10493\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10499\,
            I => \N__10490\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__10496\,
            I => \N__10485\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10485\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__10490\,
            I => \N__10482\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__10485\,
            I => \N__10479\
        );

    \I__2503\ : Sp12to4
    port map (
            O => \N__10482\,
            I => \N__10476\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__10479\,
            I => \N__10473\
        );

    \I__2501\ : Span12Mux_h
    port map (
            O => \N__10476\,
            I => \N__10470\
        );

    \I__2500\ : Sp12to4
    port map (
            O => \N__10473\,
            I => \N__10467\
        );

    \I__2499\ : Span12Mux_v
    port map (
            O => \N__10470\,
            I => \N__10462\
        );

    \I__2498\ : Span12Mux_h
    port map (
            O => \N__10467\,
            I => \N__10462\
        );

    \I__2497\ : Odrv12
    port map (
            O => \N__10462\,
            I => \CASUn_c\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10451\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10451\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10457\,
            I => \N__10448\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10445\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10442\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10448\,
            I => \N__10439\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10445\,
            I => \N__10436\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__10442\,
            I => \N__10431\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__10439\,
            I => \N__10431\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10428\
        );

    \I__2486\ : Sp12to4
    port map (
            O => \N__10431\,
            I => \N__10425\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__2484\ : Span12Mux_h
    port map (
            O => \N__10425\,
            I => \N__10419\
        );

    \I__2483\ : Sp12to4
    port map (
            O => \N__10422\,
            I => \N__10416\
        );

    \I__2482\ : Span12Mux_v
    port map (
            O => \N__10419\,
            I => \N__10411\
        );

    \I__2481\ : Span12Mux_h
    port map (
            O => \N__10416\,
            I => \N__10411\
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__10411\,
            I => \CASLn_c\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10404\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10401\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10404\,
            I => \N__10396\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10396\
        );

    \I__2475\ : Odrv12
    port map (
            O => \N__10396\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10390\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10365\
        );

    \I__2472\ : ClkMux
    port map (
            O => \N__10389\,
            I => \N__10306\
        );

    \I__2471\ : ClkMux
    port map (
            O => \N__10388\,
            I => \N__10306\
        );

    \I__2470\ : ClkMux
    port map (
            O => \N__10387\,
            I => \N__10306\
        );

    \I__2469\ : ClkMux
    port map (
            O => \N__10386\,
            I => \N__10306\
        );

    \I__2468\ : ClkMux
    port map (
            O => \N__10385\,
            I => \N__10306\
        );

    \I__2467\ : ClkMux
    port map (
            O => \N__10384\,
            I => \N__10306\
        );

    \I__2466\ : ClkMux
    port map (
            O => \N__10383\,
            I => \N__10306\
        );

    \I__2465\ : ClkMux
    port map (
            O => \N__10382\,
            I => \N__10306\
        );

    \I__2464\ : ClkMux
    port map (
            O => \N__10381\,
            I => \N__10306\
        );

    \I__2463\ : ClkMux
    port map (
            O => \N__10380\,
            I => \N__10306\
        );

    \I__2462\ : ClkMux
    port map (
            O => \N__10379\,
            I => \N__10306\
        );

    \I__2461\ : ClkMux
    port map (
            O => \N__10378\,
            I => \N__10306\
        );

    \I__2460\ : ClkMux
    port map (
            O => \N__10377\,
            I => \N__10306\
        );

    \I__2459\ : ClkMux
    port map (
            O => \N__10376\,
            I => \N__10306\
        );

    \I__2458\ : ClkMux
    port map (
            O => \N__10375\,
            I => \N__10306\
        );

    \I__2457\ : ClkMux
    port map (
            O => \N__10374\,
            I => \N__10306\
        );

    \I__2456\ : ClkMux
    port map (
            O => \N__10373\,
            I => \N__10306\
        );

    \I__2455\ : ClkMux
    port map (
            O => \N__10372\,
            I => \N__10306\
        );

    \I__2454\ : ClkMux
    port map (
            O => \N__10371\,
            I => \N__10306\
        );

    \I__2453\ : ClkMux
    port map (
            O => \N__10370\,
            I => \N__10306\
        );

    \I__2452\ : ClkMux
    port map (
            O => \N__10369\,
            I => \N__10306\
        );

    \I__2451\ : ClkMux
    port map (
            O => \N__10368\,
            I => \N__10306\
        );

    \I__2450\ : Glb2LocalMux
    port map (
            O => \N__10365\,
            I => \N__10306\
        );

    \I__2449\ : ClkMux
    port map (
            O => \N__10364\,
            I => \N__10306\
        );

    \I__2448\ : ClkMux
    port map (
            O => \N__10363\,
            I => \N__10306\
        );

    \I__2447\ : ClkMux
    port map (
            O => \N__10362\,
            I => \N__10306\
        );

    \I__2446\ : ClkMux
    port map (
            O => \N__10361\,
            I => \N__10306\
        );

    \I__2445\ : GlobalMux
    port map (
            O => \N__10306\,
            I => \CLK80_PLL\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10297\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__10294\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10286\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10283\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10280\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10272\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10272\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10280\,
            I => \N__10272\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10269\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__10272\,
            I => \N__10266\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__2431\ : Sp12to4
    port map (
            O => \N__10266\,
            I => \N__10260\
        );

    \I__2430\ : Span12Mux_v
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__2429\ : Span12Mux_h
    port map (
            O => \N__10260\,
            I => \N__10254\
        );

    \I__2428\ : Span12Mux_h
    port map (
            O => \N__10257\,
            I => \N__10249\
        );

    \I__2427\ : Span12Mux_v
    port map (
            O => \N__10254\,
            I => \N__10249\
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__10249\,
            I => \DRA_c_2\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__10246\,
            I => \N__10243\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10240\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10240\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10225\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10220\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10220\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__10228\,
            I => \N__10215\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10215\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10220\,
            I => \N__10210\
        );

    \I__2414\ : Sp12to4
    port map (
            O => \N__10215\,
            I => \N__10210\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__10210\,
            I => \N__10207\
        );

    \I__2412\ : Span12Mux_h
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__10204\,
            I => \DRA_c_5\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10198\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10198\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10190\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10184\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10184\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10181\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10178\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10175\
        );

    \I__2402\ : Span4Mux_v
    port map (
            O => \N__10181\,
            I => \N__10172\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10169\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__10175\,
            I => \N__10166\
        );

    \I__2399\ : Sp12to4
    port map (
            O => \N__10172\,
            I => \N__10163\
        );

    \I__2398\ : Span12Mux_v
    port map (
            O => \N__10169\,
            I => \N__10158\
        );

    \I__2397\ : Sp12to4
    port map (
            O => \N__10166\,
            I => \N__10158\
        );

    \I__2396\ : Span12Mux_h
    port map (
            O => \N__10163\,
            I => \N__10155\
        );

    \I__2395\ : Span12Mux_h
    port map (
            O => \N__10158\,
            I => \N__10152\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__10155\,
            I => \DRA_c_8\
        );

    \I__2393\ : Odrv12
    port map (
            O => \N__10152\,
            I => \DRA_c_8\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10144\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10144\,
            I => \N__10141\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__10141\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__10138\,
            I => \N__10133\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10130\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10127\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10124\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10130\,
            I => \N__10121\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10117\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10114\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10121\,
            I => \N__10111\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10108\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10117\,
            I => \N__10103\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__10114\,
            I => \N__10103\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__10111\,
            I => \N__10100\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10097\
        );

    \I__2376\ : Sp12to4
    port map (
            O => \N__10103\,
            I => \N__10094\
        );

    \I__2375\ : Sp12to4
    port map (
            O => \N__10100\,
            I => \N__10089\
        );

    \I__2374\ : Span12Mux_v
    port map (
            O => \N__10097\,
            I => \N__10089\
        );

    \I__2373\ : Span12Mux_v
    port map (
            O => \N__10094\,
            I => \N__10086\
        );

    \I__2372\ : Span12Mux_h
    port map (
            O => \N__10089\,
            I => \N__10083\
        );

    \I__2371\ : Span12Mux_h
    port map (
            O => \N__10086\,
            I => \N__10078\
        );

    \I__2370\ : Span12Mux_v
    port map (
            O => \N__10083\,
            I => \N__10078\
        );

    \I__2369\ : Odrv12
    port map (
            O => \N__10078\,
            I => \DRA_c_9\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10072\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10069\
        );

    \I__2366\ : Span12Mux_h
    port map (
            O => \N__10069\,
            I => \N__10066\
        );

    \I__2365\ : Odrv12
    port map (
            O => \N__10066\,
            I => \RAS0n_c\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10054\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__10051\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10044\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10041\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10044\,
            I => \N__10038\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10041\,
            I => \N__10035\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10038\,
            I => \N__10028\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10035\,
            I => \N__10028\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10025\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10022\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__10028\,
            I => \N__10019\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10025\,
            I => \N__10014\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10022\,
            I => \N__10014\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__10019\,
            I => \N__10009\
        );

    \I__2347\ : Span12Mux_v
    port map (
            O => \N__10014\,
            I => \N__10009\
        );

    \I__2346\ : Span12Mux_h
    port map (
            O => \N__10009\,
            I => \N__10006\
        );

    \I__2345\ : Odrv12
    port map (
            O => \N__10006\,
            I => \DRA_c_3\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10003\,
            I => \N__9998\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10002\,
            I => \N__9994\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9991\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9988\
        );

    \I__2340\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9985\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9980\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__9991\,
            I => \N__9980\
        );

    \I__2337\ : Span4Mux_h
    port map (
            O => \N__9988\,
            I => \N__9975\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__9985\,
            I => \N__9975\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__9980\,
            I => \N__9972\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__9975\,
            I => \N__9969\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__9972\,
            I => \N__9966\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__9969\,
            I => \N__9963\
        );

    \I__2331\ : Sp12to4
    port map (
            O => \N__9966\,
            I => \N__9960\
        );

    \I__2330\ : Sp12to4
    port map (
            O => \N__9963\,
            I => \N__9957\
        );

    \I__2329\ : Span12Mux_h
    port map (
            O => \N__9960\,
            I => \N__9954\
        );

    \I__2328\ : Span12Mux_h
    port map (
            O => \N__9957\,
            I => \N__9951\
        );

    \I__2327\ : Odrv12
    port map (
            O => \N__9954\,
            I => \DRA_c_4\
        );

    \I__2326\ : Odrv12
    port map (
            O => \N__9951\,
            I => \DRA_c_4\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__9946\,
            I => \N__9943\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9940\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__9940\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2322\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9934\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__9931\,
            I => \N__9927\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9930\,
            I => \N__9924\
        );

    \I__2318\ : Sp12to4
    port map (
            O => \N__9927\,
            I => \N__9921\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9924\,
            I => \N__9918\
        );

    \I__2316\ : Span12Mux_h
    port map (
            O => \N__9921\,
            I => \N__9915\
        );

    \I__2315\ : Span12Mux_h
    port map (
            O => \N__9918\,
            I => \N__9912\
        );

    \I__2314\ : Span12Mux_v
    port map (
            O => \N__9915\,
            I => \N__9909\
        );

    \I__2313\ : Span12Mux_v
    port map (
            O => \N__9912\,
            I => \N__9906\
        );

    \I__2312\ : Odrv12
    port map (
            O => \N__9909\,
            I => \DRA_c_0\
        );

    \I__2311\ : Odrv12
    port map (
            O => \N__9906\,
            I => \DRA_c_0\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9897\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9890\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9894\,
            I => \N__9886\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9883\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__9890\,
            I => \N__9880\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9877\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__9886\,
            I => \N__9872\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9883\,
            I => \N__9872\
        );

    \I__2301\ : Sp12to4
    port map (
            O => \N__9880\,
            I => \N__9867\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9877\,
            I => \N__9867\
        );

    \I__2299\ : Sp12to4
    port map (
            O => \N__9872\,
            I => \N__9864\
        );

    \I__2298\ : Span12Mux_h
    port map (
            O => \N__9867\,
            I => \N__9861\
        );

    \I__2297\ : Span12Mux_v
    port map (
            O => \N__9864\,
            I => \N__9858\
        );

    \I__2296\ : Span12Mux_v
    port map (
            O => \N__9861\,
            I => \N__9855\
        );

    \I__2295\ : Span12Mux_h
    port map (
            O => \N__9858\,
            I => \N__9852\
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__9855\,
            I => \DRA_c_1\
        );

    \I__2293\ : Odrv12
    port map (
            O => \N__9852\,
            I => \DRA_c_1\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9844\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9844\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__9841\,
            I => \N__9833\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9828\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9828\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9821\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9821\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9821\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9818\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9828\,
            I => \N__9809\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9809\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9809\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9803\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9803\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9800\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9797\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9803\,
            I => \N__9794\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__9800\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9797\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__9794\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9784\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__9781\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2269\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9767\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9767\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9767\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9762\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9762\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9767\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9762\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2262\ : IoInMux
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__2260\ : Span4Mux_s2_h
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__2259\ : Sp12to4
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__2258\ : Span12Mux_v
    port map (
            O => \N__9745\,
            I => \N__9742\
        );

    \I__2257\ : Span12Mux_h
    port map (
            O => \N__9742\,
            I => \N__9739\
        );

    \I__2256\ : Odrv12
    port map (
            O => \N__9739\,
            I => \CMA_c_3\
        );

    \I__2255\ : CEMux
    port map (
            O => \N__9736\,
            I => \N__9732\
        );

    \I__2254\ : CEMux
    port map (
            O => \N__9735\,
            I => \N__9729\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9722\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9719\
        );

    \I__2251\ : CEMux
    port map (
            O => \N__9728\,
            I => \N__9716\
        );

    \I__2250\ : CEMux
    port map (
            O => \N__9727\,
            I => \N__9713\
        );

    \I__2249\ : CEMux
    port map (
            O => \N__9726\,
            I => \N__9710\
        );

    \I__2248\ : CEMux
    port map (
            O => \N__9725\,
            I => \N__9707\
        );

    \I__2247\ : Span4Mux_h
    port map (
            O => \N__9722\,
            I => \N__9702\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__9719\,
            I => \N__9702\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9716\,
            I => \N__9697\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__9713\,
            I => \N__9697\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__9710\,
            I => \N__9694\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9691\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__9702\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__9697\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__9694\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__9691\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9679\,
            I => \N__9676\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__9673\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9664\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__9661\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9655\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9652\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__9652\,
            I => \N__9649\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__9649\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9643\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__9640\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9634\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__9631\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__9622\,
            I => \N__9619\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__9619\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__9607\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2211\ : IoInMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__2209\ : Span4Mux_s2_v
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__9595\,
            I => \N__9592\
        );

    \I__2207\ : Sp12to4
    port map (
            O => \N__9592\,
            I => \N__9589\
        );

    \I__2206\ : Span12Mux_h
    port map (
            O => \N__9589\,
            I => \N__9586\
        );

    \I__2205\ : Odrv12
    port map (
            O => \N__9586\,
            I => \CASn_c\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9577\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9574\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__9574\,
            I => \N__9571\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__9571\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__9568\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\
        );

    \I__2198\ : IoInMux
    port map (
            O => \N__9565\,
            I => \N__9562\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9562\,
            I => \N__9559\
        );

    \I__2196\ : Span4Mux_s3_h
    port map (
            O => \N__9559\,
            I => \N__9556\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__9556\,
            I => \N__9553\
        );

    \I__2194\ : Span12Mux_s10_v
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__2193\ : Span12Mux_h
    port map (
            O => \N__9550\,
            I => \N__9547\
        );

    \I__2192\ : Odrv12
    port map (
            O => \N__9547\,
            I => \CMA_c_6\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9541\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9541\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2189\ : IoInMux
    port map (
            O => \N__9538\,
            I => \N__9535\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9535\,
            I => \N__9532\
        );

    \I__2187\ : IoSpan4Mux
    port map (
            O => \N__9532\,
            I => \N__9529\
        );

    \I__2186\ : Span4Mux_s2_h
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__2185\ : Sp12to4
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__2184\ : Span12Mux_h
    port map (
            O => \N__9523\,
            I => \N__9520\
        );

    \I__2183\ : Odrv12
    port map (
            O => \N__9520\,
            I => \CMA_c_4\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9514\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9514\,
            I => \N__9511\
        );

    \I__2180\ : Span4Mux_h
    port map (
            O => \N__9511\,
            I => \N__9508\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__9508\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__9505\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\
        );

    \I__2177\ : IoInMux
    port map (
            O => \N__9502\,
            I => \N__9499\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9496\
        );

    \I__2175\ : IoSpan4Mux
    port map (
            O => \N__9496\,
            I => \N__9493\
        );

    \I__2174\ : Span4Mux_s2_h
    port map (
            O => \N__9493\,
            I => \N__9490\
        );

    \I__2173\ : Sp12to4
    port map (
            O => \N__9490\,
            I => \N__9487\
        );

    \I__2172\ : Span12Mux_h
    port map (
            O => \N__9487\,
            I => \N__9484\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__9484\,
            I => \CMA_c_7\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9478\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9478\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__2168\ : IoInMux
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__2166\ : IoSpan4Mux
    port map (
            O => \N__9469\,
            I => \N__9466\
        );

    \I__2165\ : Span4Mux_s2_v
    port map (
            O => \N__9466\,
            I => \N__9463\
        );

    \I__2164\ : Sp12to4
    port map (
            O => \N__9463\,
            I => \N__9460\
        );

    \I__2163\ : Odrv12
    port map (
            O => \N__9460\,
            I => \CMA_c_2\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9443\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9443\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__9455\,
            I => \N__9438\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__9454\,
            I => \N__9434\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__9453\,
            I => \N__9431\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9425\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9425\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9420\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9417\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9414\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9408\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9403\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9403\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9398\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9398\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9393\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9393\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9390\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9387\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9384\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9381\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9420\,
            I => \N__9374\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9369\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9369\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9364\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9364\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9361\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9408\,
            I => \N__9358\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9349\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9398\,
            I => \N__9349\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9349\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9390\,
            I => \N__9349\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__9387\,
            I => \N__9342\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9384\,
            I => \N__9342\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9381\,
            I => \N__9342\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9337\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9337\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9332\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9332\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__9374\,
            I => \N__9323\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__9369\,
            I => \N__9323\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9323\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9361\,
            I => \N__9323\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__9358\,
            I => \N__9320\
        );

    \I__2118\ : Span4Mux_h
    port map (
            O => \N__9349\,
            I => \N__9317\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__9342\,
            I => \N__9310\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9337\,
            I => \N__9310\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9310\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__9323\,
            I => \CPU_CYCLE\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__9320\,
            I => \CPU_CYCLE\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__9317\,
            I => \CPU_CYCLE\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__9310\,
            I => \CPU_CYCLE\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9293\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9288\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9288\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__9298\,
            I => \N__9285\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9282\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9278\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9275\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9272\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9269\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9282\,
            I => \N__9266\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__9281\,
            I => \N__9263\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9278\,
            I => \N__9256\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9256\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__9272\,
            I => \N__9240\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9240\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__9266\,
            I => \N__9233\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9228\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9228\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9225\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9256\,
            I => \N__9222\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9213\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9213\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9213\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9213\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9204\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9204\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9204\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9204\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9199\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9199\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9196\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__9240\,
            I => \N__9193\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9186\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9186\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9186\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9183\
        );

    \I__2074\ : Sp12to4
    port map (
            O => \N__9233\,
            I => \N__9168\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9168\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9225\,
            I => \N__9168\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__9222\,
            I => \N__9168\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N__9168\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9168\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9168\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9196\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__9193\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9186\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9183\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__9168\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9151\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__2059\ : IoInMux
    port map (
            O => \N__9148\,
            I => \N__9145\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__2057\ : Span4Mux_s3_v
    port map (
            O => \N__9142\,
            I => \N__9139\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__9136\,
            I => \N__9133\
        );

    \I__2054\ : Span4Mux_h
    port map (
            O => \N__9133\,
            I => \N__9130\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__9130\,
            I => \CMA_c_0\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__9127\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9121\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9121\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__9112\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9103\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__9097\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9090\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9087\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9082\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9073\
        );

    \I__2037\ : ClkMux
    port map (
            O => \N__9086\,
            I => \N__9052\
        );

    \I__2036\ : ClkMux
    port map (
            O => \N__9085\,
            I => \N__9052\
        );

    \I__2035\ : Glb2LocalMux
    port map (
            O => \N__9082\,
            I => \N__9052\
        );

    \I__2034\ : ClkMux
    port map (
            O => \N__9081\,
            I => \N__9052\
        );

    \I__2033\ : ClkMux
    port map (
            O => \N__9080\,
            I => \N__9052\
        );

    \I__2032\ : ClkMux
    port map (
            O => \N__9079\,
            I => \N__9052\
        );

    \I__2031\ : ClkMux
    port map (
            O => \N__9078\,
            I => \N__9052\
        );

    \I__2030\ : ClkMux
    port map (
            O => \N__9077\,
            I => \N__9052\
        );

    \I__2029\ : ClkMux
    port map (
            O => \N__9076\,
            I => \N__9052\
        );

    \I__2028\ : Glb2LocalMux
    port map (
            O => \N__9073\,
            I => \N__9052\
        );

    \I__2027\ : GlobalMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__2026\ : gio2CtrlBuf
    port map (
            O => \N__9049\,
            I => \CLK40_PLL_g\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9040\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9040\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9040\,
            I => \N__9033\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9028\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9028\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9025\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9022\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__9033\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9028\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9025\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9022\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__9013\,
            I => \N__9010\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9010\,
            I => \N__9007\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9007\,
            I => \U712_CYCLE_TERM.N_8\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__9004\,
            I => \N__9000\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8996\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8986\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8986\
        );

    \I__2007\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8981\
        );

    \I__2006\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8981\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8978\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8968\
        );

    \I__2003\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8968\
        );

    \I__2002\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8968\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__8986\,
            I => \N__8965\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8960\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8960\
        );

    \I__1998\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8957\
        );

    \I__1997\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8954\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8951\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8968\,
            I => \N__8946\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__8965\,
            I => \N__8937\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__8960\,
            I => \N__8937\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8937\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8954\,
            I => \N__8937\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8933\
        );

    \I__1989\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8928\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8928\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__8946\,
            I => \N__8925\
        );

    \I__1986\ : Span4Mux_v
    port map (
            O => \N__8937\,
            I => \N__8922\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8919\
        );

    \I__1984\ : Sp12to4
    port map (
            O => \N__8933\,
            I => \N__8914\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8928\,
            I => \N__8914\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__8925\,
            I => \N__8907\
        );

    \I__1981\ : Sp12to4
    port map (
            O => \N__8922\,
            I => \N__8907\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8907\
        );

    \I__1979\ : Span12Mux_v
    port map (
            O => \N__8914\,
            I => \N__8904\
        );

    \I__1978\ : Span12Mux_h
    port map (
            O => \N__8907\,
            I => \N__8901\
        );

    \I__1977\ : Span12Mux_h
    port map (
            O => \N__8904\,
            I => \N__8898\
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__8901\,
            I => \RESETn_c\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__8898\,
            I => \RESETn_c\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8888\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8885\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8882\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8888\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8885\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8882\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8871\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8868\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8871\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8868\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__8863\,
            I => \N__8858\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__8862\,
            I => \N__8855\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8851\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8848\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8845\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8842\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8851\,
            I => \N__8838\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8848\,
            I => \N__8835\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8845\,
            I => \N__8830\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8842\,
            I => \N__8830\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8827\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__8838\,
            I => \N__8824\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__8835\,
            I => \N__8821\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__8830\,
            I => \N__8818\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8827\,
            I => \CPU_TACK\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__8824\,
            I => \CPU_TACK\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__8821\,
            I => \CPU_TACK\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__8818\,
            I => \CPU_TACK\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__8809\,
            I => \U712_CYCLE_TERM.N_227_i_0_0_cascade_\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__8806\,
            I => \N__8801\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8796\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8793\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8790\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8785\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8785\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8796\,
            I => \N__8780\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8780\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8790\,
            I => \REG_TACK\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8785\,
            I => \REG_TACK\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8780\,
            I => \REG_TACK\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__8773\,
            I => \U712_CYCLE_TERM.N_227_i_0_en_cascade_\
        );

    \I__1933\ : IoInMux
    port map (
            O => \N__8770\,
            I => \N__8767\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8764\
        );

    \I__1931\ : Span12Mux_s1_v
    port map (
            O => \N__8764\,
            I => \N__8760\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8757\
        );

    \I__1929\ : Odrv12
    port map (
            O => \N__8760\,
            I => \RESETn_c_i\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8757\,
            I => \RESETn_c_i\
        );

    \I__1927\ : CEMux
    port map (
            O => \N__8752\,
            I => \N__8749\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8746\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__8746\,
            I => \U712_CYCLE_TERM.N_227_i_0_en_0\
        );

    \I__1924\ : IoInMux
    port map (
            O => \N__8743\,
            I => \N__8740\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8740\,
            I => \N__8737\
        );

    \I__1922\ : Span4Mux_s2_v
    port map (
            O => \N__8737\,
            I => \N__8734\
        );

    \I__1921\ : Sp12to4
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__1920\ : Span12Mux_h
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__1919\ : Odrv12
    port map (
            O => \N__8728\,
            I => \CRCSn_c\
        );

    \I__1918\ : IoInMux
    port map (
            O => \N__8725\,
            I => \N__8722\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__1916\ : Span4Mux_s2_v
    port map (
            O => \N__8719\,
            I => \N__8716\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__8713\,
            I => \N__8710\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__8710\,
            I => \N__8707\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__8707\,
            I => \CMA_c_10\
        );

    \I__1911\ : IoInMux
    port map (
            O => \N__8704\,
            I => \N__8700\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8697\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8700\,
            I => \N__8694\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8691\
        );

    \I__1907\ : Span12Mux_s11_v
    port map (
            O => \N__8694\,
            I => \N__8688\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__8691\,
            I => \N__8685\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__8688\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__8685\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8677\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8677\,
            I => \N__8674\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__8674\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8668\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8668\,
            I => \N__8665\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__8665\,
            I => \N__8662\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__8662\,
            I => \N__8659\
        );

    \I__1896\ : Sp12to4
    port map (
            O => \N__8659\,
            I => \N__8656\
        );

    \I__1895\ : Span12Mux_h
    port map (
            O => \N__8656\,
            I => \N__8653\
        );

    \I__1894\ : Odrv12
    port map (
            O => \N__8653\,
            I => \A_c_6\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8647\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1891\ : Span12Mux_v
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1890\ : Span12Mux_h
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1889\ : Odrv12
    port map (
            O => \N__8638\,
            I => \A_c_13\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__8635\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__8632\,
            I => \N__8629\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8626\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8626\,
            I => \N__8623\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__8623\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8615\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8612\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8608\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8601\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8612\,
            I => \N__8601\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8597\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8594\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8591\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8588\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__8601\,
            I => \N__8585\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8582\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8597\,
            I => \N__8575\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__8594\,
            I => \N__8575\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8575\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8588\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__8585\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8582\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8575\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__8566\,
            I => \N__8561\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8558\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__8564\,
            I => \N__8555\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8551\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8548\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8545\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__8554\,
            I => \N__8542\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8538\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__8548\,
            I => \N__8535\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8532\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8529\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8526\
        );

    \I__1853\ : Span12Mux_h
    port map (
            O => \N__8538\,
            I => \N__8523\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__8535\,
            I => \N__8520\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8532\,
            I => \N__8515\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8515\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8526\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1848\ : Odrv12
    port map (
            O => \N__8523\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__8520\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__8515\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8501\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8498\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8494\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8501\,
            I => \N__8486\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8486\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8483\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8480\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8475\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8475\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8472\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__8486\,
            I => \N__8469\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8483\,
            I => \N__8460\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__8480\,
            I => \N__8460\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8460\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8460\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__8469\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__8460\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__8455\,
            I => \N__8450\
        );

    \I__1827\ : IoInMux
    port map (
            O => \N__8454\,
            I => \N__8447\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8442\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8442\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8447\,
            I => \N__8439\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8442\,
            I => \N__8436\
        );

    \I__1822\ : Span12Mux_s3_h
    port map (
            O => \N__8439\,
            I => \N__8433\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__8436\,
            I => \N__8430\
        );

    \I__1820\ : Span12Mux_v
    port map (
            O => \N__8433\,
            I => \N__8427\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__1818\ : Span12Mux_h
    port map (
            O => \N__8427\,
            I => \N__8421\
        );

    \I__1817\ : Span12Mux_v
    port map (
            O => \N__8424\,
            I => \N__8418\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__8421\,
            I => \CLK40_PLL\
        );

    \I__1815\ : Odrv12
    port map (
            O => \N__8418\,
            I => \CLK40_PLL\
        );

    \I__1814\ : IoInMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__1812\ : IoSpan4Mux
    port map (
            O => \N__8407\,
            I => \N__8404\
        );

    \I__1811\ : Span4Mux_s2_h
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__1810\ : Sp12to4
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__1809\ : Span12Mux_h
    port map (
            O => \N__8398\,
            I => \N__8394\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8391\
        );

    \I__1807\ : Odrv12
    port map (
            O => \N__8394\,
            I => \TACK_OUTn\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8391\,
            I => \TACK_OUTn\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8382\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8379\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8382\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8379\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8366\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8363\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8360\
        );

    \I__1797\ : Odrv12
    port map (
            O => \N__8366\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8363\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8360\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8350\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8341\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8341\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8335\,
            I => \TACK_EN_i_ess\
        );

    \I__1787\ : IoInMux
    port map (
            O => \N__8332\,
            I => \N__8329\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__1785\ : IoSpan4Mux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__1784\ : Sp12to4
    port map (
            O => \N__8323\,
            I => \N__8320\
        );

    \I__1783\ : Span12Mux_s9_v
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__8317\,
            I => \RASn_c\
        );

    \I__1781\ : IoInMux
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8308\
        );

    \I__1779\ : Span12Mux_s4_h
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__8302\,
            I => \WEn_c\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__8299\,
            I => \N__8295\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8290\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8290\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__8287\,
            I => \N__8282\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8277\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8277\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__8282\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8277\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8269\,
            I => \N__8266\
        );

    \I__1765\ : Sp12to4
    port map (
            O => \N__8266\,
            I => \N__8263\
        );

    \I__1764\ : Span12Mux_v
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1763\ : Span12Mux_h
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__8257\,
            I => \A_c_19\
        );

    \I__1761\ : IoInMux
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8251\,
            I => \N__8248\
        );

    \I__1759\ : Span12Mux_s5_h
    port map (
            O => \N__8248\,
            I => \N__8245\
        );

    \I__1758\ : Span12Mux_h
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__1757\ : Odrv12
    port map (
            O => \N__8242\,
            I => \CMA_c_9\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8236\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8236\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1754\ : IoInMux
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1752\ : IoSpan4Mux
    port map (
            O => \N__8227\,
            I => \N__8224\
        );

    \I__1751\ : Span4Mux_s3_h
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1750\ : Sp12to4
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__1749\ : Span12Mux_h
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__8215\,
            I => \CMA_c_5\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8209\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8203\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8197\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8188\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8182\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8182\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1736\ : IoInMux
    port map (
            O => \N__8179\,
            I => \N__8176\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__1734\ : Span4Mux_s3_v
    port map (
            O => \N__8173\,
            I => \N__8170\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__8170\,
            I => \N__8167\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__8164\,
            I => \CMA_c_1\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__8155\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__8146\,
            I => \N__8143\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__8143\,
            I => \DBRn_c_i\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8136\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8133\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8136\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8133\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8124\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8121\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8124\,
            I => \N__8117\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8114\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8111\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8117\,
            I => \N__8108\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__8114\,
            I => \N__8103\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8111\,
            I => \N__8103\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8108\,
            I => \N__8098\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8103\,
            I => \N__8098\
        );

    \I__1709\ : Sp12to4
    port map (
            O => \N__8098\,
            I => \N__8095\
        );

    \I__1708\ : Span12Mux_h
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__8092\,
            I => \DBRn_c\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8086\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8086\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_0\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8079\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8075\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8079\,
            I => \N__8072\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__8078\,
            I => \N__8069\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8064\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__8072\,
            I => \N__8064\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8069\,
            I => \N__8061\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__8064\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8061\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8049\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8052\,
            I => \N__8046\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8049\,
            I => \N__8042\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N__8039\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8036\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__8042\,
            I => \REG_CYCLE\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__8039\,
            I => \REG_CYCLE\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8036\,
            I => \REG_CYCLE\
        );

    \I__1686\ : IoInMux
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8026\,
            I => \N__8023\
        );

    \I__1684\ : Span4Mux_s0_v
    port map (
            O => \N__8023\,
            I => \N__8020\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__8017\,
            I => \N__8014\
        );

    \I__1681\ : Sp12to4
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__1680\ : Span12Mux_s11_h
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8008\,
            I => \DRDENn_c\
        );

    \I__1678\ : IoInMux
    port map (
            O => \N__8005\,
            I => \N__8002\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1676\ : IoSpan4Mux
    port map (
            O => \N__7999\,
            I => \N__7996\
        );

    \I__1675\ : Span4Mux_s3_v
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__7990\,
            I => \N_118_i\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7978\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7975\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7972\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7969\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7964\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7964\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7961\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7957\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7975\,
            I => \N__7950\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7972\,
            I => \N__7950\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7969\,
            I => \N__7950\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7964\,
            I => \N__7945\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7945\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7942\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7957\,
            I => \N__7937\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__7950\,
            I => \N__7937\
        );

    \I__1656\ : Span4Mux_h
    port map (
            O => \N__7945\,
            I => \N__7932\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7942\,
            I => \N__7932\
        );

    \I__1654\ : Span4Mux_h
    port map (
            O => \N__7937\,
            I => \N__7929\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7932\,
            I => \N__7926\
        );

    \I__1652\ : Sp12to4
    port map (
            O => \N__7929\,
            I => \N__7921\
        );

    \I__1651\ : Sp12to4
    port map (
            O => \N__7926\,
            I => \N__7921\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__7921\,
            I => \A_c_0\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__7918\,
            I => \N__7915\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__1647\ : Span4Mux_s3_v
    port map (
            O => \N__7912\,
            I => \N__7909\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__7906\,
            I => \U712_BYTE_ENABLE_UUBE_i\
        );

    \I__1644\ : IoInMux
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1642\ : Span4Mux_s2_v
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__7888\,
            I => \LLBEn_c\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7881\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7878\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7871\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7871\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7866\
        );

    \I__1633\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7866\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__7871\,
            I => \N__7861\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7861\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__7861\,
            I => \N_386\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__7858\,
            I => \N__7854\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7851\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7854\,
            I => \N__7848\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7851\,
            I => \N__7840\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7848\,
            I => \N__7840\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7835\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7835\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7832\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__7840\,
            I => \N__7826\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7826\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7832\,
            I => \N__7823\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7820\
        );

    \I__1617\ : Span4Mux_h
    port map (
            O => \N__7826\,
            I => \N__7817\
        );

    \I__1616\ : Span12Mux_h
    port map (
            O => \N__7823\,
            I => \N__7814\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7811\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__7817\,
            I => \N__7808\
        );

    \I__1613\ : Span12Mux_v
    port map (
            O => \N__7814\,
            I => \N__7805\
        );

    \I__1612\ : Span12Mux_v
    port map (
            O => \N__7811\,
            I => \N__7800\
        );

    \I__1611\ : Sp12to4
    port map (
            O => \N__7808\,
            I => \N__7800\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__7805\,
            I => \SIZ_c_0\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__7800\,
            I => \SIZ_c_0\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7787\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7794\,
            I => \N__7780\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7780\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7780\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__7791\,
            I => \N__7776\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__7790\,
            I => \N__7773\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7770\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7767\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7760\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7760\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7760\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__7770\,
            I => \N__7757\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__7767\,
            I => \N__7754\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7751\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__7757\,
            I => \N__7747\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7754\,
            I => \N__7742\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__7751\,
            I => \N__7742\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7739\
        );

    \I__1590\ : Sp12to4
    port map (
            O => \N__7747\,
            I => \N__7732\
        );

    \I__1589\ : Sp12to4
    port map (
            O => \N__7742\,
            I => \N__7732\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7739\,
            I => \N__7732\
        );

    \I__1587\ : Span12Mux_h
    port map (
            O => \N__7732\,
            I => \N__7729\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__7729\,
            I => \A_c_1\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7719\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7716\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__7719\,
            I => \N__7712\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7716\,
            I => \N__7705\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7702\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__7712\,
            I => \N__7699\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7696\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7693\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7688\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7688\
        );

    \I__1574\ : Sp12to4
    port map (
            O => \N__7705\,
            I => \N__7683\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7702\,
            I => \N__7683\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__7699\,
            I => \N__7680\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7673\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7693\,
            I => \N__7673\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7673\
        );

    \I__1568\ : Span12Mux_h
    port map (
            O => \N__7683\,
            I => \N__7670\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__7680\,
            I => \N__7665\
        );

    \I__1566\ : Span12Mux_v
    port map (
            O => \N__7673\,
            I => \N__7665\
        );

    \I__1565\ : Span12Mux_v
    port map (
            O => \N__7670\,
            I => \N__7660\
        );

    \I__1564\ : Span12Mux_h
    port map (
            O => \N__7665\,
            I => \N__7660\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__7660\,
            I => \SIZ_c_1\
        );

    \I__1562\ : IoInMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__1560\ : Span4Mux_s2_v
    port map (
            O => \N__7651\,
            I => \N__7648\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__7648\,
            I => \N__7645\
        );

    \I__1558\ : Sp12to4
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__7642\,
            I => \UMBEn_c\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7636\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7636\,
            I => \N__7633\
        );

    \I__1554\ : Sp12to4
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__1553\ : Span12Mux_v
    port map (
            O => \N__7630\,
            I => \N__7627\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__7627\,
            I => \N__7624\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7624\,
            I => \A_c_17\
        );

    \I__1550\ : IoInMux
    port map (
            O => \N__7621\,
            I => \N__7618\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7618\,
            I => \N__7615\
        );

    \I__1548\ : IoSpan4Mux
    port map (
            O => \N__7615\,
            I => \N__7612\
        );

    \I__1547\ : Span4Mux_s3_h
    port map (
            O => \N__7612\,
            I => \N__7609\
        );

    \I__1546\ : Sp12to4
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1545\ : Span12Mux_h
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1544\ : Odrv12
    port map (
            O => \N__7603\,
            I => \CMA_c_8\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__7600\,
            I => \N__7596\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7590\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7587\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7584\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7581\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7593\,
            I => \N__7578\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7590\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7587\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7584\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7581\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7578\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7563\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7559\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7563\,
            I => \N__7556\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7552\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7549\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__7556\,
            I => \N__7546\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7543\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7552\,
            I => \N__7540\
        );

    \I__1524\ : Sp12to4
    port map (
            O => \N__7549\,
            I => \N__7533\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__7546\,
            I => \N__7533\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7543\,
            I => \N__7533\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7540\,
            I => \N__7530\
        );

    \I__1520\ : Span12Mux_h
    port map (
            O => \N__7533\,
            I => \N__7527\
        );

    \I__1519\ : Sp12to4
    port map (
            O => \N__7530\,
            I => \N__7524\
        );

    \I__1518\ : Span12Mux_v
    port map (
            O => \N__7527\,
            I => \N__7521\
        );

    \I__1517\ : Span12Mux_h
    port map (
            O => \N__7524\,
            I => \N__7518\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__7521\,
            I => \RnW_c\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__7518\,
            I => \RnW_c\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__7507\,
            I => \U712_REG_SM.UDSn_7_iv_i_0\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7501\,
            I => \U712_REG_SM.N_245\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7495\,
            I => \U712_REG_SM.un15_0_i_0_0_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7487\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7482\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7482\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7487\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7482\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7468\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7473\,
            I => \N__7463\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7472\,
            I => \N__7459\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7456\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7468\,
            I => \N__7453\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7448\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7448\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7445\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7440\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7440\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7456\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__7453\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7448\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7445\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7440\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__7429\,
            I => \N__7424\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7421\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7418\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7415\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7421\,
            I => \N__7412\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7418\,
            I => \U712_REG_SM.N_209\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7415\,
            I => \U712_REG_SM.N_209\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__7412\,
            I => \U712_REG_SM.N_209\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7397\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7394\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7391\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7397\,
            I => \U712_REG_SM.N_229\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7394\,
            I => \U712_REG_SM.N_229\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7391\,
            I => \U712_REG_SM.N_229\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__7384\,
            I => \N__7378\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__7383\,
            I => \N__7373\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7369\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7366\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7363\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7360\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7355\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7355\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7352\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7369\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7360\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7355\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7352\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7331\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7328\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7325\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7331\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7328\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7325\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1449\ : IoInMux
    port map (
            O => \N__7318\,
            I => \N__7315\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7315\,
            I => \N__7312\
        );

    \I__1447\ : Span4Mux_s1_h
    port map (
            O => \N__7312\,
            I => \N__7309\
        );

    \I__1446\ : Sp12to4
    port map (
            O => \N__7309\,
            I => \N__7306\
        );

    \I__1445\ : Span12Mux_v
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__1444\ : Span12Mux_h
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__7300\,
            I => \N_858_i\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7297\,
            I => \N__7294\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7285\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7282\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7277\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7277\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7272\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7272\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7269\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7285\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7282\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7277\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7272\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7269\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7247\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7242\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7242\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7237\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7237\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7234\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7247\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7242\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7237\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7234\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__7225\,
            I => \N__7220\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7224\,
            I => \N__7213\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7210\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7207\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7204\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7197\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7197\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7197\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7194\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7191\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7204\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7197\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7194\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__7191\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7177\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7177\,
            I => \N__7172\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7169\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7166\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__7172\,
            I => \U712_REG_SM.REG_TACK_0_sqmuxa\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7169\,
            I => \U712_REG_SM.REG_TACK_0_sqmuxa\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7166\,
            I => \U712_REG_SM.REG_TACK_0_sqmuxa\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__7159\,
            I => \U712_BYTE_ENABLE.N_319_cascade_\
        );

    \I__1395\ : IoInMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1393\ : IoSpan4Mux
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__1392\ : Span4Mux_s2_h
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1391\ : Span4Mux_h
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1390\ : Sp12to4
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1389\ : Span12Mux_h
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1388\ : Span12Mux_v
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1387\ : Odrv12
    port map (
            O => \N__7132\,
            I => \N_58_i\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7126\,
            I => \U712_BYTE_ENABLE.N_320\
        );

    \I__1384\ : IoInMux
    port map (
            O => \N__7123\,
            I => \N__7120\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7117\
        );

    \I__1382\ : Span4Mux_s3_h
    port map (
            O => \N__7117\,
            I => \N__7114\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__7114\,
            I => \N__7111\
        );

    \I__1380\ : Sp12to4
    port map (
            O => \N__7111\,
            I => \N__7108\
        );

    \I__1379\ : Span12Mux_h
    port map (
            O => \N__7108\,
            I => \N__7105\
        );

    \I__1378\ : Span12Mux_v
    port map (
            O => \N__7105\,
            I => \N__7102\
        );

    \I__1377\ : Odrv12
    port map (
            O => \N__7102\,
            I => \N_56_i\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7093\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7093\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7093\,
            I => \U712_BYTE_ENABLE.N_318\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__7090\,
            I => \U712_BYTE_ENABLE.N_323_cascade_\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7081\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7081\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\
        );

    \I__1369\ : IoInMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1367\ : Span4Mux_s1_v
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1365\ : Span4Mux_v
    port map (
            O => \N__7066\,
            I => \N__7063\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__7057\,
            I => \N_54_i\
        );

    \I__1361\ : IoInMux
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7047\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__7050\,
            I => \N__7041\
        );

    \I__1358\ : IoSpan4Mux
    port map (
            O => \N__7047\,
            I => \N__7038\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7029\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7029\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7029\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7029\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__7038\,
            I => \N__7026\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7029\,
            I => \N__7023\
        );

    \I__1351\ : Span12Mux_s7_v
    port map (
            O => \N__7026\,
            I => \N__7019\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__7023\,
            I => \N__7016\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7013\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__7019\,
            I => \DBENn_c\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7016\,
            I => \DBENn_c\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7013\,
            I => \DBENn_c\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7006\,
            I => \N__6997\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7005\,
            I => \N__6997\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6992\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6992\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6989\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6982\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6982\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6989\,
            I => \N__6978\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6975\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__6987\,
            I => \N__6972\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__6982\,
            I => \N__6967\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6964\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__6978\,
            I => \N__6961\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6975\,
            I => \N__6958\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6951\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6951\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6951\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__6967\,
            I => \DMA_CYCLE\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6964\,
            I => \DMA_CYCLE\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__6961\,
            I => \DMA_CYCLE\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__6958\,
            I => \DMA_CYCLE\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6951\,
            I => \DMA_CYCLE\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__6940\,
            I => \U712_BYTE_ENABLE.N_315_cascade_\
        );

    \I__1322\ : IoInMux
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6934\,
            I => \N__6931\
        );

    \I__1320\ : IoSpan4Mux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1318\ : Span12Mux_s9_h
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1317\ : Span12Mux_v
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__6919\,
            I => \N_60_i\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__1312\ : Span12Mux_h
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__6904\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6894\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6894\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6891\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6894\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6891\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6883\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6883\,
            I => \N__6878\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6875\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6872\
        );

    \I__1301\ : Span4Mux_h
    port map (
            O => \N__6878\,
            I => \N__6869\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6875\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6872\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__6869\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6858\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6855\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6852\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6855\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__6852\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6838\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__6843\,
            I => \N__6832\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6829\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6826\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6838\,
            I => \N__6823\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6820\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6836\,
            I => \N__6817\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6809\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6809\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6829\,
            I => \N__6806\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6826\,
            I => \N__6803\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__6823\,
            I => \N__6798\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6798\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6791\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6791\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6791\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6788\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6809\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__6806\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__6803\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6798\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6788\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6770\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6767\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6762\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6757\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6757\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6754\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6751\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6748\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__6757\,
            I => \N__6745\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6754\,
            I => \U712_CHIP_RAM.N_198\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6751\,
            I => \U712_CHIP_RAM.N_198\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__6748\,
            I => \U712_CHIP_RAM.N_198\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__6745\,
            I => \U712_CHIP_RAM.N_198\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6731\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6725\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6725\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6731\,
            I => \N__6722\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6719\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6716\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__6722\,
            I => \N__6713\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6710\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__6716\,
            I => \N__6707\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__6713\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__6710\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__6707\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__6700\,
            I => \U712_CHIP_RAM.N_313_cascade_\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__6691\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\
        );

    \I__1239\ : CEMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__6676\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6669\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6666\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6669\,
            I => \N__6663\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6666\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__6663\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6654\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6651\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6654\,
            I => \N__6648\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6651\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__6648\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6637\,
            I => \N__6633\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6630\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__6633\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6630\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__6619\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__6616\,
            I => \N__6610\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6607\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6601\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6598\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6595\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6589\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6601\,
            I => \N__6589\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6598\,
            I => \N__6583\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__6595\,
            I => \N__6583\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6580\
        );

    \I__1204\ : Span4Mux_h
    port map (
            O => \N__6589\,
            I => \N__6577\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6574\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__6583\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6580\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__6577\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6574\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6562\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6553\,
            I => \N__6549\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__6552\,
            I => \N__6545\
        );

    \I__1192\ : Span4Mux_h
    port map (
            O => \N__6549\,
            I => \N__6538\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6535\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6530\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6530\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6525\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6525\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6522\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__6538\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6535\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6525\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__6505\,
            I => \N__6501\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6498\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6501\,
            I => \LATCH_RAM\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6498\,
            I => \LATCH_RAM\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6488\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6484\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6481\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6478\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__6487\,
            I => \N__6475\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6468\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6468\
        );

    \I__1167\ : Span4Mux_h
    port map (
            O => \N__6478\,
            I => \N__6468\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6465\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__6468\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6465\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6457\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__6454\,
            I => \N__6450\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6447\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6447\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6439\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6436\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6433\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6430\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1152\ : ClkMux
    port map (
            O => \N__6427\,
            I => \N__6409\
        );

    \I__1151\ : ClkMux
    port map (
            O => \N__6426\,
            I => \N__6409\
        );

    \I__1150\ : ClkMux
    port map (
            O => \N__6425\,
            I => \N__6409\
        );

    \I__1149\ : ClkMux
    port map (
            O => \N__6424\,
            I => \N__6409\
        );

    \I__1148\ : ClkMux
    port map (
            O => \N__6423\,
            I => \N__6409\
        );

    \I__1147\ : ClkMux
    port map (
            O => \N__6422\,
            I => \N__6409\
        );

    \I__1146\ : GlobalMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1145\ : gio2CtrlBuf
    port map (
            O => \N__6406\,
            I => \C1_c_g\
        );

    \I__1144\ : SRMux
    port map (
            O => \N__6403\,
            I => \N__6400\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__1142\ : Span4Mux_h
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__6394\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__1138\ : Span4Mux_s2_v
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1136\ : Span12Mux_h
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__6376\,
            I => \BANK0_c\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6370\,
            I => \N__6367\
        );

    \I__1132\ : Span12Mux_v
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1131\ : Span12Mux_h
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__6361\,
            I => \A_c_20\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \N__6348\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__6351\,
            I => \N__6345\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6342\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6338\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6342\,
            I => \N__6334\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6331\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6328\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6324\
        );

    \I__1119\ : Sp12to4
    port map (
            O => \N__6334\,
            I => \N__6321\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6316\
        );

    \I__1117\ : Span4Mux_h
    port map (
            O => \N__6328\,
            I => \N__6316\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6313\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1114\ : Odrv12
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__6316\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6313\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6301\,
            I => \U712_CHIP_RAM.N_405\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6287\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6287\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6287\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6281\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6278\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6287\,
            I => \N__6275\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6271\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6265\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6265\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6281\,
            I => \N__6262\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6278\,
            I => \N__6259\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__6275\,
            I => \N__6256\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6253\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6271\,
            I => \N__6250\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6247\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6265\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__6262\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6256\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6253\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__6250\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6247\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \U712_CHIP_RAM.N_405_cascade_\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6225\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6221\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6218\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__6224\,
            I => \N__6211\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6207\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6204\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6201\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6198\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6194\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6191\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6188\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__6210\,
            I => \N__6185\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__6207\,
            I => \N__6178\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__6204\,
            I => \N__6173\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6173\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6198\,
            I => \N__6170\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6167\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6194\,
            I => \N__6160\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6160\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6160\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6155\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6155\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6148\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6148\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6148\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__6178\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__6173\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6167\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1057\ : Odrv4
    port map (
            O => \N__6160\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6155\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6148\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__6133\,
            I => \U712_CHIP_RAM.N_303_cascade_\
        );

    \I__1053\ : CEMux
    port map (
            O => \N__6130\,
            I => \N__6127\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__6124\,
            I => \N__6121\
        );

    \I__1050\ : Span4Mux_h
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6118\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6109\,
            I => \U712_CHIP_RAM.N_136\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6100\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6100\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__1042\ : Span12Mux_v
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1041\ : Span12Mux_h
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1040\ : Odrv12
    port map (
            O => \N__6091\,
            I => \A_c_10\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6085\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6082\,
            I => \bfn_10_8_0_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6075\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6072\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6072\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6067\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6060\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6057\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6060\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6052\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6045\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6042\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6045\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6042\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6037\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__6034\,
            I => \U712_REG_SM.N_209_cascade_\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6028\,
            I => \N__6025\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__6025\,
            I => \U712_REG_SM.LDSn_7_iv_i_0\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6022\,
            I => \U712_REG_SM.N_297_cascade_\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1014\ : Span12Mux_s11_v
    port map (
            O => \N__6013\,
            I => \N__6010\
        );

    \I__1013\ : Span12Mux_h
    port map (
            O => \N__6010\,
            I => \N__6005\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6000\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6000\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__6005\,
            I => \LDSn_c\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6000\,
            I => \LDSn_c\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__5995\,
            I => \U712_REG_SM.N_295_cascade_\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5986\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5986\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5986\,
            I => \U712_REG_SM.N_153\
        );

    \I__1004\ : IoInMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5977\
        );

    \I__1002\ : Span4Mux_s0_v
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__1000\ : Sp12to4
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__999\ : Span12Mux_h
    port map (
            O => \N__5968\,
            I => \N__5963\
        );

    \I__998\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5958\
        );

    \I__997\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5958\
        );

    \I__996\ : Odrv12
    port map (
            O => \N__5963\,
            I => \UDSn_c\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5958\,
            I => \UDSn_c\
        );

    \I__994\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5949\
        );

    \I__993\ : IoInMux
    port map (
            O => \N__5952\,
            I => \N__5946\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5949\,
            I => \N__5943\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5940\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__5943\,
            I => \N__5937\
        );

    \I__989\ : IoSpan4Mux
    port map (
            O => \N__5940\,
            I => \N__5934\
        );

    \I__988\ : Sp12to4
    port map (
            O => \N__5937\,
            I => \N__5931\
        );

    \I__987\ : IoSpan4Mux
    port map (
            O => \N__5934\,
            I => \N__5928\
        );

    \I__986\ : Span12Mux_h
    port map (
            O => \N__5931\,
            I => \N__5925\
        );

    \I__985\ : IoSpan4Mux
    port map (
            O => \N__5928\,
            I => \N__5922\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__5925\,
            I => \C1_c\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__5922\,
            I => \C1_c\
        );

    \I__982\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5911\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__5911\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__979\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5905\,
            I => \N__5902\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__976\ : Sp12to4
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__975\ : Span12Mux_h
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__974\ : Span12Mux_v
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__973\ : Odrv12
    port map (
            O => \N__5890\,
            I => \REGSPACEn_c\
        );

    \I__972\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5884\,
            I => \N__5880\
        );

    \I__970\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__969\ : Span4Mux_v
    port map (
            O => \N__5880\,
            I => \N__5874\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5877\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__5874\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__965\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5859\
        );

    \I__963\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5856\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__5859\,
            I => \N__5853\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5850\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__5853\,
            I => \N__5847\
        );

    \I__959\ : Span4Mux_v
    port map (
            O => \N__5850\,
            I => \N__5844\
        );

    \I__958\ : Sp12to4
    port map (
            O => \N__5847\,
            I => \N__5839\
        );

    \I__957\ : Sp12to4
    port map (
            O => \N__5844\,
            I => \N__5839\
        );

    \I__956\ : Span12Mux_h
    port map (
            O => \N__5839\,
            I => \N__5836\
        );

    \I__955\ : Odrv12
    port map (
            O => \N__5836\,
            I => \TSn_c\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__5833\,
            I => \N__5829\
        );

    \I__953\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5825\
        );

    \I__952\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5822\
        );

    \I__951\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5819\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5825\,
            I => \N__5816\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5822\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5819\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__5816\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__946\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__5803\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__5800\,
            I => \U712_REG_SM.N_229_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5788\
        );

    \I__941\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5788\
        );

    \I__940\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5783\
        );

    \I__939\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5783\
        );

    \I__938\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5780\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5788\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5783\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__934\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5768\
        );

    \I__933\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5765\
        );

    \I__932\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5762\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5768\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5765\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5762\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5749\,
            I => \U712_REG_SM.REG_CPU_CYCLE_e_1\
        );

    \I__925\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5743\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5743\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__923\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U712_REG_SM.N_224\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5734\,
            I => \U712_REG_SM.N_224_cascade_\
        );

    \I__920\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5728\,
            I => \U712_CHIP_RAM.N_234\
        );

    \I__918\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5719\
        );

    \I__917\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5719\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5719\,
            I => \N__5715\
        );

    \I__915\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5712\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__5715\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5712\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0\
        );

    \I__912\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5702\
        );

    \I__911\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5698\
        );

    \I__910\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5695\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5692\
        );

    \I__908\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5688\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5698\,
            I => \N__5684\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5695\,
            I => \N__5681\
        );

    \I__905\ : Span4Mux_h
    port map (
            O => \N__5692\,
            I => \N__5678\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__5691\,
            I => \N__5675\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5671\
        );

    \I__902\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5668\
        );

    \I__901\ : Span4Mux_v
    port map (
            O => \N__5684\,
            I => \N__5661\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__5681\,
            I => \N__5661\
        );

    \I__899\ : Span4Mux_h
    port map (
            O => \N__5678\,
            I => \N__5661\
        );

    \I__898\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5656\
        );

    \I__897\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5656\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__5671\,
            I => \WRITE_CYCLE\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5668\,
            I => \WRITE_CYCLE\
        );

    \I__894\ : Odrv4
    port map (
            O => \N__5661\,
            I => \WRITE_CYCLE\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5656\,
            I => \WRITE_CYCLE\
        );

    \I__892\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5638\
        );

    \I__891\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5635\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__5645\,
            I => \N__5632\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5644\,
            I => \N__5626\
        );

    \I__888\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5622\
        );

    \I__887\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5619\
        );

    \I__886\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5615\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5638\,
            I => \N__5610\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5635\,
            I => \N__5610\
        );

    \I__883\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5607\
        );

    \I__882\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5604\
        );

    \I__881\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5601\
        );

    \I__880\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5596\
        );

    \I__879\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5596\
        );

    \I__878\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5593\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5588\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5619\,
            I => \N__5588\
        );

    \I__875\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5585\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5615\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5610\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5607\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5604\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5601\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5588\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5585\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__865\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5563\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5560\,
            I => \N__5557\
        );

    \I__862\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5554\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5554\,
            I => \U712_CHIP_RAM.N_292\
        );

    \I__860\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.N_19\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__856\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5536\,
            I => \U712_BYTE_ENABLE.N_185_i\
        );

    \I__854\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5530\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_5\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__5527\,
            I => \U712_CHIP_RAM.N_391_cascade_\
        );

    \I__851\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5521\,
            I => \U712_CHIP_RAM.N_387\
        );

    \I__849\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5514\
        );

    \I__848\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5511\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5514\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5511\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5506\,
            I => \N__5502\
        );

    \I__844\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5496\
        );

    \I__843\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5493\
        );

    \I__842\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5488\
        );

    \I__841\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5488\
        );

    \I__840\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5484\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5480\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5493\,
            I => \N__5475\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5488\,
            I => \N__5475\
        );

    \I__836\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5472\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5484\,
            I => \N__5469\
        );

    \I__834\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5466\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5475\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5472\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__5469\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5466\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__828\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__827\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5446\
        );

    \I__826\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5435\
        );

    \I__825\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5435\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5430\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5430\
        );

    \I__822\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5423\
        );

    \I__821\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5423\
        );

    \I__820\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5423\
        );

    \I__819\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5418\
        );

    \I__818\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5418\
        );

    \I__817\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5415\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5435\,
            I => \N__5412\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5418\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5415\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__5412\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__5401\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_\
        );

    \I__809\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5386\
        );

    \I__808\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5386\
        );

    \I__807\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5378\
        );

    \I__806\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5371\
        );

    \I__805\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5371\
        );

    \I__804\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5371\
        );

    \I__803\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5368\
        );

    \I__802\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5365\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5362\
        );

    \I__800\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5355\
        );

    \I__799\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5355\
        );

    \I__798\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5355\
        );

    \I__797\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5350\
        );

    \I__796\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5350\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5378\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5371\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5368\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5355\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__788\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5329\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__5329\,
            I => \N__5325\
        );

    \I__785\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5322\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__5325\,
            I => \N__5317\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5317\
        );

    \I__782\ : Span12Mux_h
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__781\ : Span12Mux_v
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__780\ : Odrv12
    port map (
            O => \N__5311\,
            I => \AWEn_c\
        );

    \I__779\ : IoInMux
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__777\ : Span4Mux_s2_v
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__776\ : Span4Mux_v
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__5296\,
            I => \N__5293\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__5293\,
            I => \N__5289\
        );

    \I__773\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5286\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__5289\,
            I => \DBDIR_c\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5286\,
            I => \DBDIR_c\
        );

    \I__770\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5278\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__768\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5269\
        );

    \I__767\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5269\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5269\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0\
        );

    \I__765\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__763\ : Span4Mux_h
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__5257\,
            I => \U712_CHIP_RAM.N_399\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \U712_CHIP_RAM.N_399_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__5242\,
            I => \U712_CHIP_RAM.N_277\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__5239\,
            I => \U712_CHIP_RAM.N_277_cascade_\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__5236\,
            I => \U712_CHIP_RAM.N_347_cascade_\
        );

    \I__754\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5229\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__5232\,
            I => \N__5226\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5229\,
            I => \N__5221\
        );

    \I__751\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5218\
        );

    \I__750\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5215\
        );

    \I__749\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5212\
        );

    \I__748\ : Span4Mux_h
    port map (
            O => \N__5221\,
            I => \N__5209\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5218\,
            I => \U712_CHIP_RAM.N_353\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5215\,
            I => \U712_CHIP_RAM.N_353\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5212\,
            I => \U712_CHIP_RAM.N_353\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__5209\,
            I => \U712_CHIP_RAM.N_353\
        );

    \I__743\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5192\
        );

    \I__741\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5188\
        );

    \I__740\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5185\
        );

    \I__739\ : Span4Mux_h
    port map (
            O => \N__5192\,
            I => \N__5182\
        );

    \I__738\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5179\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5188\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__5182\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5179\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__5170\,
            I => \N__5164\
        );

    \I__732\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5161\
        );

    \I__731\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5158\
        );

    \I__730\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5155\
        );

    \I__729\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5152\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5161\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5143\,
            I => \N__5138\
        );

    \I__723\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5134\
        );

    \I__722\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5131\
        );

    \I__721\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5128\
        );

    \I__720\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5125\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5134\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5131\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5128\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5125\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__715\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__714\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5110\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5106\
        );

    \I__712\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5103\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__5106\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5103\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__5098\,
            I => \U712_CHIP_RAM.N_343_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5083\
        );

    \I__707\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5083\
        );

    \I__706\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5083\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5080\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__5091\,
            I => \N__5077\
        );

    \I__703\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5071\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5068\
        );

    \I__701\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5065\
        );

    \I__700\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5062\
        );

    \I__699\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5059\
        );

    \I__698\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5054\
        );

    \I__697\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5054\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__5068\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5065\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__690\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5031\
        );

    \I__689\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5028\
        );

    \I__688\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5025\
        );

    \I__687\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5022\
        );

    \I__686\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5019\
        );

    \I__685\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5014\
        );

    \I__684\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5014\
        );

    \I__683\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5011\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5022\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5019\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5011\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__675\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4991\
        );

    \I__674\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4988\
        );

    \I__673\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4985\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4981\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4978\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4985\,
            I => \N__4975\
        );

    \I__669\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4972\
        );

    \I__668\ : Span4Mux_h
    port map (
            O => \N__4981\,
            I => \N__4969\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__4978\,
            I => \U712_CHIP_RAM.N_391\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__4975\,
            I => \U712_CHIP_RAM.N_391\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4972\,
            I => \U712_CHIP_RAM.N_391\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__4969\,
            I => \U712_CHIP_RAM.N_391\
        );

    \I__663\ : IoInMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__661\ : IoSpan4Mux
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__660\ : Span4Mux_s0_h
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__659\ : Span4Mux_h
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__657\ : Span12Mux_v
    port map (
            O => \N__4942\,
            I => \N__4938\
        );

    \I__656\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__655\ : Span12Mux_h
    port map (
            O => \N__4938\,
            I => \N__4932\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4929\
        );

    \I__653\ : Span12Mux_h
    port map (
            O => \N__4932\,
            I => \N__4926\
        );

    \I__652\ : Span12Mux_h
    port map (
            O => \N__4929\,
            I => \N__4923\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__4926\,
            I => \C3_c\
        );

    \I__650\ : Odrv12
    port map (
            O => \N__4923\,
            I => \C3_c\
        );

    \I__649\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4915\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__4906\,
            I => \A_c_9\
        );

    \I__644\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4900\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__641\ : Sp12to4
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__640\ : Span12Mux_h
    port map (
            O => \N__4891\,
            I => \N__4888\
        );

    \I__639\ : Span12Mux_v
    port map (
            O => \N__4888\,
            I => \N__4885\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__4885\,
            I => \A_c_2\
        );

    \I__637\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4879\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__4876\,
            I => \N__4873\
        );

    \I__634\ : Sp12to4
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__633\ : Span12Mux_h
    port map (
            O => \N__4870\,
            I => \N__4867\
        );

    \I__632\ : Odrv12
    port map (
            O => \N__4867\,
            I => \A_c_12\
        );

    \I__631\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4861\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4861\,
            I => \N__4858\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__4858\,
            I => \N__4855\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__4855\,
            I => \N__4852\
        );

    \I__627\ : Sp12to4
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__626\ : Odrv12
    port map (
            O => \N__4849\,
            I => \A_c_5\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__624\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__621\ : Span12Mux_v
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__4831\,
            I => \A_c_3\
        );

    \I__619\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4825\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4825\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\
        );

    \I__617\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__615\ : Span4Mux_h
    port map (
            O => \N__4816\,
            I => \N__4813\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__613\ : Span4Mux_v
    port map (
            O => \N__4810\,
            I => \N__4807\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__4804\,
            I => \RAMSPACEn_c\
        );

    \I__610\ : IoInMux
    port map (
            O => \N__4801\,
            I => \N__4797\
        );

    \I__609\ : IoInMux
    port map (
            O => \N__4800\,
            I => \N__4794\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4791\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4788\
        );

    \I__606\ : Span12Mux_s3_h
    port map (
            O => \N__4791\,
            I => \N__4785\
        );

    \I__605\ : Span4Mux_s3_v
    port map (
            O => \N__4788\,
            I => \N__4782\
        );

    \I__604\ : Span12Mux_v
    port map (
            O => \N__4785\,
            I => \N__4779\
        );

    \I__603\ : Span4Mux_h
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__602\ : Span12Mux_h
    port map (
            O => \N__4779\,
            I => \N__4773\
        );

    \I__601\ : Sp12to4
    port map (
            O => \N__4776\,
            I => \N__4770\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__4773\,
            I => \N_246\
        );

    \I__599\ : Odrv12
    port map (
            O => \N__4770\,
            I => \N_246\
        );

    \I__598\ : IoInMux
    port map (
            O => \N__4765\,
            I => \N__4762\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__596\ : IoSpan4Mux
    port map (
            O => \N__4759\,
            I => \N__4756\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__594\ : Span12Mux_v
    port map (
            O => \N__4753\,
            I => \N__4749\
        );

    \I__593\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__4749\,
            I => \REGENn_c\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4746\,
            I => \REGENn_c\
        );

    \I__590\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4737\
        );

    \I__589\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4734\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4737\,
            I => \LATCH_REG\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4734\,
            I => \LATCH_REG\
        );

    \I__586\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4726\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__584\ : Span12Mux_v
    port map (
            O => \N__4723\,
            I => \N__4719\
        );

    \I__583\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4716\
        );

    \I__582\ : Odrv12
    port map (
            O => \N__4719\,
            I => \REG_CPU_CYCLE\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4716\,
            I => \REG_CPU_CYCLE\
        );

    \I__580\ : IoInMux
    port map (
            O => \N__4711\,
            I => \N__4708\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4708\,
            I => \N__4705\
        );

    \I__578\ : Span4Mux_s3_v
    port map (
            O => \N__4705\,
            I => \N__4702\
        );

    \I__577\ : Span4Mux_h
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__576\ : Sp12to4
    port map (
            O => \N__4699\,
            I => \N__4696\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__4696\,
            I => \N__4692\
        );

    \I__574\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4689\
        );

    \I__573\ : Odrv12
    port map (
            O => \N__4692\,
            I => \ASn_c\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4689\,
            I => \ASn_c\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__4684\,
            I => \U712_CHIP_RAM.N_400_cascade_\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__569\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4674\
        );

    \I__568\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4671\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4666\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4666\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__4663\,
            I => \U712_CHIP_RAM.N_266\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__4660\,
            I => \U712_CHIP_RAM.N_304_cascade_\
        );

    \I__562\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4654\,
            I => \U712_CHIP_RAM.N_249\
        );

    \I__560\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4646\
        );

    \I__559\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4643\
        );

    \I__558\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4639\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4646\,
            I => \N__4636\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4643\,
            I => \N__4633\
        );

    \I__555\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4630\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4639\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__4636\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4633\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__550\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4617\
        );

    \I__549\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4614\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4610\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4607\
        );

    \I__546\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4604\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__4610\,
            I => \U712_CHIP_RAM.N_350_0\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__4607\,
            I => \U712_CHIP_RAM.N_350_0\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4604\,
            I => \U712_CHIP_RAM.N_350_0\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4597\,
            I => \U712_CHIP_RAM.N_291_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4591\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0\
        );

    \I__539\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\
        );

    \I__537\ : InMux
    port map (
            O => \N__4582\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__536\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__534\ : InMux
    port map (
            O => \N__4573\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__533\ : InMux
    port map (
            O => \N__4570\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__532\ : InMux
    port map (
            O => \N__4567\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__531\ : InMux
    port map (
            O => \N__4564\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__530\ : InMux
    port map (
            O => \N__4561\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__529\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4551\
        );

    \I__528\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4551\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__4556\,
            I => \N__4543\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4540\
        );

    \I__525\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4533\
        );

    \I__524\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4533\
        );

    \I__523\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4533\
        );

    \I__522\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4526\
        );

    \I__521\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4526\
        );

    \I__520\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4526\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__4540\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4533\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4526\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__516\ : InMux
    port map (
            O => \N__4519\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__515\ : CEMux
    port map (
            O => \N__4516\,
            I => \N__4512\
        );

    \I__514\ : CEMux
    port map (
            O => \N__4515\,
            I => \N__4509\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4512\,
            I => \N__4506\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4509\,
            I => \N__4503\
        );

    \I__511\ : Span4Mux_v
    port map (
            O => \N__4506\,
            I => \N__4500\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__4503\,
            I => \N__4497\
        );

    \I__509\ : Span4Mux_h
    port map (
            O => \N__4500\,
            I => \N__4494\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__4497\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4494\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__506\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4481\
        );

    \I__505\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4481\
        );

    \I__504\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4476\
        );

    \I__503\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4476\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4481\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4476\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__4471\,
            I => \N__4467\
        );

    \I__499\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4460\
        );

    \I__498\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4460\
        );

    \I__497\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4455\
        );

    \I__496\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4455\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4460\,
            I => \U712_CHIP_RAM.N_280\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4455\,
            I => \U712_CHIP_RAM.N_280\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4450\,
            I => \U712_CHIP_RAM.N_301_cascade_\
        );

    \I__492\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4443\
        );

    \I__491\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4440\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4443\,
            I => \U712_CHIP_RAM.N_280_2\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4440\,
            I => \U712_CHIP_RAM.N_280_2\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__487\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4429\,
            I => \U712_CHIP_RAM.N_192\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__4426\,
            I => \U712_CHIP_RAM.N_192_cascade_\
        );

    \I__484\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4420\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4420\,
            I => \U712_CHIP_RAM.N_215\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__4417\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_\
        );

    \I__481\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4411\,
            I => \U712_CHIP_RAM.N_345\
        );

    \I__479\ : IoInMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__477\ : IoSpan4Mux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__476\ : Span4Mux_s2_v
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__475\ : Sp12to4
    port map (
            O => \N__4396\,
            I => \N__4393\
        );

    \I__474\ : Odrv12
    port map (
            O => \N__4393\,
            I => \LATCH_CLK_0_i\
        );

    \I__473\ : IoInMux
    port map (
            O => \N__4390\,
            I => \N__4386\
        );

    \I__472\ : IoInMux
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4377\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4383\,
            I => \N__4377\
        );

    \I__469\ : IoInMux
    port map (
            O => \N__4382\,
            I => \N__4374\
        );

    \I__468\ : IoSpan4Mux
    port map (
            O => \N__4377\,
            I => \N__4371\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4368\
        );

    \I__466\ : Sp12to4
    port map (
            O => \N__4371\,
            I => \N__4365\
        );

    \I__465\ : Span4Mux_s3_h
    port map (
            O => \N__4368\,
            I => \N__4362\
        );

    \I__464\ : Span12Mux_v
    port map (
            O => \N__4365\,
            I => \N__4359\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__462\ : Span12Mux_h
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__4356\,
            I => \N__4350\
        );

    \I__460\ : Odrv12
    port map (
            O => \N__4353\,
            I => \CLK40_PLL_iso_i\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__4350\,
            I => \CLK40_PLL_iso_i\
        );

    \I__458\ : IoInMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__456\ : Span12Mux_s5_v
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4336\,
            I => \VBENn_c\
        );

    \I__454\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__452\ : Span12Mux_h
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__4324\,
            I => \A_c_11\
        );

    \I__450\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__448\ : Span4Mux_h
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__447\ : Sp12to4
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__4309\,
            I => \N__4306\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__4306\,
            I => \A_c_4\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4303\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\
        );

    \I__443\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4297\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__441\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4291\,
            I => \U712_CHIP_RAM.N_283\
        );

    \I__439\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4284\
        );

    \I__438\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4284\,
            I => \N__4276\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N__4276\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__4276\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0\
        );

    \I__434\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4268\
        );

    \I__433\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4263\
        );

    \I__432\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4263\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4268\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4263\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \U712_CHIP_RAM.N_389_cascade_\
        );

    \I__428\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4252\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4249\,
            I => \U712_CHIP_RAM.N_348_cascade_\
        );

    \I__425\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4243\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0\
        );

    \I__423\ : IoInMux
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__421\ : IoSpan4Mux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__419\ : Span12Mux_s9_h
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__418\ : Span12Mux_h
    port map (
            O => \N__4225\,
            I => \N__4221\
        );

    \I__417\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__4221\,
            I => \CLK_EN_c\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__4218\,
            I => \CLK_EN_c\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__4213\,
            I => \DBRn_c_i_cascade_\
        );

    \I__413\ : IoInMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__411\ : Span12Mux_s5_h
    port map (
            O => \N__4204\,
            I => \N__4201\
        );

    \I__410\ : Odrv12
    port map (
            O => \N__4201\,
            I => \DBRn_c_i_0\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__4198\,
            I => \U712_CHIP_RAM.N_288_cascade_\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__4195\,
            I => \U712_CHIP_RAM.N_325_cascade_\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__4192\,
            I => \U712_CHIP_RAM.N_308_cascade_\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4189\,
            I => \U712_CHIP_RAM.N_350_0_cascade_\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__4186\,
            I => \U712_CHIP_RAM.N_355_cascade_\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__402\ : Span4Mux_s2_v
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__400\ : Span4Mux_h
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__4168\,
            I => \CLK80_PLL_i_i\
        );

    \I__398\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__393\ : Odrv12
    port map (
            O => \N__4150\,
            I => \A_c_14\
        );

    \I__392\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__388\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__387\ : Odrv12
    port map (
            O => \N__4132\,
            I => \A_c_7\
        );

    \I__386\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__384\ : Span4Mux_v
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__383\ : Span4Mux_v
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__382\ : Sp12to4
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__4114\,
            I => \A_c_16\
        );

    \I__380\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__4096\,
            I => \A_c_18\
        );

    \I__374\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__372\ : Sp12to4
    port map (
            O => \N__4087\,
            I => \N__4084\
        );

    \I__371\ : Span12Mux_v
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__4081\,
            I => \A_c_15\
        );

    \I__369\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__4075\,
            I => \N__4072\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__4069\,
            I => \N__4066\
        );

    \I__365\ : Sp12to4
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__4063\,
            I => \A_c_8\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__4060\,
            I => \U712_CHIP_RAM.N_350_cascade_\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__4057\,
            I => \U712_CHIP_RAM.N_376_cascade_\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__4054\,
            I => \U712_CHIP_RAM.N_280_cascade_\
        );

    \I__360\ : IoInMux
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__4048\,
            I => \N__4045\
        );

    \I__358\ : Span4Mux_s0_v
    port map (
            O => \N__4045\,
            I => \N__4042\
        );

    \I__357\ : Span4Mux_v
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__356\ : Sp12to4
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__355\ : Span12Mux_h
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__354\ : Span12Mux_v
    port map (
            O => \N__4033\,
            I => \N__4030\
        );

    \I__353\ : Odrv12
    port map (
            O => \N__4030\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__6422\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__6423\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__6424\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__6426\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__6425\
        );

    \INVU712_REG_SM.DBR_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.DBR_SYNC_0C_net\,
            I => \N__9081\
        );

    \INVU712_REG_SM.REG_TACKC\ : INV
    port map (
            O => \INVU712_REG_SM.REG_TACKC_net\,
            I => \N__9077\
        );

    \INVU712_REG_SM.C1_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.C1_SYNC_0C_net\,
            I => \N__9086\
        );

    \INVU712_REG_SM.C3_SYNC_1C\ : INV
    port map (
            O => \INVU712_REG_SM.C3_SYNC_1C_net\,
            I => \N__9080\
        );

    \INVU712_REG_SM.STATE_COUNTER_0C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_0C_net\,
            I => \N__9078\
        );

    \INVU712_REG_SM.CYCLE_RUNC\ : INV
    port map (
            O => \INVU712_REG_SM.CYCLE_RUNC_net\,
            I => \N__9076\
        );

    \INVU712_REG_SM.ASnC\ : INV
    port map (
            O => \INVU712_REG_SM.ASnC_net\,
            I => \N__9085\
        );

    \INVU712_REG_SM.REGENnC\ : INV
    port map (
            O => \INVU712_REG_SM.REGENnC_net\,
            I => \N__9079\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \CLK40_PLL_derived_clock_RNIIOT\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8454\,
            GLOBALBUFFEROUTPUT => \CLK40_PLL_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8770\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5952\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4210\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4960\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10393\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4165\,
            in1 => \N__4147\,
            in2 => \_gnd_net_\,
            in3 => \N__9237\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9238\,
            in1 => \N__4129\,
            in2 => \_gnd_net_\,
            in3 => \N__4111\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9239\,
            in1 => \N__4093\,
            in2 => \_gnd_net_\,
            in3 => \N__4078\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILSBFD_4_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__5094\,
            in1 => \N__5233\,
            in2 => \N__9003\,
            in3 => \N__4423\,
            lcout => \U712_CHIP_RAM.N_350\,
            ltout => \U712_CHIP_RAM.N_350_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4060\,
            in3 => \N__4271\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__4465\,
            in1 => \N__4489\,
            in2 => \N__4057\,
            in3 => \N__8541\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__6493\,
            in1 => \N__6613\,
            in2 => \N__6352\,
            in3 => \N__4446\,
            lcout => \U712_CHIP_RAM.N_280\,
            ltout => \U712_CHIP_RAM.N_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1RLTB_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5093\,
            in1 => \N__4677\,
            in2 => \N__4054\,
            in3 => \N__4287\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__8995\,
            in2 => \N__4435\,
            in3 => \N__5095\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4272\,
            in1 => \N__6614\,
            in2 => \N__4198\,
            in3 => \N__4447\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__4488\,
            in1 => \N__4466\,
            in2 => \N__4195\,
            in3 => \N__9245\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISJJB2_7_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5452\,
            in2 => \_gnd_net_\,
            in3 => \N__8992\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVENA4_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5453\,
            in1 => \N__5382\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILAVHF_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4255\,
            in1 => \N__8993\,
            in2 => \N__4192\,
            in3 => \N__6837\,
            lcout => \U712_CHIP_RAM.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7BNR1_7_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5191\,
            in1 => \N__5137\,
            in2 => \N__5170\,
            in3 => \N__5381\,
            lcout => \U712_CHIP_RAM.N_350_0\,
            ltout => \U712_CHIP_RAM.N_350_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5631\,
            in2 => \N__4189\,
            in3 => \N__6543\,
            lcout => \U712_CHIP_RAM.N_355\,
            ltout => \U712_CHIP_RAM.N_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__8991\,
            in1 => \_gnd_net_\,
            in2 => \N__4186\,
            in3 => \N__6881\,
            lcout => \U712_CHIP_RAM.N_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4613\,
            in1 => \N__5483\,
            in2 => \_gnd_net_\,
            in3 => \N__6542\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => \U712_CHIP_RAM.N_389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__5707\,
            in1 => \N__4996\,
            in2 => \N__4258\,
            in3 => \N__4642\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6181\,
            in1 => \N__5074\,
            in2 => \_gnd_net_\,
            in3 => \N__5035\,
            lcout => \U712_CHIP_RAM.N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__6183\,
            in1 => \N__4995\,
            in2 => \_gnd_net_\,
            in3 => \N__4649\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10382\,
            ce => 'H',
            sr => \N__10645\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6182\,
            lcout => \U712_CHIP_RAM.N_348\,
            ltout => \U712_CHIP_RAM.N_348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRD202_3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__6988\,
            in1 => \N__5036\,
            in2 => \N__4249\,
            in3 => \N__5646\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__7022\,
            in1 => \N__5517\,
            in2 => \N__6847\,
            in3 => \N__9628\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10386\,
            ce => 'H',
            sr => \N__10640\
        );

    \U712_CHIP_RAM.CLK_EN_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__5266\,
            in1 => \N__4224\,
            in2 => \N__5506\,
            in3 => \N__5251\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10386\,
            ce => 'H',
            sr => \N__10640\
        );

    \DBRn_ibuf_RNIBAB_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => \DBRn_c_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4213\,
            in3 => \N__10663\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.LATCH_CLK_0_i_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6511\,
            lcout => \LATCH_CLK_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9094\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9450\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__4321\,
            in2 => \_gnd_net_\,
            in3 => \N__9236\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4294\,
            in1 => \N__4621\,
            in2 => \N__9004\,
            in3 => \N__5505\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4994\,
            in1 => \N__8999\,
            in2 => \N__4303\,
            in3 => \N__4651\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__4300\,
            in1 => \N__4487\,
            in2 => \N__4471\,
            in3 => \N__8606\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__4594\,
            in2 => \_gnd_net_\,
            in3 => \N__5443\,
            lcout => \U712_CHIP_RAM.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__4288\,
            in1 => \N__4273\,
            in2 => \N__4681\,
            in3 => \N__5706\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__4470\,
            in2 => \N__4450\,
            in3 => \N__8497\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10372\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__8994\,
            in2 => \N__6224\,
            in3 => \N__6814\,
            lcout => \U712_CHIP_RAM.N_280_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__5394\,
            in1 => \N__5444\,
            in2 => \N__5645\,
            in3 => \N__4414\,
            lcout => \U712_CHIP_RAM.N_192\,
            ltout => \U712_CHIP_RAM.N_192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__5445\,
            in1 => \N__6214\,
            in2 => \N__4426\,
            in3 => \N__5395\,
            lcout => \U712_CHIP_RAM.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__4546\,
            in1 => \N__8703\,
            in2 => \N__6552\,
            in3 => \N__4828\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10375\,
            ce => \N__4516\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__5391\,
            in2 => \N__5644\,
            in3 => \N__6544\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__5195\,
            in2 => \N__4417\,
            in3 => \N__5168\,
            lcout => \U712_CHIP_RAM.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__4588\,
            in2 => \N__5232\,
            in3 => \N__4547\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10375\,
            ce => \N__4516\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__5225\,
            in1 => \N__4579\,
            in2 => \N__4556\,
            in3 => \N__5725\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10375\,
            ce => \N__4516\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_4_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5629\,
            in1 => \N__8977\,
            in2 => \N__5092\,
            in3 => \N__6197\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6548\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5396\,
            in2 => \_gnd_net_\,
            in3 => \N__4582\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5641\,
            in2 => \_gnd_net_\,
            in3 => \N__4573\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__5041\,
            in2 => \_gnd_net_\,
            in3 => \N__4570\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10379\,
            ce => \N__4515\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4557\,
            in1 => \N__5090\,
            in2 => \_gnd_net_\,
            in3 => \N__4567\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10379\,
            ce => \N__4515\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__5169\,
            in2 => \_gnd_net_\,
            in3 => \N__4564\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10379\,
            ce => \N__4515\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4558\,
            in1 => \N__5196\,
            in2 => \_gnd_net_\,
            in3 => \N__4561\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10379\,
            ce => \N__4515\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4550\,
            in1 => \N__5142\,
            in2 => \_gnd_net_\,
            in3 => \N__4519\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10379\,
            ce => \N__4515\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPI372_4_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__5115\,
            in2 => \N__5091\,
            in3 => \N__5397\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILMBG3_4_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4684\,
            in3 => \N__5487\,
            lcout => \U712_CHIP_RAM.N_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBO8O5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4657\,
            in1 => \N__5454\,
            in2 => \N__6210\,
            in3 => \N__5398\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => \U712_CHIP_RAM.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI34JU9_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__5687\,
            in1 => \N__6730\,
            in2 => \N__4660\,
            in3 => \N__5643\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIC6723_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6274\,
            in1 => \N__5116\,
            in2 => \_gnd_net_\,
            in3 => \N__5524\,
            lcout => \U712_CHIP_RAM.N_249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6882\,
            in1 => \N__4650\,
            in2 => \_gnd_net_\,
            in3 => \N__5040\,
            lcout => \U712_CHIP_RAM.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101100"
        )
    port map (
            in0 => \N__8936\,
            in1 => \N__6285\,
            in2 => \N__6916\,
            in3 => \N__7002\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6765\,
            in1 => \N__4620\,
            in2 => \_gnd_net_\,
            in3 => \N__5500\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__5501\,
            in1 => \N__5455\,
            in2 => \N__4597\,
            in3 => \N__5647\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMQBQ1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__6861\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__7567\,
            in1 => \N__5328\,
            in2 => \_gnd_net_\,
            in3 => \N__6284\,
            lcout => \U712_CHIP_RAM.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__4822\,
            in1 => \N__9411\,
            in2 => \N__5869\,
            in3 => \N__6337\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10389\,
            ce => 'H',
            sr => \N__10618\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7726\,
            lcout => \U712_BYTE_ENABLE.N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__7599\,
            in1 => \N__8052\,
            in2 => \_gnd_net_\,
            in3 => \N__5701\,
            lcout => \N_246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__4752\,
            in1 => \N__7339\,
            in2 => \_gnd_net_\,
            in3 => \N__5794\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REGENnC_net\,
            ce => 'H',
            sr => \N__10610\
        );

    \U712_REG_SM.LATCH_REG_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__6900\,
            in1 => \N__5795\,
            in2 => \N__7600\,
            in3 => \N__4740\,
            lcout => \LATCH_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REGENnC_net\,
            ce => 'H',
            sr => \N__10610\
        );

    \U712_REG_SM.STATE_COUNTER_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6901\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REGENnC_net\,
            ce => 'H',
            sr => \N__10610\
        );

    \U712_REG_SM.REG_CPU_CYCLE_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000000101"
        )
    port map (
            in0 => \N__5772\,
            in1 => \N__4722\,
            in2 => \N__7477\,
            in3 => \N__5752\,
            lcout => \REG_CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REGENnC_net\,
            ce => 'H',
            sr => \N__10610\
        );

    \U712_REG_SM.ASn_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__5797\,
            in1 => \N__5740\,
            in2 => \N__7297\,
            in3 => \N__4695\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.ASnC_net\,
            ce => 'H',
            sr => \N__10608\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4941\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.ASnC_net\,
            ce => 'H',
            sr => \N__10608\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__5796\,
            in1 => \N__8045\,
            in2 => \_gnd_net_\,
            in3 => \N__7180\,
            lcout => \REG_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.ASnC_net\,
            ce => 'H',
            sr => \N__10608\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4918\,
            in1 => \N__4903\,
            in2 => \_gnd_net_\,
            in3 => \N__9248\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8600\,
            in2 => \_gnd_net_\,
            in3 => \N__8492\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8493\,
            in1 => \N__8611\,
            in2 => \_gnd_net_\,
            in3 => \N__9249\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9250\,
            in1 => \N__4882\,
            in2 => \_gnd_net_\,
            in3 => \N__4864\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9378\,
            in1 => \N__9251\,
            in2 => \N__4846\,
            in3 => \N__9658\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4843\,
            in1 => \N__9377\,
            in2 => \_gnd_net_\,
            in3 => \N__9682\,
            lcout => \U712_CHIP_RAM.N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__5224\,
            in1 => \N__6294\,
            in2 => \N__6229\,
            in3 => \N__6615\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5442\,
            in2 => \_gnd_net_\,
            in3 => \N__5385\,
            lcout => \U712_CHIP_RAM.N_399\,
            ltout => \U712_CHIP_RAM.N_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6773\,
            in1 => \N__9379\,
            in2 => \N__5254\,
            in3 => \N__4984\,
            lcout => \U712_CHIP_RAM.N_277\,
            ltout => \U712_CHIP_RAM.N_277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__9380\,
            in1 => \N__5039\,
            in2 => \N__5239\,
            in3 => \N__5705\,
            lcout => \U712_CHIP_RAM.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5034\,
            in2 => \_gnd_net_\,
            in3 => \N__5618\,
            lcout => \U712_CHIP_RAM.N_347\,
            ltout => \U712_CHIP_RAM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8976\,
            in1 => \N__5441\,
            in2 => \N__5236\,
            in3 => \N__5384\,
            lcout => \U712_CHIP_RAM.N_353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ANR1_7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5200\,
            in1 => \N__5167\,
            in2 => \N__5143\,
            in3 => \N__6541\,
            lcout => \U712_CHIP_RAM.N_343\,
            ltout => \U712_CHIP_RAM.N_343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5109\,
            in2 => \N__5098\,
            in3 => \N__5383\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5076\,
            in2 => \_gnd_net_\,
            in3 => \N__5037\,
            lcout => \U712_CHIP_RAM.N_391\,
            ltout => \U712_CHIP_RAM.N_391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNI0TLK1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6970\,
            in2 => \N__5527\,
            in3 => \N__5625\,
            lcout => \U712_CHIP_RAM.N_387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5274\,
            in1 => \N__6835\,
            in2 => \N__6987\,
            in3 => \N__5518\,
            lcout => \DMA_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10376\,
            ce => 'H',
            sr => \N__10632\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5630\,
            in1 => \N__5499\,
            in2 => \_gnd_net_\,
            in3 => \N__6971\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5440\,
            in2 => \N__5401\,
            in3 => \N__5392\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__5335\,
            in1 => \N__5292\,
            in2 => \N__6843\,
            in3 => \N__5275\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10376\,
            ce => 'H',
            sr => \N__10632\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6341\,
            in1 => \N__6492\,
            in2 => \N__6616\,
            in3 => \N__6842\,
            lcout => \CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10380\,
            ce => \N__6130\,
            sr => \N__10625\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__6766\,
            in1 => \N__6736\,
            in2 => \_gnd_net_\,
            in3 => \N__5281\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6228\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__6270\,
            in1 => \N__6588\,
            in2 => \N__6487\,
            in3 => \N__6327\,
            lcout => \U712_CHIP_RAM.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__5718\,
            in2 => \N__5691\,
            in3 => \N__6841\,
            lcout => \WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10383\,
            ce => 'H',
            sr => \N__10619\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5674\,
            in2 => \_gnd_net_\,
            in3 => \N__5642\,
            lcout => \U712_CHIP_RAM.N_198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__5566\,
            in1 => \N__8841\,
            in2 => \N__5560\,
            in3 => \N__5551\,
            lcout => \CPU_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10383\,
            ce => 'H',
            sr => \N__10619\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__7981\,
            in2 => \N__5542\,
            in3 => \N__7795\,
            lcout => \U712_BYTE_ENABLE.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__7845\,
            in1 => \N__7715\,
            in2 => \_gnd_net_\,
            in3 => \N__9413\,
            lcout => \U712_BYTE_ENABLE.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.CYCLE_RUN_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__7334\,
            in1 => \N__7401\,
            in2 => \N__7384\,
            in3 => \N__5883\,
            lcout => \U712_REG_SM.CYCLE_RUNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.CYCLE_RUNC_net\,
            ce => 'H',
            sr => \N__10611\
        );

    \U712_REG_SM.STATE_COUNTER_5_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.CYCLE_RUNC_net\,
            ce => 'H',
            sr => \N__10611\
        );

    \U712_REG_SM.STATE_COUNTER_6_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5533\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.CYCLE_RUNC_net\,
            ce => 'H',
            sr => \N__10611\
        );

    \U712_REG_SM.STATE_COUNTER_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8083\,
            in1 => \N__7428\,
            in2 => \_gnd_net_\,
            in3 => \N__7219\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.CYCLE_RUNC_net\,
            ce => 'H',
            sr => \N__10611\
        );

    \U712_REG_SM.REG_WRITE_CYCLE_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100010111001100"
        )
    port map (
            in0 => \N__7555\,
            in1 => \N__7595\,
            in2 => \N__7405\,
            in3 => \N__7382\,
            lcout => \REG_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.CYCLE_RUNC_net\,
            ce => 'H',
            sr => \N__10611\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__5832\,
            in1 => \N__7292\,
            in2 => \_gnd_net_\,
            in3 => \N__7254\,
            lcout => \U712_REG_SM.N_229\,
            ltout => \U712_REG_SM.N_229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7376\,
            in2 => \N__5800\,
            in3 => \N__5793\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__10609\
        );

    \U712_REG_SM.LDSn_RNO_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__7467\,
            in1 => \N__7885\,
            in2 => \N__7383\,
            in3 => \N__7562\,
            lcout => \U712_REG_SM.LDSn_7_iv_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5917\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__10609\
        );

    \U712_REG_SM.C3_SYNC_RNIELLV_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7466\,
            in1 => \N__7291\,
            in2 => \_gnd_net_\,
            in3 => \N__7253\,
            lcout => \U712_REG_SM.LATCH_REG_0_sqmuxa\,
            ltout => \U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__7594\,
            in1 => \N__5771\,
            in2 => \N__5755\,
            in3 => \N__7175\,
            lcout => \U712_REG_SM.REG_CPU_CYCLE_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5746\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__10604\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__7377\,
            in1 => \N__5828\,
            in2 => \N__7473\,
            in3 => \N__7252\,
            lcout => \U712_REG_SM.N_224\,
            ltout => \U712_REG_SM.N_224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNI5ITS1_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__7290\,
            in1 => \_gnd_net_\,
            in2 => \N__5734\,
            in3 => \N__7216\,
            lcout => \U712_REG_SM.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7289\,
            in2 => \_gnd_net_\,
            in3 => \N__7251\,
            lcout => \U712_REG_SM.N_209\,
            ltout => \U712_REG_SM.N_209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__7884\,
            in1 => \N__6008\,
            in2 => \N__6034\,
            in3 => \N__7218\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__6009\,
            in1 => \N__6031\,
            in2 => \N__6022\,
            in3 => \N__5992\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__10604\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__5966\,
            in1 => \N__7217\,
            in2 => \N__7429\,
            in3 => \N__7960\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__7513\,
            in1 => \N__5967\,
            in2 => \N__5995\,
            in3 => \N__5991\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__10604\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10602\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110101"
        )
    port map (
            in0 => \N__5908\,
            in1 => \N__5887\,
            in2 => \N__5833\,
            in3 => \N__5862\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10602\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9423\,
            in1 => \N__5809\,
            in2 => \N__9298\,
            in3 => \N__9616\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001110010"
        )
    port map (
            in0 => \N__9808\,
            in1 => \N__9247\,
            in2 => \N__6115\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011111111"
        )
    port map (
            in0 => \N__6106\,
            in1 => \N__9109\,
            in2 => \N__9453\,
            in3 => \N__8285\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__6048\,
            in1 => \N__6078\,
            in2 => \N__6454\,
            in3 => \N__6063\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__6105\,
            in1 => \N__9108\,
            in2 => \N__9454\,
            in3 => \N__8286\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__8607\,
            in2 => \N__8554\,
            in3 => \N__9246\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6088\,
            in2 => \_gnd_net_\,
            in3 => \N__6082\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6079\,
            in2 => \_gnd_net_\,
            in3 => \N__6067\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6064\,
            in2 => \_gnd_net_\,
            in3 => \N__6052\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6049\,
            in2 => \_gnd_net_\,
            in3 => \N__6037\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6453\,
            in2 => \_gnd_net_\,
            in3 => \N__6439\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6657\,
            in2 => \_gnd_net_\,
            in3 => \N__6436\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6672\,
            in2 => \_gnd_net_\,
            in3 => \N__6433\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6636\,
            in2 => \_gnd_net_\,
            in3 => \N__6430\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6427\,
            ce => 'H',
            sr => \N__6403\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__6298\,
            in1 => \N__6358\,
            in2 => \N__6836\,
            in3 => \N__8139\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10373\,
            ce => \N__6688\,
            sr => \N__10626\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6373\,
            in1 => \N__6297\,
            in2 => \N__10993\,
            in3 => \N__6304\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6815\,
            in1 => \N__6594\,
            in2 => \N__6351\,
            in3 => \N__6491\,
            lcout => \U712_CHIP_RAM.N_405\,
            ltout => \U712_CHIP_RAM.N_405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6296\,
            in2 => \N__6232\,
            in3 => \N__6216\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__10662\,
            in1 => \N__6775\,
            in2 => \N__6133\,
            in3 => \N__6735\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6886\,
            in1 => \N__6862\,
            in2 => \_gnd_net_\,
            in3 => \N__6816\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__6734\,
            in2 => \N__6700\,
            in3 => \N__6697\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6691\,
            in3 => \N__10661\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6673\,
            in1 => \N__6658\,
            in2 => \N__6643\,
            in3 => \N__6625\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10377\,
            ce => 'H',
            sr => \N__10620\
        );

    \U712_CHIP_RAM.LATCH_RAM_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__6981\,
            in1 => \N__6565\,
            in2 => \N__6559\,
            in3 => \N__6504\,
            lcout => \LATCH_RAM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10377\,
            ce => 'H',
            sr => \N__10620\
        );

    \DBR_SYNC_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6460\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10381\,
            ce => 'H',
            sr => \N__10614\
        );

    \DBR_SYNC_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10381\,
            ce => 'H',
            sr => \N__10614\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_1_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10459\,
            in1 => \N__7006\,
            in2 => \_gnd_net_\,
            in3 => \N__7046\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_58_i_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__7793\,
            in1 => \N__7099\,
            in2 => \N__7159\,
            in3 => \N__7087\,
            lcout => \N_58_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7722\,
            in1 => \N__9448\,
            in2 => \_gnd_net_\,
            in3 => \N__7982\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_56_i_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__7129\,
            in1 => \N__10509\,
            in2 => \N__7050\,
            in3 => \N__7003\,
            lcout => \N_56_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10458\,
            in1 => \N__7005\,
            in2 => \_gnd_net_\,
            in3 => \N__7045\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_54_i_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__7792\,
            in1 => \N__7098\,
            in2 => \N__7090\,
            in3 => \N__7086\,
            lcout => \N_54_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9449\,
            in1 => \N__7794\,
            in2 => \_gnd_net_\,
            in3 => \N__7983\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_60_i_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__7044\,
            in1 => \N__7004\,
            in2 => \N__6940\,
            in3 => \N__10510\,
            lcout => \N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8353\,
            in2 => \_gnd_net_\,
            in3 => \N__10407\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7491\,
            in1 => \N__7462\,
            in2 => \_gnd_net_\,
            in3 => \N__6899\,
            lcout => \U712_REG_SM.un15_0_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__7490\,
            in1 => \_gnd_net_\,
            in2 => \N__7224\,
            in3 => \N__7593\,
            lcout => \U712_REG_SM.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110000"
        )
    port map (
            in0 => \N__7566\,
            in1 => \N__7987\,
            in2 => \N__7472\,
            in3 => \N__7372\,
            lcout => \U712_REG_SM.UDSn_7_iv_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__7504\,
            in1 => \N__7176\,
            in2 => \N__8806\,
            in3 => \N__7498\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_TACKC_net\,
            ce => 'H',
            sr => \N__10605\
        );

    \U712_REG_SM.STATE_COUNTER_7_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__7471\,
            in1 => \N__7293\,
            in2 => \N__7258\,
            in3 => \N__7492\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_TACKC_net\,
            ce => 'H',
            sr => \N__10605\
        );

    \U712_REG_SM.STATE_COUNTER_2_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__8082\,
            in1 => \N__7427\,
            in2 => \N__7225\,
            in3 => \N__7335\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_TACKC_net\,
            ce => 'H',
            sr => \N__10605\
        );

    \U712_REG_SM.STATE_COUNTER_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7400\,
            in2 => \_gnd_net_\,
            in3 => \N__7381\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_TACKC_net\,
            ce => 'H',
            sr => \N__10605\
        );

    \TACKn_obuft_RNO_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_858_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7288\,
            in1 => \N__7250\,
            in2 => \N__8078\,
            in3 => \N__7223\,
            lcout => \U712_REG_SM.REG_TACK_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8120\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.DBR_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10601\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8089\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.DBR_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10601\
        );

    \U712_BYTE_ENABLE.LLBE_0_0_a2_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7857\,
            in1 => \N__7984\,
            in2 => \_gnd_net_\,
            in3 => \N__7711\,
            lcout => \N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10456\,
            in1 => \N__10502\,
            in2 => \_gnd_net_\,
            in3 => \N__8056\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_118_i_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__7710\,
            in1 => \N__7985\,
            in2 => \N__7858\,
            in3 => \N__7750\,
            lcout => \N_118_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7986\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7779\,
            lcout => \U712_BYTE_ENABLE_UUBE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101110"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__7846\,
            in2 => \N__7790\,
            in3 => \N__7708\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_0_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011101010"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__7847\,
            in2 => \N__7791\,
            in3 => \N__7709\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__7639\,
            in1 => \N__9456\,
            in2 => \N__8299\,
            in3 => \N__8161\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10363\,
            ce => \N__9728\,
            sr => \N__10646\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__8298\,
            in1 => \N__8272\,
            in2 => \N__10063\,
            in3 => \N__9457\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10363\,
            ce => \N__9728\,
            sr => \N__10646\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8212\,
            in1 => \N__8206\,
            in2 => \_gnd_net_\,
            in3 => \N__8239\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10368\,
            ce => \N__9735\,
            sr => \N__10641\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001001010"
        )
    port map (
            in0 => \N__9816\,
            in1 => \N__10302\,
            in2 => \N__9281\,
            in3 => \N__9437\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111011"
        )
    port map (
            in0 => \N__10303\,
            in1 => \N__9262\,
            in2 => \N__9455\,
            in3 => \N__9817\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__8200\,
            in1 => \_gnd_net_\,
            in2 => \N__8194\,
            in3 => \N__8185\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10370\,
            ce => \N__9725\,
            sr => \N__10633\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10137\,
            in1 => \N__10195\,
            in2 => \_gnd_net_\,
            in3 => \N__10992\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10717\,
            ce => \N__10688\,
            sr => \N__10627\
        );

    \U712_CHIP_RAM.DMA_A20_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8152\,
            in1 => \N__10988\,
            in2 => \N__10138\,
            in3 => \N__8140\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10615\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8453\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9045\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10378\,
            ce => 'H',
            sr => \N__10612\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8386\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10378\,
            ce => 'H',
            sr => \N__10612\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__8397\,
            in1 => \N__8370\,
            in2 => \N__8455\,
            in3 => \N__9046\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10378\,
            ce => 'H',
            sr => \N__10612\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8385\,
            in1 => \N__9037\,
            in2 => \N__8863\,
            in3 => \N__8369\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__9039\,
            in1 => \N__8861\,
            in2 => \N__9013\,
            in3 => \N__8800\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10384\,
            ce => 'H',
            sr => \N__10606\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8374\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10384\,
            ce => 'H',
            sr => \N__10606\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10408\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10384\,
            ce => 'H',
            sr => \N__10606\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__9038\,
            in1 => \N__8875\,
            in2 => \N__8347\,
            in3 => \N__8799\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10384\,
            ce => 'H',
            sr => \N__10606\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__8975\,
            in1 => \N__8805\,
            in2 => \N__8862\,
            in3 => \N__8893\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10388\,
            ce => \N__8752\,
            sr => \N__10603\
        );

    \U712_CHIP_RAM.RASn_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8619\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10361\,
            ce => 'H',
            sr => \N__10644\
        );

    \U712_CHIP_RAM.WEn_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8506\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10361\,
            ce => 'H',
            sr => \N__10644\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8565\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10361\,
            ce => 'H',
            sr => \N__10644\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8620\,
            in1 => \N__9296\,
            in2 => \N__8566\,
            in3 => \N__8505\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10362\,
            ce => \N__9727\,
            sr => \N__10639\
        );

    \CONSTANT_ONE_LUT4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9424\,
            in1 => \N__8680\,
            in2 => \N__9301\,
            in3 => \N__9118\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8671\,
            in1 => \N__9253\,
            in2 => \_gnd_net_\,
            in3 => \N__8650\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9255\,
            in1 => \N__9442\,
            in2 => \N__8635\,
            in3 => \N__9637\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9254\,
            in1 => \N__9441\,
            in2 => \N__8632\,
            in3 => \N__9124\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__8618\,
            in1 => \N__9252\,
            in2 => \N__8564\,
            in3 => \N__8504\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10660\,
            in1 => \_gnd_net_\,
            in2 => \N__9127\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9901\,
            in1 => \N__10291\,
            in2 => \_gnd_net_\,
            in3 => \N__10980\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10691\,
            sr => \N__10617\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10048\,
            in1 => \N__10002\,
            in2 => \_gnd_net_\,
            in3 => \N__10981\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10691\,
            sr => \N__10617\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10983\,
            in1 => \N__9889\,
            in2 => \_gnd_net_\,
            in3 => \N__10290\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10715\,
            ce => \N__10689\,
            sr => \N__10613\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__9093\,
            in1 => \N__9036\,
            in2 => \_gnd_net_\,
            in3 => \N__8892\,
            lcout => \U712_CYCLE_TERM.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8949\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8950\,
            in2 => \_gnd_net_\,
            in3 => \N__8891\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_227_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__8874\,
            in1 => \N__8854\,
            in2 => \N__8809\,
            in3 => \N__8804\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_227_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8773\,
            in3 => \N__8763\,
            lcout => \U712_CYCLE_TERM.N_227_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9297\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10364\,
            ce => 'H',
            sr => \N__10647\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9451\,
            in1 => \N__9300\,
            in2 => \N__9583\,
            in3 => \N__9646\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__9839\,
            in1 => \N__9777\,
            in2 => \N__9568\,
            in3 => \N__10729\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10369\,
            ce => \N__9736\,
            sr => \N__10642\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9776\,
            in1 => \N__10201\,
            in2 => \N__9841\,
            in3 => \N__9544\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10369\,
            ce => \N__9736\,
            sr => \N__10642\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9299\,
            in1 => \N__9517\,
            in2 => \N__9670\,
            in3 => \N__9452\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__9778\,
            in1 => \N__10147\,
            in2 => \N__9505\,
            in3 => \N__9840\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10369\,
            ce => \N__9736\,
            sr => \N__10642\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__9774\,
            in1 => \N__9838\,
            in2 => \N__10246\,
            in3 => \N__9481\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10371\,
            ce => \N__9726\,
            sr => \N__10634\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9430\,
            in2 => \_gnd_net_\,
            in3 => \N__9261\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__9847\,
            in1 => \N__9837\,
            in2 => \N__9157\,
            in3 => \N__9154\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10371\,
            ce => \N__9726\,
            sr => \N__10634\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__9836\,
            in1 => \N__9787\,
            in2 => \N__9946\,
            in3 => \N__9775\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10371\,
            ce => \N__9726\,
            sr => \N__10634\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10984\,
            in1 => \N__10289\,
            in2 => \_gnd_net_\,
            in3 => \N__10047\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10693\,
            sr => \N__10628\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__10136\,
            in2 => \_gnd_net_\,
            in3 => \N__10194\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10693\,
            sr => \N__10628\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10237\,
            in1 => \N__10001\,
            in2 => \_gnd_net_\,
            in3 => \N__10985\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10693\,
            sr => \N__10628\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10193\,
            in1 => \N__10777\,
            in2 => \_gnd_net_\,
            in3 => \N__10986\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10693\,
            sr => \N__10628\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10828\,
            in1 => \N__10233\,
            in2 => \_gnd_net_\,
            in3 => \N__10982\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10692\,
            sr => \N__10621\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9893\,
            in1 => \N__10954\,
            in2 => \_gnd_net_\,
            in3 => \N__9930\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10690\,
            sr => \N__10616\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__10970\,
            in1 => \N__10822\,
            in2 => \N__10765\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10690\,
            sr => \N__10616\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10457\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10385\,
            ce => 'H',
            sr => \N__10607\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10827\,
            in1 => \N__10232\,
            in2 => \_gnd_net_\,
            in3 => \N__10926\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10716\,
            ce => \N__10695\,
            sr => \N__10643\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10924\,
            in1 => \N__10034\,
            in2 => \_gnd_net_\,
            in3 => \N__10279\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10716\,
            ce => \N__10695\,
            sr => \N__10643\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10003\,
            in1 => \N__10231\,
            in2 => \_gnd_net_\,
            in3 => \N__10925\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10716\,
            ce => \N__10695\,
            sr => \N__10643\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10927\,
            in1 => \N__10776\,
            in2 => \_gnd_net_\,
            in3 => \N__10189\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10716\,
            ce => \N__10695\,
            sr => \N__10643\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10922\,
            in1 => \N__10120\,
            in2 => \_gnd_net_\,
            in3 => \N__10075\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10713\,
            ce => \N__10694\,
            sr => \N__10635\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10033\,
            in1 => \N__9997\,
            in2 => \_gnd_net_\,
            in3 => \N__10921\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10713\,
            ce => \N__10694\,
            sr => \N__10635\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9937\,
            in1 => \N__9900\,
            in2 => \_gnd_net_\,
            in3 => \N__10920\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10713\,
            ce => \N__10694\,
            sr => \N__10635\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10923\,
            in1 => \N__10826\,
            in2 => \_gnd_net_\,
            in3 => \N__10775\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10714\,
            ce => \N__10696\,
            sr => \N__10648\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 4 2025 21:50:11

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_LL_AMIGA,
    D_LM_AMIGA,
    D_UU_AMIGA,
    D_UM_AMIGA,
    D_LL_040,
    D_UU_040,
    D_UM_040,
    D_LM_040,
    A_AMIGA,
    A_040,
    SIZ,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LL_040;
    inout [7:0] D_UU_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LM_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    output CLK40B;
    output TBI_CPUn;
    output TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    input TACKn;
    input BGn;

    wire N__8315;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8290;
    wire N__8289;
    wire N__8288;
    wire N__8281;
    wire N__8280;
    wire N__8279;
    wire N__8272;
    wire N__8271;
    wire N__8270;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8254;
    wire N__8253;
    wire N__8252;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8218;
    wire N__8217;
    wire N__8216;
    wire N__8209;
    wire N__8208;
    wire N__8207;
    wire N__8200;
    wire N__8199;
    wire N__8198;
    wire N__8191;
    wire N__8190;
    wire N__8189;
    wire N__8182;
    wire N__8181;
    wire N__8180;
    wire N__8173;
    wire N__8172;
    wire N__8171;
    wire N__8164;
    wire N__8163;
    wire N__8162;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8146;
    wire N__8145;
    wire N__8144;
    wire N__8137;
    wire N__8136;
    wire N__8135;
    wire N__8128;
    wire N__8127;
    wire N__8126;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8110;
    wire N__8109;
    wire N__8108;
    wire N__8101;
    wire N__8100;
    wire N__8099;
    wire N__8092;
    wire N__8091;
    wire N__8090;
    wire N__8083;
    wire N__8082;
    wire N__8081;
    wire N__8074;
    wire N__8073;
    wire N__8072;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8056;
    wire N__8055;
    wire N__8054;
    wire N__8047;
    wire N__8046;
    wire N__8045;
    wire N__8038;
    wire N__8037;
    wire N__8036;
    wire N__8029;
    wire N__8028;
    wire N__8027;
    wire N__8020;
    wire N__8019;
    wire N__8018;
    wire N__8011;
    wire N__8010;
    wire N__8009;
    wire N__8002;
    wire N__8001;
    wire N__8000;
    wire N__7993;
    wire N__7992;
    wire N__7991;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7975;
    wire N__7974;
    wire N__7973;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7957;
    wire N__7956;
    wire N__7955;
    wire N__7948;
    wire N__7947;
    wire N__7946;
    wire N__7939;
    wire N__7938;
    wire N__7937;
    wire N__7930;
    wire N__7929;
    wire N__7928;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7912;
    wire N__7911;
    wire N__7910;
    wire N__7903;
    wire N__7902;
    wire N__7901;
    wire N__7894;
    wire N__7893;
    wire N__7892;
    wire N__7885;
    wire N__7884;
    wire N__7883;
    wire N__7876;
    wire N__7875;
    wire N__7874;
    wire N__7867;
    wire N__7866;
    wire N__7865;
    wire N__7858;
    wire N__7857;
    wire N__7856;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7840;
    wire N__7839;
    wire N__7838;
    wire N__7831;
    wire N__7830;
    wire N__7829;
    wire N__7822;
    wire N__7821;
    wire N__7820;
    wire N__7813;
    wire N__7812;
    wire N__7811;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7795;
    wire N__7794;
    wire N__7793;
    wire N__7786;
    wire N__7785;
    wire N__7784;
    wire N__7777;
    wire N__7776;
    wire N__7775;
    wire N__7768;
    wire N__7767;
    wire N__7766;
    wire N__7759;
    wire N__7758;
    wire N__7757;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7741;
    wire N__7740;
    wire N__7739;
    wire N__7732;
    wire N__7731;
    wire N__7730;
    wire N__7723;
    wire N__7722;
    wire N__7721;
    wire N__7714;
    wire N__7713;
    wire N__7712;
    wire N__7705;
    wire N__7704;
    wire N__7703;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7687;
    wire N__7686;
    wire N__7685;
    wire N__7678;
    wire N__7677;
    wire N__7676;
    wire N__7669;
    wire N__7668;
    wire N__7667;
    wire N__7660;
    wire N__7659;
    wire N__7658;
    wire N__7651;
    wire N__7650;
    wire N__7649;
    wire N__7642;
    wire N__7641;
    wire N__7640;
    wire N__7633;
    wire N__7632;
    wire N__7631;
    wire N__7624;
    wire N__7623;
    wire N__7622;
    wire N__7615;
    wire N__7614;
    wire N__7613;
    wire N__7606;
    wire N__7605;
    wire N__7604;
    wire N__7597;
    wire N__7596;
    wire N__7595;
    wire N__7588;
    wire N__7587;
    wire N__7586;
    wire N__7579;
    wire N__7578;
    wire N__7577;
    wire N__7570;
    wire N__7569;
    wire N__7568;
    wire N__7561;
    wire N__7560;
    wire N__7559;
    wire N__7552;
    wire N__7551;
    wire N__7550;
    wire N__7543;
    wire N__7542;
    wire N__7541;
    wire N__7534;
    wire N__7533;
    wire N__7532;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7516;
    wire N__7515;
    wire N__7514;
    wire N__7507;
    wire N__7506;
    wire N__7505;
    wire N__7498;
    wire N__7497;
    wire N__7496;
    wire N__7479;
    wire N__7478;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7470;
    wire N__7469;
    wire N__7468;
    wire N__7467;
    wire N__7466;
    wire N__7465;
    wire N__7464;
    wire N__7463;
    wire N__7462;
    wire N__7461;
    wire N__7460;
    wire N__7457;
    wire N__7450;
    wire N__7445;
    wire N__7440;
    wire N__7435;
    wire N__7430;
    wire N__7427;
    wire N__7426;
    wire N__7425;
    wire N__7424;
    wire N__7423;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7411;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7384;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7368;
    wire N__7365;
    wire N__7360;
    wire N__7357;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7301;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7245;
    wire N__7244;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7233;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7212;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6995;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6950;
    wire N__6947;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6663;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6578;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6509;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6446;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6398;
    wire N__6395;
    wire N__6394;
    wire N__6393;
    wire N__6392;
    wire N__6389;
    wire N__6388;
    wire N__6387;
    wire N__6386;
    wire N__6385;
    wire N__6382;
    wire N__6377;
    wire N__6374;
    wire N__6369;
    wire N__6362;
    wire N__6351;
    wire N__6350;
    wire N__6347;
    wire N__6346;
    wire N__6343;
    wire N__6342;
    wire N__6341;
    wire N__6336;
    wire N__6331;
    wire N__6328;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6284;
    wire N__6283;
    wire N__6282;
    wire N__6281;
    wire N__6280;
    wire N__6277;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6261;
    wire N__6254;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6233;
    wire N__6232;
    wire N__6231;
    wire N__6230;
    wire N__6229;
    wire N__6228;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6224;
    wire N__6221;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6132;
    wire N__6129;
    wire N__6128;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6093;
    wire N__6090;
    wire N__6089;
    wire N__6088;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6076;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6041;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5984;
    wire N__5983;
    wire N__5982;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5964;
    wire N__5955;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5939;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5935;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5833;
    wire N__5832;
    wire N__5831;
    wire N__5830;
    wire N__5825;
    wire N__5822;
    wire N__5821;
    wire N__5820;
    wire N__5817;
    wire N__5812;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5760;
    wire N__5753;
    wire N__5750;
    wire N__5749;
    wire N__5748;
    wire N__5745;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5702;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5636;
    wire N__5635;
    wire N__5632;
    wire N__5631;
    wire N__5628;
    wire N__5623;
    wire N__5618;
    wire N__5613;
    wire N__5610;
    wire N__5609;
    wire N__5602;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5561;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5477;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5450;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5430;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5388;
    wire N__5387;
    wire N__5386;
    wire N__5381;
    wire N__5380;
    wire N__5379;
    wire N__5378;
    wire N__5375;
    wire N__5374;
    wire N__5373;
    wire N__5372;
    wire N__5369;
    wire N__5368;
    wire N__5367;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5356;
    wire N__5353;
    wire N__5352;
    wire N__5349;
    wire N__5348;
    wire N__5345;
    wire N__5344;
    wire N__5343;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5338;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5323;
    wire N__5322;
    wire N__5321;
    wire N__5318;
    wire N__5313;
    wire N__5310;
    wire N__5309;
    wire N__5308;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5281;
    wire N__5276;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5251;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5229;
    wire N__5228;
    wire N__5223;
    wire N__5216;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5198;
    wire N__5195;
    wire N__5190;
    wire N__5185;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5158;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5140;
    wire N__5137;
    wire N__5132;
    wire N__5123;
    wire N__5112;
    wire N__5111;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5093;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5072;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5039;
    wire N__5036;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4566;
    wire N__4565;
    wire N__4564;
    wire N__4563;
    wire N__4562;
    wire N__4561;
    wire N__4560;
    wire N__4559;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4526;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4496;
    wire N__4493;
    wire N__4492;
    wire N__4487;
    wire N__4482;
    wire N__4481;
    wire N__4480;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4466;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4453;
    wire N__4452;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4448;
    wire N__4445;
    wire N__4440;
    wire N__4439;
    wire N__4438;
    wire N__4431;
    wire N__4428;
    wire N__4427;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4409;
    wire N__4404;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4392;
    wire N__4387;
    wire N__4382;
    wire N__4379;
    wire N__4374;
    wire N__4367;
    wire N__4364;
    wire N__4363;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4347;
    wire N__4342;
    wire N__4341;
    wire N__4338;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4290;
    wire N__4287;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3342;
    wire N__3339;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3306;
    wire N__3303;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2565;
    wire N__2562;
    wire N__2559;
    wire N__2558;
    wire N__2557;
    wire N__2556;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2545;
    wire N__2544;
    wire N__2543;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2535;
    wire N__2534;
    wire N__2527;
    wire N__2524;
    wire N__2521;
    wire N__2518;
    wire N__2515;
    wire N__2514;
    wire N__2513;
    wire N__2512;
    wire N__2511;
    wire N__2510;
    wire N__2509;
    wire N__2508;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2473;
    wire N__2472;
    wire N__2471;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2460;
    wire N__2459;
    wire N__2454;
    wire N__2451;
    wire N__2440;
    wire N__2437;
    wire N__2434;
    wire N__2431;
    wire N__2428;
    wire N__2427;
    wire N__2426;
    wire N__2423;
    wire N__2418;
    wire N__2415;
    wire N__2412;
    wire N__2411;
    wire N__2410;
    wire N__2409;
    wire N__2408;
    wire N__2407;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2374;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2362;
    wire N__2359;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2343;
    wire N__2332;
    wire N__2327;
    wire N__2322;
    wire N__2317;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire VCCG0;
    wire GNDG0;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire A_040_c_1;
    wire D_LL_AMIGA_in_2;
    wire un1_D_LL_AMIGA_2;
    wire RnW_c_i_0;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_LM_AMIGA_in_1;
    wire un1_D_LM_AMIGA_1;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire D_UM_040_in_4;
    wire D_LL_040_in_4;
    wire un1_D_UM_040_4;
    wire D_UU_040_in_3;
    wire D_LM_040_in_3;
    wire un1_D_UU_040_3;
    wire D_LM_040_in_6;
    wire D_UU_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LL_AMIGA_in_7;
    wire un1_D_LL_AMIGA_7;
    wire D_LL_040_in_1;
    wire D_UM_040_in_1;
    wire un1_D_UM_040_1;
    wire D_UU_040_in_7;
    wire D_LM_040_in_7;
    wire un1_D_UU_040_7;
    wire D_LL_AMIGA_in_4;
    wire un1_D_LL_AMIGA_4;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire D_LM_AMIGA_in_3;
    wire un1_D_LM_AMIGA_3;
    wire D_LM_AMIGA_in_5;
    wire un1_D_LM_AMIGA_5;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_LL_AMIGA_in_0;
    wire un1_D_LL_AMIGA_0;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire D_LM_AMIGA_in_2;
    wire un1_D_LM_AMIGA_2;
    wire D_LM_AMIGA_in_6;
    wire un1_D_LM_AMIGA_6;
    wire D_UU_040_in_1;
    wire D_LM_040_in_1;
    wire un1_D_UU_040_1;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_LL_AMIGA_in_6;
    wire un1_D_LL_AMIGA_6;
    wire D_LL_040_in_3;
    wire D_UM_040_in_3;
    wire un1_D_UM_040_3;
    wire D_LL_AMIGA_in_3;
    wire un1_D_LL_AMIGA_3;
    wire D_LL_AMIGA_in_1;
    wire un1_D_LL_AMIGA_1;
    wire D_LL_AMIGA_in_5;
    wire un1_D_LL_AMIGA_5;
    wire D_LM_AMIGA_in_0;
    wire un1_D_LM_AMIGA_0;
    wire un1_D_UM_AMIGA_0;
    wire \INVU111_CYCLE_SM.TA_ENC_net ;
    wire \U111_CYCLE_SM.RESETn_c_i ;
    wire \INVU111_CYCLE_SM.A_OUTC_net ;
    wire \U111_CYCLE_SM.A_OUTZ0 ;
    wire \U111_CYCLE_SM.A_OUT_0 ;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ;
    wire D_LM_AMIGA_in_4;
    wire un1_D_LM_AMIGA_4;
    wire \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ;
    wire CONSTANT_ONE_NET;
    wire D_LM_AMIGA_in_7;
    wire un1_D_LM_AMIGA_7;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire un1_D_UM_040_5;
    wire D_UU_040_in_5;
    wire D_LM_040_in_5;
    wire A_AMIGA_c_1;
    wire un1_D_UU_040_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire un1_D_UU_AMIGA_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire \U111_CYCLE_SM.TA_ENZ0 ;
    wire U111_CYCLE_SM_TAn_0_i;
    wire \U111_CYCLE_SM.un1_LW_TRANS_1_0 ;
    wire PORTSIZE_c;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ;
    wire \INVU111_CYCLE_SM.TS_ENC_net ;
    wire TS_CPUn_c;
    wire \U111_CYCLE_SM.TS_EN_5 ;
    wire \U111_CYCLE_SM.N_69_0 ;
    wire CLK40;
    wire \U111_CYCLE_SM.N_91_cascade_ ;
    wire \INVU111_CYCLE_SM.CYCLE_STATE_0C_net ;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire un1_D_UM_AMIGA_6;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ;
    wire RnW_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ;
    wire \U111_CYCLE_SM.LW_CYCLE_STARTZ0 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ;
    wire \INVU111_CYCLE_SM.LW_CYCLEC_net ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire TACKn_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.LW_CYCLE_0 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire D_UM_AMIGA_in_1;
    wire un1_D_UM_AMIGA_1;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire D_UU_AMIGA_in_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire un1_D_UU_AMIGA_3;
    wire un1_D_UM_AMIGA_2;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ;
    wire \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire un1_D_UU_AMIGA_1;
    wire D_UM_AMIGA_in_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire \U111_CYCLE_SM.LW_CYCLEZ0 ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__4989),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__8315));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__8315),
            .PACKAGEPIN(CLK40_IN));
    defparam D_UM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__8299),
            .DIN(N__8298),
            .DOUT(N__8297),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__8299),
            .PADOUT(N__8298),
            .PADIN(N__8297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5832),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__6801),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__8290),
            .DIN(N__8289),
            .DOUT(N__8288),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__8290),
            .PADOUT(N__8289),
            .PADIN(N__8288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2460),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__2802),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__8281),
            .DIN(N__8280),
            .DOUT(N__8279),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__8281),
            .PADOUT(N__8280),
            .PADIN(N__8279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2558),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__4278),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_ibuf_iopad (
            .OE(N__8272),
            .DIN(N__8271),
            .DOUT(N__8270),
            .PACKAGEPIN(TACKn));
    defparam TACKn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TACKn_ibuf_preio (
            .PADOEN(N__8272),
            .PADOUT(N__8271),
            .PADIN(N__8270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TACKn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__8263),
            .DIN(N__8262),
            .DOUT(N__8261),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__8263),
            .PADOUT(N__8262),
            .PADIN(N__8261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5936),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__4206),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__8254),
            .DIN(N__8253),
            .DOUT(N__8252),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__8254),
            .PADOUT(N__8253),
            .PADIN(N__8252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__8245),
            .DIN(N__8244),
            .DOUT(N__8243),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__8245),
            .PADOUT(N__8244),
            .PADIN(N__8243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5948),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__2823),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__8236),
            .DIN(N__8235),
            .DOUT(N__8234),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__8236),
            .PADOUT(N__8235),
            .PADIN(N__8234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2459),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__3069),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__8227),
            .DIN(N__8226),
            .DOUT(N__8225),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8227),
            .PADOUT(N__8226),
            .PADIN(N__8225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2543),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__3732),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__8218),
            .DIN(N__8217),
            .DOUT(N__8216),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__8218),
            .PADOUT(N__8217),
            .PADIN(N__8216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5885),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__6486),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__8209),
            .DIN(N__8208),
            .DOUT(N__8207),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__8209),
            .PADOUT(N__8208),
            .PADIN(N__8207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4990),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__8200),
            .DIN(N__8199),
            .DOUT(N__8198),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__8200),
            .PADOUT(N__8199),
            .PADIN(N__8198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__8191),
            .DIN(N__8190),
            .DOUT(N__8189),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8191),
            .PADOUT(N__8190),
            .PADIN(N__8189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2427),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__2985),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__8182),
            .DIN(N__8181),
            .DOUT(N__8180),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__8182),
            .PADOUT(N__8181),
            .PADIN(N__8180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5949),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__4176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__8173),
            .DIN(N__8172),
            .DOUT(N__8171),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8173),
            .PADOUT(N__8172),
            .PADIN(N__8171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2557),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__3108),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__8164),
            .DIN(N__8163),
            .DOUT(N__8162),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8164),
            .PADOUT(N__8163),
            .PADIN(N__8162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2472),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__3381),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__8155),
            .DIN(N__8154),
            .DOUT(N__8153),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__8155),
            .PADOUT(N__8154),
            .PADIN(N__8153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__8146),
            .DIN(N__8145),
            .DOUT(N__8144),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__8146),
            .PADOUT(N__8145),
            .PADIN(N__8144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5749),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__4920),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__8137),
            .DIN(N__8136),
            .DOUT(N__8135),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__8137),
            .PADOUT(N__8136),
            .PADIN(N__8135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5886),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__6639),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__8128),
            .DIN(N__8127),
            .DOUT(N__8126),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__8128),
            .PADOUT(N__8127),
            .PADIN(N__8126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5478),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__8119),
            .DIN(N__8118),
            .DOUT(N__8117),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__8119),
            .PADOUT(N__8118),
            .PADIN(N__8117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2407),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__4743),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__8110),
            .DIN(N__8109),
            .DOUT(N__8108),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__8110),
            .PADOUT(N__8109),
            .PADIN(N__8108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__8101),
            .DIN(N__8100),
            .DOUT(N__8099),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8101),
            .PADOUT(N__8100),
            .PADIN(N__8099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2409),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__4797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__8092),
            .DIN(N__8091),
            .DOUT(N__8090),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__8092),
            .PADOUT(N__8091),
            .PADIN(N__8090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5830),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__6882),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__8083),
            .DIN(N__8082),
            .DOUT(N__8081),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__8083),
            .PADOUT(N__8082),
            .PADIN(N__8081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5430),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__8074),
            .DIN(N__8073),
            .DOUT(N__8072),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__8074),
            .PADOUT(N__8073),
            .PADIN(N__8072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5477),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__8065),
            .DIN(N__8064),
            .DOUT(N__8063),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__8065),
            .PADOUT(N__8064),
            .PADIN(N__8063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5911),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__3459),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__8056),
            .DIN(N__8055),
            .DOUT(N__8054),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__8056),
            .PADOUT(N__8055),
            .PADIN(N__8054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5983),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__3573),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__8047),
            .DIN(N__8046),
            .DOUT(N__8045),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__8047),
            .PADOUT(N__8046),
            .PADIN(N__8045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2408),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__4875),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__8038),
            .DIN(N__8037),
            .DOUT(N__8036),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__8038),
            .PADOUT(N__8037),
            .PADIN(N__8036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2555),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__2655),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__8029),
            .DIN(N__8028),
            .DOUT(N__8027),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__8029),
            .PADOUT(N__8028),
            .PADIN(N__8027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5967),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__8020),
            .DIN(N__8019),
            .DOUT(N__8018),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__8020),
            .PADOUT(N__8019),
            .PADIN(N__8018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2511),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__4617),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__8011),
            .DIN(N__8010),
            .DOUT(N__8009),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__8011),
            .PADOUT(N__8010),
            .PADIN(N__8009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5939),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__6900),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__8002),
            .DIN(N__8001),
            .DOUT(N__8000),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__8002),
            .PADOUT(N__8001),
            .PADIN(N__8000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__7993),
            .DIN(N__7992),
            .DOUT(N__7991),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__7993),
            .PADOUT(N__7992),
            .PADIN(N__7991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5744),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__3228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__7984),
            .DIN(N__7983),
            .DOUT(N__7982),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__7984),
            .PADOUT(N__7983),
            .PADIN(N__7982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5887),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__6981),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__7975),
            .DIN(N__7974),
            .DOUT(N__7973),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__7975),
            .PADOUT(N__7974),
            .PADIN(N__7973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__7966),
            .DIN(N__7965),
            .DOUT(N__7964),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__7966),
            .PADOUT(N__7965),
            .PADIN(N__7964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5982),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__3654),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__7957),
            .DIN(N__7956),
            .DOUT(N__7955),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__7957),
            .PADOUT(N__7956),
            .PADIN(N__7955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2508),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__3800),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__7948),
            .DIN(N__7947),
            .DOUT(N__7946),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__7948),
            .PADOUT(N__7947),
            .PADIN(N__7946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2535),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__4659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__7939),
            .DIN(N__7938),
            .DOUT(N__7937),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__7939),
            .PADOUT(N__7938),
            .PADIN(N__7937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5833),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__7059),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__7930),
            .DIN(N__7929),
            .DOUT(N__7928),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__7930),
            .PADOUT(N__7929),
            .PADIN(N__7928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2559),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__2940),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__7921),
            .DIN(N__7920),
            .DOUT(N__7919),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7921),
            .PADOUT(N__7920),
            .PADIN(N__7919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2426),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__3987),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__7912),
            .DIN(N__7911),
            .DOUT(N__7910),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__7912),
            .PADOUT(N__7911),
            .PADIN(N__7910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5947),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__3264),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__7903),
            .DIN(N__7902),
            .DOUT(N__7901),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__7903),
            .PADOUT(N__7902),
            .PADIN(N__7901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5950),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__3612),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__7894),
            .DIN(N__7893),
            .DOUT(N__7892),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__7894),
            .PADOUT(N__7893),
            .PADIN(N__7892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2410),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__3156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__7885),
            .DIN(N__7884),
            .DOUT(N__7883),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__7885),
            .PADOUT(N__7884),
            .PADIN(N__7883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2556),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__2856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__7876),
            .DIN(N__7875),
            .DOUT(N__7874),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__7876),
            .PADOUT(N__7875),
            .PADIN(N__7874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2512),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__2736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__7867),
            .DIN(N__7866),
            .DOUT(N__7865),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__7867),
            .PADOUT(N__7866),
            .PADIN(N__7865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5888),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__6561),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__7858),
            .DIN(N__7857),
            .DOUT(N__7856),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__7858),
            .PADOUT(N__7857),
            .PADIN(N__7856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6195),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__7849),
            .DIN(N__7848),
            .DOUT(N__7847),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__7849),
            .PADOUT(N__7848),
            .PADIN(N__7847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5777),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__6465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__7840),
            .DIN(N__7839),
            .DOUT(N__7838),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__7840),
            .PADOUT(N__7839),
            .PADIN(N__7838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5968),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__2583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__7831),
            .DIN(N__7830),
            .DOUT(N__7829),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__7831),
            .PADOUT(N__7830),
            .PADIN(N__7829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__7822),
            .DIN(N__7821),
            .DOUT(N__7820),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__7822),
            .PADOUT(N__7821),
            .PADIN(N__7820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6188),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__7813),
            .DIN(N__7812),
            .DOUT(N__7811),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__7813),
            .PADOUT(N__7812),
            .PADIN(N__7811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2509),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__3534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__7804),
            .DIN(N__7803),
            .DOUT(N__7802),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__7804),
            .PADOUT(N__7803),
            .PADIN(N__7802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2545),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__3027),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__7795),
            .DIN(N__7794),
            .DOUT(N__7793),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__7795),
            .PADOUT(N__7794),
            .PADIN(N__7793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2406),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__3867),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7786),
            .DIN(N__7785),
            .DOUT(N__7784),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7786),
            .PADOUT(N__7785),
            .PADIN(N__7784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__7777),
            .DIN(N__7776),
            .DOUT(N__7775),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__7777),
            .PADOUT(N__7776),
            .PADIN(N__7775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2514),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__2919),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RnW_ibuf_iopad.PULLUP=1'b1;
    IO_PAD RnW_ibuf_iopad (
            .OE(N__7768),
            .DIN(N__7767),
            .DOUT(N__7766),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__7768),
            .PADOUT(N__7767),
            .PADIN(N__7766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__7759),
            .DIN(N__7758),
            .DOUT(N__7757),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__7759),
            .PADOUT(N__7758),
            .PADIN(N__7757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5821),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__7750),
            .DIN(N__7749),
            .DOUT(N__7748),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__7750),
            .PADOUT(N__7749),
            .PADIN(N__7748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5748),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__6009),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TAn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TAn_obuf_iopad (
            .OE(N__7741),
            .DIN(N__7740),
            .DOUT(N__7739),
            .PACKAGEPIN(TAn));
    defparam TAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TAn_obuf_preio (
            .PADOEN(N__7741),
            .PADOUT(N__7740),
            .PADIN(N__7739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5429),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__7732),
            .DIN(N__7731),
            .DOUT(N__7730),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__7732),
            .PADOUT(N__7731),
            .PADIN(N__7730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4998),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_6_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__7723),
            .DIN(N__7722),
            .DOUT(N__7721),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__7723),
            .PADOUT(N__7722),
            .PADIN(N__7721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5951),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__3825),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_5_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__7714),
            .DIN(N__7713),
            .DOUT(N__7712),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__7714),
            .PADOUT(N__7713),
            .PADIN(N__7712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2411),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__4725),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__7705),
            .DIN(N__7704),
            .DOUT(N__7703),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__7705),
            .PADOUT(N__7704),
            .PADIN(N__7703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2471),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__2238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__7696),
            .DIN(N__7695),
            .DOUT(N__7694),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__7696),
            .PADOUT(N__7695),
            .PADIN(N__7694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5938),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__5493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__7687),
            .DIN(N__7686),
            .DOUT(N__7685),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7687),
            .PADOUT(N__7686),
            .PADIN(N__7685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2470),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__3905),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__7678),
            .DIN(N__7677),
            .DOUT(N__7676),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__7678),
            .PADOUT(N__7677),
            .PADIN(N__7676),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_3_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__7669),
            .DIN(N__7668),
            .DOUT(N__7667),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__7669),
            .PADOUT(N__7668),
            .PADIN(N__7667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5984),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__3693),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__7660),
            .DIN(N__7659),
            .DOUT(N__7658),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__7660),
            .PADOUT(N__7659),
            .PADIN(N__7658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5946),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__3195),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TSn_obuf_iopad.PULLUP=1'b1;
    IO_PAD TSn_obuf_iopad (
            .OE(N__7651),
            .DIN(N__7650),
            .DOUT(N__7649),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__7651),
            .PADOUT(N__7650),
            .PADIN(N__7649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3291),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__7642),
            .DIN(N__7641),
            .DOUT(N__7640),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7642),
            .PADOUT(N__7641),
            .PADIN(N__7640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2544),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__4830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_AMIGA_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__7633),
            .DIN(N__7632),
            .DOUT(N__7631),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__7633),
            .PADOUT(N__7632),
            .PADIN(N__7631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2513),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__2700),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__7624),
            .DIN(N__7623),
            .DOUT(N__7622),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__7624),
            .PADOUT(N__7623),
            .PADIN(N__7622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__7615),
            .DIN(N__7614),
            .DOUT(N__7613),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__7615),
            .PADOUT(N__7614),
            .PADIN(N__7613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2622),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LM_040_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__7606),
            .DIN(N__7605),
            .DOUT(N__7604),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__7606),
            .PADOUT(N__7605),
            .PADIN(N__7604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5866),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__4032),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__7597),
            .DIN(N__7596),
            .DOUT(N__7595),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__7597),
            .PADOUT(N__7596),
            .PADIN(N__7595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5831),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__6717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7588),
            .DIN(N__7587),
            .DOUT(N__7586),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7588),
            .PADOUT(N__7587),
            .PADIN(N__7586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_1_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__7579),
            .DIN(N__7578),
            .DOUT(N__7577),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__7579),
            .PADOUT(N__7578),
            .PADIN(N__7577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2542),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__3945),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__7570),
            .DIN(N__7569),
            .DOUT(N__7568),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__7570),
            .PADOUT(N__7569),
            .PADIN(N__7568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5476),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__7561),
            .DIN(N__7560),
            .DOUT(N__7559),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__7561),
            .PADOUT(N__7560),
            .PADIN(N__7559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5820),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__4155),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_AMIGA_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__7552),
            .DIN(N__7551),
            .DOUT(N__7550),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__7552),
            .PADOUT(N__7551),
            .PADIN(N__7550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2510),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__2283),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_AMIGA_iobuf_4_iopad.PULLUP=1'b1;
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__7543),
            .DIN(N__7542),
            .DOUT(N__7541),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__7543),
            .PADOUT(N__7542),
            .PADIN(N__7541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2534),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__3342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_7_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__7534),
            .DIN(N__7533),
            .DOUT(N__7532),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__7534),
            .PADOUT(N__7533),
            .PADIN(N__7532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5935),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__7290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SIZ_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7525),
            .DIN(N__7524),
            .DOUT(N__7523),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7525),
            .PADOUT(N__7524),
            .PADIN(N__7523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_LL_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__7516),
            .DIN(N__7515),
            .DOUT(N__7514),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__7516),
            .PADOUT(N__7515),
            .PADIN(N__7514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5985),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__3312),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UM_AMIGA_iobuf_2_iopad.PULLUP=1'b1;
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__7507),
            .DIN(N__7506),
            .DOUT(N__7505),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__7507),
            .PADOUT(N__7506),
            .PADIN(N__7505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2473),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__3492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam D_UU_040_iobuf_0_iopad.PULLUP=1'b1;
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__7498),
            .DIN(N__7497),
            .DOUT(N__7496),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__7498),
            .PADOUT(N__7497),
            .PADIN(N__7496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5937),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__7134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1948 (
            .O(N__7479),
            .I(N__7473));
    InMux I__1947 (
            .O(N__7478),
            .I(N__7473));
    LocalMux I__1946 (
            .O(N__7473),
            .I(N__7457));
    InMux I__1945 (
            .O(N__7472),
            .I(N__7450));
    InMux I__1944 (
            .O(N__7471),
            .I(N__7450));
    InMux I__1943 (
            .O(N__7470),
            .I(N__7450));
    InMux I__1942 (
            .O(N__7469),
            .I(N__7445));
    InMux I__1941 (
            .O(N__7468),
            .I(N__7445));
    InMux I__1940 (
            .O(N__7467),
            .I(N__7440));
    InMux I__1939 (
            .O(N__7466),
            .I(N__7440));
    InMux I__1938 (
            .O(N__7465),
            .I(N__7435));
    InMux I__1937 (
            .O(N__7464),
            .I(N__7435));
    InMux I__1936 (
            .O(N__7463),
            .I(N__7430));
    InMux I__1935 (
            .O(N__7462),
            .I(N__7430));
    InMux I__1934 (
            .O(N__7461),
            .I(N__7427));
    CascadeMux I__1933 (
            .O(N__7460),
            .I(N__7420));
    Sp12to4 I__1932 (
            .O(N__7457),
            .I(N__7416));
    LocalMux I__1931 (
            .O(N__7450),
            .I(N__7411));
    LocalMux I__1930 (
            .O(N__7445),
            .I(N__7411));
    LocalMux I__1929 (
            .O(N__7440),
            .I(N__7404));
    LocalMux I__1928 (
            .O(N__7435),
            .I(N__7404));
    LocalMux I__1927 (
            .O(N__7430),
            .I(N__7404));
    LocalMux I__1926 (
            .O(N__7427),
            .I(N__7401));
    InMux I__1925 (
            .O(N__7426),
            .I(N__7398));
    InMux I__1924 (
            .O(N__7425),
            .I(N__7395));
    CascadeMux I__1923 (
            .O(N__7424),
            .I(N__7392));
    InMux I__1922 (
            .O(N__7423),
            .I(N__7389));
    InMux I__1921 (
            .O(N__7420),
            .I(N__7384));
    InMux I__1920 (
            .O(N__7419),
            .I(N__7384));
    Span12Mux_v I__1919 (
            .O(N__7416),
            .I(N__7380));
    Span4Mux_v I__1918 (
            .O(N__7411),
            .I(N__7377));
    Span4Mux_v I__1917 (
            .O(N__7404),
            .I(N__7368));
    Span4Mux_v I__1916 (
            .O(N__7401),
            .I(N__7368));
    LocalMux I__1915 (
            .O(N__7398),
            .I(N__7368));
    LocalMux I__1914 (
            .O(N__7395),
            .I(N__7368));
    InMux I__1913 (
            .O(N__7392),
            .I(N__7365));
    LocalMux I__1912 (
            .O(N__7389),
            .I(N__7360));
    LocalMux I__1911 (
            .O(N__7384),
            .I(N__7360));
    InMux I__1910 (
            .O(N__7383),
            .I(N__7357));
    Odrv12 I__1909 (
            .O(N__7380),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1908 (
            .O(N__7377),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1907 (
            .O(N__7368),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1906 (
            .O(N__7365),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    Odrv4 I__1905 (
            .O(N__7360),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    LocalMux I__1904 (
            .O(N__7357),
            .I(\U111_CYCLE_SM.LW_CYCLEZ0 ));
    InMux I__1903 (
            .O(N__7344),
            .I(N__7341));
    LocalMux I__1902 (
            .O(N__7341),
            .I(N__7338));
    Odrv12 I__1901 (
            .O(N__7338),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__1900 (
            .O(N__7335),
            .I(N__7331));
    InMux I__1899 (
            .O(N__7334),
            .I(N__7328));
    LocalMux I__1898 (
            .O(N__7331),
            .I(N__7324));
    LocalMux I__1897 (
            .O(N__7328),
            .I(N__7321));
    InMux I__1896 (
            .O(N__7327),
            .I(N__7318));
    Span4Mux_v I__1895 (
            .O(N__7324),
            .I(N__7315));
    Span4Mux_v I__1894 (
            .O(N__7321),
            .I(N__7312));
    LocalMux I__1893 (
            .O(N__7318),
            .I(N__7309));
    Span4Mux_h I__1892 (
            .O(N__7315),
            .I(N__7306));
    Span4Mux_v I__1891 (
            .O(N__7312),
            .I(N__7301));
    Span4Mux_v I__1890 (
            .O(N__7309),
            .I(N__7301));
    Sp12to4 I__1889 (
            .O(N__7306),
            .I(N__7296));
    Sp12to4 I__1888 (
            .O(N__7301),
            .I(N__7296));
    Span12Mux_h I__1887 (
            .O(N__7296),
            .I(N__7293));
    Odrv12 I__1886 (
            .O(N__7293),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1885 (
            .O(N__7290),
            .I(N__7287));
    LocalMux I__1884 (
            .O(N__7287),
            .I(N__7284));
    Span12Mux_s11_v I__1883 (
            .O(N__7284),
            .I(N__7281));
    Span12Mux_h I__1882 (
            .O(N__7281),
            .I(N__7278));
    Odrv12 I__1881 (
            .O(N__7278),
            .I(un1_D_UU_AMIGA_7));
    CEMux I__1880 (
            .O(N__7275),
            .I(N__7268));
    CEMux I__1879 (
            .O(N__7274),
            .I(N__7265));
    CEMux I__1878 (
            .O(N__7273),
            .I(N__7262));
    CEMux I__1877 (
            .O(N__7272),
            .I(N__7259));
    CEMux I__1876 (
            .O(N__7271),
            .I(N__7256));
    LocalMux I__1875 (
            .O(N__7268),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    LocalMux I__1874 (
            .O(N__7265),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    LocalMux I__1873 (
            .O(N__7262),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    LocalMux I__1872 (
            .O(N__7259),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    LocalMux I__1871 (
            .O(N__7256),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ));
    SRMux I__1870 (
            .O(N__7245),
            .I(N__7240));
    SRMux I__1869 (
            .O(N__7244),
            .I(N__7237));
    SRMux I__1868 (
            .O(N__7243),
            .I(N__7233));
    LocalMux I__1867 (
            .O(N__7240),
            .I(N__7229));
    LocalMux I__1866 (
            .O(N__7237),
            .I(N__7226));
    SRMux I__1865 (
            .O(N__7236),
            .I(N__7223));
    LocalMux I__1864 (
            .O(N__7233),
            .I(N__7220));
    SRMux I__1863 (
            .O(N__7232),
            .I(N__7217));
    Span4Mux_v I__1862 (
            .O(N__7229),
            .I(N__7212));
    Span4Mux_v I__1861 (
            .O(N__7226),
            .I(N__7212));
    LocalMux I__1860 (
            .O(N__7223),
            .I(N__7205));
    Span4Mux_v I__1859 (
            .O(N__7220),
            .I(N__7205));
    LocalMux I__1858 (
            .O(N__7217),
            .I(N__7205));
    Span4Mux_h I__1857 (
            .O(N__7212),
            .I(N__7202));
    Span4Mux_v I__1856 (
            .O(N__7205),
            .I(N__7199));
    Odrv4 I__1855 (
            .O(N__7202),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    Odrv4 I__1854 (
            .O(N__7199),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ));
    InMux I__1853 (
            .O(N__7194),
            .I(N__7191));
    LocalMux I__1852 (
            .O(N__7191),
            .I(N__7188));
    Odrv12 I__1851 (
            .O(N__7188),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    CascadeMux I__1850 (
            .O(N__7185),
            .I(N__7182));
    InMux I__1849 (
            .O(N__7182),
            .I(N__7179));
    LocalMux I__1848 (
            .O(N__7179),
            .I(N__7175));
    InMux I__1847 (
            .O(N__7178),
            .I(N__7172));
    Span4Mux_v I__1846 (
            .O(N__7175),
            .I(N__7168));
    LocalMux I__1845 (
            .O(N__7172),
            .I(N__7165));
    InMux I__1844 (
            .O(N__7171),
            .I(N__7162));
    Span4Mux_v I__1843 (
            .O(N__7168),
            .I(N__7159));
    Span4Mux_v I__1842 (
            .O(N__7165),
            .I(N__7154));
    LocalMux I__1841 (
            .O(N__7162),
            .I(N__7154));
    Sp12to4 I__1840 (
            .O(N__7159),
            .I(N__7151));
    Sp12to4 I__1839 (
            .O(N__7154),
            .I(N__7148));
    Span12Mux_h I__1838 (
            .O(N__7151),
            .I(N__7145));
    Span12Mux_v I__1837 (
            .O(N__7148),
            .I(N__7142));
    Span12Mux_v I__1836 (
            .O(N__7145),
            .I(N__7137));
    Span12Mux_h I__1835 (
            .O(N__7142),
            .I(N__7137));
    Odrv12 I__1834 (
            .O(N__7137),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1833 (
            .O(N__7134),
            .I(N__7131));
    LocalMux I__1832 (
            .O(N__7131),
            .I(N__7128));
    Span4Mux_s3_v I__1831 (
            .O(N__7128),
            .I(N__7125));
    Span4Mux_h I__1830 (
            .O(N__7125),
            .I(N__7122));
    Sp12to4 I__1829 (
            .O(N__7122),
            .I(N__7119));
    Span12Mux_s8_v I__1828 (
            .O(N__7119),
            .I(N__7116));
    Odrv12 I__1827 (
            .O(N__7116),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1826 (
            .O(N__7113),
            .I(N__7110));
    LocalMux I__1825 (
            .O(N__7110),
            .I(N__7106));
    InMux I__1824 (
            .O(N__7109),
            .I(N__7103));
    Span4Mux_v I__1823 (
            .O(N__7106),
            .I(N__7099));
    LocalMux I__1822 (
            .O(N__7103),
            .I(N__7096));
    InMux I__1821 (
            .O(N__7102),
            .I(N__7093));
    Span4Mux_v I__1820 (
            .O(N__7099),
            .I(N__7090));
    Span4Mux_v I__1819 (
            .O(N__7096),
            .I(N__7085));
    LocalMux I__1818 (
            .O(N__7093),
            .I(N__7085));
    Span4Mux_v I__1817 (
            .O(N__7090),
            .I(N__7082));
    Span4Mux_v I__1816 (
            .O(N__7085),
            .I(N__7079));
    Sp12to4 I__1815 (
            .O(N__7082),
            .I(N__7074));
    Sp12to4 I__1814 (
            .O(N__7079),
            .I(N__7074));
    Span12Mux_h I__1813 (
            .O(N__7074),
            .I(N__7071));
    Odrv12 I__1812 (
            .O(N__7071),
            .I(D_UU_AMIGA_in_1));
    InMux I__1811 (
            .O(N__7068),
            .I(N__7065));
    LocalMux I__1810 (
            .O(N__7065),
            .I(N__7062));
    Odrv12 I__1809 (
            .O(N__7062),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    IoInMux I__1808 (
            .O(N__7059),
            .I(N__7056));
    LocalMux I__1807 (
            .O(N__7056),
            .I(N__7053));
    IoSpan4Mux I__1806 (
            .O(N__7053),
            .I(N__7050));
    IoSpan4Mux I__1805 (
            .O(N__7050),
            .I(N__7047));
    Span4Mux_s2_h I__1804 (
            .O(N__7047),
            .I(N__7044));
    Sp12to4 I__1803 (
            .O(N__7044),
            .I(N__7041));
    Odrv12 I__1802 (
            .O(N__7041),
            .I(un1_D_UU_AMIGA_1));
    InMux I__1801 (
            .O(N__7038),
            .I(N__7035));
    LocalMux I__1800 (
            .O(N__7035),
            .I(N__7031));
    InMux I__1799 (
            .O(N__7034),
            .I(N__7027));
    Span4Mux_v I__1798 (
            .O(N__7031),
            .I(N__7024));
    InMux I__1797 (
            .O(N__7030),
            .I(N__7021));
    LocalMux I__1796 (
            .O(N__7027),
            .I(N__7018));
    Sp12to4 I__1795 (
            .O(N__7024),
            .I(N__7015));
    LocalMux I__1794 (
            .O(N__7021),
            .I(N__7012));
    Span12Mux_v I__1793 (
            .O(N__7018),
            .I(N__7009));
    Span12Mux_h I__1792 (
            .O(N__7015),
            .I(N__7006));
    Span12Mux_s7_v I__1791 (
            .O(N__7012),
            .I(N__7003));
    Span12Mux_h I__1790 (
            .O(N__7009),
            .I(N__7000));
    Span12Mux_v I__1789 (
            .O(N__7006),
            .I(N__6995));
    Span12Mux_h I__1788 (
            .O(N__7003),
            .I(N__6995));
    Odrv12 I__1787 (
            .O(N__7000),
            .I(D_UM_AMIGA_in_5));
    Odrv12 I__1786 (
            .O(N__6995),
            .I(D_UM_AMIGA_in_5));
    InMux I__1785 (
            .O(N__6990),
            .I(N__6987));
    LocalMux I__1784 (
            .O(N__6987),
            .I(N__6984));
    Odrv12 I__1783 (
            .O(N__6984),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    IoInMux I__1782 (
            .O(N__6981),
            .I(N__6978));
    LocalMux I__1781 (
            .O(N__6978),
            .I(N__6975));
    Span4Mux_s2_v I__1780 (
            .O(N__6975),
            .I(N__6972));
    Span4Mux_h I__1779 (
            .O(N__6972),
            .I(N__6969));
    Span4Mux_v I__1778 (
            .O(N__6969),
            .I(N__6966));
    Sp12to4 I__1777 (
            .O(N__6966),
            .I(N__6963));
    Odrv12 I__1776 (
            .O(N__6963),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1775 (
            .O(N__6960),
            .I(N__6957));
    LocalMux I__1774 (
            .O(N__6957),
            .I(N__6954));
    Odrv12 I__1773 (
            .O(N__6954),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    CascadeMux I__1772 (
            .O(N__6951),
            .I(N__6947));
    InMux I__1771 (
            .O(N__6950),
            .I(N__6943));
    InMux I__1770 (
            .O(N__6947),
            .I(N__6940));
    InMux I__1769 (
            .O(N__6946),
            .I(N__6937));
    LocalMux I__1768 (
            .O(N__6943),
            .I(N__6934));
    LocalMux I__1767 (
            .O(N__6940),
            .I(N__6931));
    LocalMux I__1766 (
            .O(N__6937),
            .I(N__6928));
    Span4Mux_v I__1765 (
            .O(N__6934),
            .I(N__6925));
    Span4Mux_v I__1764 (
            .O(N__6931),
            .I(N__6922));
    Span4Mux_v I__1763 (
            .O(N__6928),
            .I(N__6919));
    Sp12to4 I__1762 (
            .O(N__6925),
            .I(N__6914));
    Sp12to4 I__1761 (
            .O(N__6922),
            .I(N__6914));
    Sp12to4 I__1760 (
            .O(N__6919),
            .I(N__6911));
    Span12Mux_h I__1759 (
            .O(N__6914),
            .I(N__6908));
    Span12Mux_h I__1758 (
            .O(N__6911),
            .I(N__6905));
    Odrv12 I__1757 (
            .O(N__6908),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__1756 (
            .O(N__6905),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1755 (
            .O(N__6900),
            .I(N__6897));
    LocalMux I__1754 (
            .O(N__6897),
            .I(N__6894));
    Span4Mux_s3_v I__1753 (
            .O(N__6894),
            .I(N__6891));
    Span4Mux_h I__1752 (
            .O(N__6891),
            .I(N__6888));
    Span4Mux_h I__1751 (
            .O(N__6888),
            .I(N__6885));
    Odrv4 I__1750 (
            .O(N__6885),
            .I(un1_D_UU_AMIGA_4));
    IoInMux I__1749 (
            .O(N__6882),
            .I(N__6879));
    LocalMux I__1748 (
            .O(N__6879),
            .I(N__6876));
    IoSpan4Mux I__1747 (
            .O(N__6876),
            .I(N__6873));
    Span4Mux_s2_h I__1746 (
            .O(N__6873),
            .I(N__6870));
    Sp12to4 I__1745 (
            .O(N__6870),
            .I(N__6867));
    Span12Mux_h I__1744 (
            .O(N__6867),
            .I(N__6864));
    Odrv12 I__1743 (
            .O(N__6864),
            .I(un1_D_UM_AMIGA_1));
    CascadeMux I__1742 (
            .O(N__6861),
            .I(N__6858));
    InMux I__1741 (
            .O(N__6858),
            .I(N__6855));
    LocalMux I__1740 (
            .O(N__6855),
            .I(N__6850));
    InMux I__1739 (
            .O(N__6854),
            .I(N__6847));
    InMux I__1738 (
            .O(N__6853),
            .I(N__6844));
    Span4Mux_v I__1737 (
            .O(N__6850),
            .I(N__6841));
    LocalMux I__1736 (
            .O(N__6847),
            .I(N__6836));
    LocalMux I__1735 (
            .O(N__6844),
            .I(N__6836));
    Span4Mux_v I__1734 (
            .O(N__6841),
            .I(N__6833));
    Span4Mux_v I__1733 (
            .O(N__6836),
            .I(N__6830));
    Sp12to4 I__1732 (
            .O(N__6833),
            .I(N__6827));
    Span4Mux_v I__1731 (
            .O(N__6830),
            .I(N__6824));
    Span12Mux_h I__1730 (
            .O(N__6827),
            .I(N__6821));
    Sp12to4 I__1729 (
            .O(N__6824),
            .I(N__6818));
    Span12Mux_v I__1728 (
            .O(N__6821),
            .I(N__6813));
    Span12Mux_h I__1727 (
            .O(N__6818),
            .I(N__6813));
    Odrv12 I__1726 (
            .O(N__6813),
            .I(D_UM_AMIGA_in_3));
    InMux I__1725 (
            .O(N__6810),
            .I(N__6807));
    LocalMux I__1724 (
            .O(N__6807),
            .I(N__6804));
    Odrv4 I__1723 (
            .O(N__6804),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1722 (
            .O(N__6801),
            .I(N__6798));
    LocalMux I__1721 (
            .O(N__6798),
            .I(N__6795));
    Span4Mux_s0_h I__1720 (
            .O(N__6795),
            .I(N__6792));
    Span4Mux_h I__1719 (
            .O(N__6792),
            .I(N__6789));
    Sp12to4 I__1718 (
            .O(N__6789),
            .I(N__6786));
    Span12Mux_s11_v I__1717 (
            .O(N__6786),
            .I(N__6783));
    Span12Mux_h I__1716 (
            .O(N__6783),
            .I(N__6780));
    Odrv12 I__1715 (
            .O(N__6780),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1714 (
            .O(N__6777),
            .I(N__6773));
    CascadeMux I__1713 (
            .O(N__6776),
            .I(N__6770));
    LocalMux I__1712 (
            .O(N__6773),
            .I(N__6767));
    InMux I__1711 (
            .O(N__6770),
            .I(N__6763));
    Span4Mux_v I__1710 (
            .O(N__6767),
            .I(N__6760));
    InMux I__1709 (
            .O(N__6766),
            .I(N__6757));
    LocalMux I__1708 (
            .O(N__6763),
            .I(N__6754));
    Span4Mux_v I__1707 (
            .O(N__6760),
            .I(N__6749));
    LocalMux I__1706 (
            .O(N__6757),
            .I(N__6749));
    Span4Mux_v I__1705 (
            .O(N__6754),
            .I(N__6746));
    Span4Mux_v I__1704 (
            .O(N__6749),
            .I(N__6743));
    Sp12to4 I__1703 (
            .O(N__6746),
            .I(N__6740));
    Sp12to4 I__1702 (
            .O(N__6743),
            .I(N__6737));
    Span12Mux_v I__1701 (
            .O(N__6740),
            .I(N__6734));
    Span12Mux_h I__1700 (
            .O(N__6737),
            .I(N__6731));
    Odrv12 I__1699 (
            .O(N__6734),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1698 (
            .O(N__6731),
            .I(D_UM_AMIGA_in_7));
    InMux I__1697 (
            .O(N__6726),
            .I(N__6723));
    LocalMux I__1696 (
            .O(N__6723),
            .I(N__6720));
    Odrv12 I__1695 (
            .O(N__6720),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1694 (
            .O(N__6717),
            .I(N__6714));
    LocalMux I__1693 (
            .O(N__6714),
            .I(N__6711));
    IoSpan4Mux I__1692 (
            .O(N__6711),
            .I(N__6708));
    Span4Mux_s3_h I__1691 (
            .O(N__6708),
            .I(N__6705));
    Span4Mux_h I__1690 (
            .O(N__6705),
            .I(N__6702));
    Span4Mux_h I__1689 (
            .O(N__6702),
            .I(N__6699));
    Span4Mux_h I__1688 (
            .O(N__6699),
            .I(N__6696));
    Odrv4 I__1687 (
            .O(N__6696),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1686 (
            .O(N__6693),
            .I(N__6690));
    LocalMux I__1685 (
            .O(N__6690),
            .I(N__6687));
    Odrv12 I__1684 (
            .O(N__6687),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1683 (
            .O(N__6684),
            .I(N__6681));
    LocalMux I__1682 (
            .O(N__6681),
            .I(N__6678));
    Span4Mux_v I__1681 (
            .O(N__6678),
            .I(N__6675));
    Span4Mux_v I__1680 (
            .O(N__6675),
            .I(N__6671));
    InMux I__1679 (
            .O(N__6674),
            .I(N__6668));
    Span4Mux_v I__1678 (
            .O(N__6671),
            .I(N__6663));
    LocalMux I__1677 (
            .O(N__6668),
            .I(N__6663));
    Span4Mux_h I__1676 (
            .O(N__6663),
            .I(N__6659));
    InMux I__1675 (
            .O(N__6662),
            .I(N__6656));
    Span4Mux_v I__1674 (
            .O(N__6659),
            .I(N__6651));
    LocalMux I__1673 (
            .O(N__6656),
            .I(N__6651));
    Span4Mux_v I__1672 (
            .O(N__6651),
            .I(N__6648));
    Sp12to4 I__1671 (
            .O(N__6648),
            .I(N__6645));
    Span12Mux_h I__1670 (
            .O(N__6645),
            .I(N__6642));
    Odrv12 I__1669 (
            .O(N__6642),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1668 (
            .O(N__6639),
            .I(N__6636));
    LocalMux I__1667 (
            .O(N__6636),
            .I(N__6633));
    Span4Mux_s3_v I__1666 (
            .O(N__6633),
            .I(N__6630));
    Span4Mux_v I__1665 (
            .O(N__6630),
            .I(N__6627));
    Sp12to4 I__1664 (
            .O(N__6627),
            .I(N__6624));
    Span12Mux_h I__1663 (
            .O(N__6624),
            .I(N__6621));
    Odrv12 I__1662 (
            .O(N__6621),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1661 (
            .O(N__6618),
            .I(N__6615));
    LocalMux I__1660 (
            .O(N__6615),
            .I(N__6612));
    Odrv12 I__1659 (
            .O(N__6612),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    CascadeMux I__1658 (
            .O(N__6609),
            .I(N__6605));
    InMux I__1657 (
            .O(N__6608),
            .I(N__6602));
    InMux I__1656 (
            .O(N__6605),
            .I(N__6599));
    LocalMux I__1655 (
            .O(N__6602),
            .I(N__6596));
    LocalMux I__1654 (
            .O(N__6599),
            .I(N__6592));
    Span4Mux_v I__1653 (
            .O(N__6596),
            .I(N__6589));
    InMux I__1652 (
            .O(N__6595),
            .I(N__6586));
    Span4Mux_v I__1651 (
            .O(N__6592),
            .I(N__6583));
    Span4Mux_v I__1650 (
            .O(N__6589),
            .I(N__6578));
    LocalMux I__1649 (
            .O(N__6586),
            .I(N__6578));
    Span4Mux_v I__1648 (
            .O(N__6583),
            .I(N__6573));
    Span4Mux_h I__1647 (
            .O(N__6578),
            .I(N__6573));
    Span4Mux_v I__1646 (
            .O(N__6573),
            .I(N__6570));
    Span4Mux_h I__1645 (
            .O(N__6570),
            .I(N__6567));
    Sp12to4 I__1644 (
            .O(N__6567),
            .I(N__6564));
    Odrv12 I__1643 (
            .O(N__6564),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1642 (
            .O(N__6561),
            .I(N__6558));
    LocalMux I__1641 (
            .O(N__6558),
            .I(N__6555));
    IoSpan4Mux I__1640 (
            .O(N__6555),
            .I(N__6552));
    IoSpan4Mux I__1639 (
            .O(N__6552),
            .I(N__6549));
    Sp12to4 I__1638 (
            .O(N__6549),
            .I(N__6546));
    Span12Mux_s6_v I__1637 (
            .O(N__6546),
            .I(N__6543));
    Odrv12 I__1636 (
            .O(N__6543),
            .I(un1_D_UU_AMIGA_5));
    CascadeMux I__1635 (
            .O(N__6540),
            .I(N__6537));
    InMux I__1634 (
            .O(N__6537),
            .I(N__6534));
    LocalMux I__1633 (
            .O(N__6534),
            .I(N__6530));
    InMux I__1632 (
            .O(N__6533),
            .I(N__6527));
    Span4Mux_v I__1631 (
            .O(N__6530),
            .I(N__6523));
    LocalMux I__1630 (
            .O(N__6527),
            .I(N__6520));
    InMux I__1629 (
            .O(N__6526),
            .I(N__6517));
    Span4Mux_v I__1628 (
            .O(N__6523),
            .I(N__6514));
    Span4Mux_v I__1627 (
            .O(N__6520),
            .I(N__6509));
    LocalMux I__1626 (
            .O(N__6517),
            .I(N__6509));
    Span4Mux_v I__1625 (
            .O(N__6514),
            .I(N__6504));
    Span4Mux_v I__1624 (
            .O(N__6509),
            .I(N__6504));
    Sp12to4 I__1623 (
            .O(N__6504),
            .I(N__6501));
    Span12Mux_h I__1622 (
            .O(N__6501),
            .I(N__6498));
    Odrv12 I__1621 (
            .O(N__6498),
            .I(D_UU_AMIGA_in_3));
    InMux I__1620 (
            .O(N__6495),
            .I(N__6492));
    LocalMux I__1619 (
            .O(N__6492),
            .I(N__6489));
    Odrv12 I__1618 (
            .O(N__6489),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    IoInMux I__1617 (
            .O(N__6486),
            .I(N__6483));
    LocalMux I__1616 (
            .O(N__6483),
            .I(N__6480));
    Span4Mux_s2_v I__1615 (
            .O(N__6480),
            .I(N__6477));
    Span4Mux_h I__1614 (
            .O(N__6477),
            .I(N__6474));
    Span4Mux_v I__1613 (
            .O(N__6474),
            .I(N__6471));
    Sp12to4 I__1612 (
            .O(N__6471),
            .I(N__6468));
    Odrv12 I__1611 (
            .O(N__6468),
            .I(un1_D_UU_AMIGA_3));
    IoInMux I__1610 (
            .O(N__6465),
            .I(N__6462));
    LocalMux I__1609 (
            .O(N__6462),
            .I(N__6459));
    IoSpan4Mux I__1608 (
            .O(N__6459),
            .I(N__6456));
    Span4Mux_s2_h I__1607 (
            .O(N__6456),
            .I(N__6453));
    Sp12to4 I__1606 (
            .O(N__6453),
            .I(N__6450));
    Odrv12 I__1605 (
            .O(N__6450),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1604 (
            .O(N__6447),
            .I(N__6442));
    InMux I__1603 (
            .O(N__6446),
            .I(N__6439));
    CascadeMux I__1602 (
            .O(N__6445),
            .I(N__6436));
    LocalMux I__1601 (
            .O(N__6442),
            .I(N__6431));
    LocalMux I__1600 (
            .O(N__6439),
            .I(N__6431));
    InMux I__1599 (
            .O(N__6436),
            .I(N__6428));
    Span4Mux_v I__1598 (
            .O(N__6431),
            .I(N__6425));
    LocalMux I__1597 (
            .O(N__6428),
            .I(N__6422));
    Sp12to4 I__1596 (
            .O(N__6425),
            .I(N__6419));
    Span12Mux_v I__1595 (
            .O(N__6422),
            .I(N__6416));
    Span12Mux_h I__1594 (
            .O(N__6419),
            .I(N__6413));
    Odrv12 I__1593 (
            .O(N__6416),
            .I(D_UM_AMIGA_in_2));
    Odrv12 I__1592 (
            .O(N__6413),
            .I(D_UM_AMIGA_in_2));
    InMux I__1591 (
            .O(N__6408),
            .I(N__6405));
    LocalMux I__1590 (
            .O(N__6405),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    CascadeMux I__1589 (
            .O(N__6402),
            .I(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ));
    InMux I__1588 (
            .O(N__6399),
            .I(N__6395));
    CascadeMux I__1587 (
            .O(N__6398),
            .I(N__6389));
    LocalMux I__1586 (
            .O(N__6395),
            .I(N__6382));
    InMux I__1585 (
            .O(N__6394),
            .I(N__6377));
    InMux I__1584 (
            .O(N__6393),
            .I(N__6377));
    InMux I__1583 (
            .O(N__6392),
            .I(N__6374));
    InMux I__1582 (
            .O(N__6389),
            .I(N__6369));
    InMux I__1581 (
            .O(N__6388),
            .I(N__6369));
    InMux I__1580 (
            .O(N__6387),
            .I(N__6362));
    InMux I__1579 (
            .O(N__6386),
            .I(N__6362));
    InMux I__1578 (
            .O(N__6385),
            .I(N__6362));
    Odrv4 I__1577 (
            .O(N__6382),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1576 (
            .O(N__6377),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1575 (
            .O(N__6374),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1574 (
            .O(N__6369),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1573 (
            .O(N__6362),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    CascadeMux I__1572 (
            .O(N__6351),
            .I(N__6347));
    CascadeMux I__1571 (
            .O(N__6350),
            .I(N__6343));
    InMux I__1570 (
            .O(N__6347),
            .I(N__6336));
    InMux I__1569 (
            .O(N__6346),
            .I(N__6336));
    InMux I__1568 (
            .O(N__6343),
            .I(N__6331));
    InMux I__1567 (
            .O(N__6342),
            .I(N__6331));
    InMux I__1566 (
            .O(N__6341),
            .I(N__6328));
    LocalMux I__1565 (
            .O(N__6336),
            .I(N__6323));
    LocalMux I__1564 (
            .O(N__6331),
            .I(N__6323));
    LocalMux I__1563 (
            .O(N__6328),
            .I(N__6320));
    Span4Mux_v I__1562 (
            .O(N__6323),
            .I(N__6317));
    Span4Mux_h I__1561 (
            .O(N__6320),
            .I(N__6314));
    Sp12to4 I__1560 (
            .O(N__6317),
            .I(N__6311));
    Span4Mux_v I__1559 (
            .O(N__6314),
            .I(N__6308));
    Span12Mux_h I__1558 (
            .O(N__6311),
            .I(N__6305));
    Span4Mux_v I__1557 (
            .O(N__6308),
            .I(N__6302));
    Span12Mux_v I__1556 (
            .O(N__6305),
            .I(N__6299));
    Span4Mux_v I__1555 (
            .O(N__6302),
            .I(N__6296));
    Odrv12 I__1554 (
            .O(N__6299),
            .I(TACKn_c));
    Odrv4 I__1553 (
            .O(N__6296),
            .I(TACKn_c));
    InMux I__1552 (
            .O(N__6291),
            .I(N__6285));
    CascadeMux I__1551 (
            .O(N__6290),
            .I(N__6277));
    InMux I__1550 (
            .O(N__6289),
            .I(N__6272));
    InMux I__1549 (
            .O(N__6288),
            .I(N__6272));
    LocalMux I__1548 (
            .O(N__6285),
            .I(N__6269));
    InMux I__1547 (
            .O(N__6284),
            .I(N__6266));
    InMux I__1546 (
            .O(N__6283),
            .I(N__6261));
    InMux I__1545 (
            .O(N__6282),
            .I(N__6261));
    InMux I__1544 (
            .O(N__6281),
            .I(N__6254));
    InMux I__1543 (
            .O(N__6280),
            .I(N__6254));
    InMux I__1542 (
            .O(N__6277),
            .I(N__6254));
    LocalMux I__1541 (
            .O(N__6272),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv4 I__1540 (
            .O(N__6269),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1539 (
            .O(N__6266),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1538 (
            .O(N__6261),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1537 (
            .O(N__6254),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1536 (
            .O(N__6243),
            .I(N__6240));
    LocalMux I__1535 (
            .O(N__6240),
            .I(\U111_CYCLE_SM.LW_CYCLE_0 ));
    InMux I__1534 (
            .O(N__6237),
            .I(N__6234));
    LocalMux I__1533 (
            .O(N__6234),
            .I(N__6221));
    ClkMux I__1532 (
            .O(N__6233),
            .I(N__6198));
    ClkMux I__1531 (
            .O(N__6232),
            .I(N__6198));
    ClkMux I__1530 (
            .O(N__6231),
            .I(N__6198));
    ClkMux I__1529 (
            .O(N__6230),
            .I(N__6198));
    ClkMux I__1528 (
            .O(N__6229),
            .I(N__6198));
    ClkMux I__1527 (
            .O(N__6228),
            .I(N__6198));
    ClkMux I__1526 (
            .O(N__6227),
            .I(N__6198));
    ClkMux I__1525 (
            .O(N__6226),
            .I(N__6198));
    ClkMux I__1524 (
            .O(N__6225),
            .I(N__6198));
    ClkMux I__1523 (
            .O(N__6224),
            .I(N__6198));
    Glb2LocalMux I__1522 (
            .O(N__6221),
            .I(N__6198));
    GlobalMux I__1521 (
            .O(N__6198),
            .I(CLK80));
    IoInMux I__1520 (
            .O(N__6195),
            .I(N__6192));
    LocalMux I__1519 (
            .O(N__6192),
            .I(N__6189));
    IoSpan4Mux I__1518 (
            .O(N__6189),
            .I(N__6184));
    IoInMux I__1517 (
            .O(N__6188),
            .I(N__6181));
    IoInMux I__1516 (
            .O(N__6187),
            .I(N__6178));
    IoSpan4Mux I__1515 (
            .O(N__6184),
            .I(N__6173));
    LocalMux I__1514 (
            .O(N__6181),
            .I(N__6173));
    LocalMux I__1513 (
            .O(N__6178),
            .I(N__6170));
    IoSpan4Mux I__1512 (
            .O(N__6173),
            .I(N__6167));
    IoSpan4Mux I__1511 (
            .O(N__6170),
            .I(N__6164));
    Span4Mux_s2_v I__1510 (
            .O(N__6167),
            .I(N__6161));
    Span4Mux_s2_h I__1509 (
            .O(N__6164),
            .I(N__6158));
    Sp12to4 I__1508 (
            .O(N__6161),
            .I(N__6155));
    Sp12to4 I__1507 (
            .O(N__6158),
            .I(N__6152));
    Span12Mux_s9_v I__1506 (
            .O(N__6155),
            .I(N__6149));
    Span12Mux_h I__1505 (
            .O(N__6152),
            .I(N__6146));
    Odrv12 I__1504 (
            .O(N__6149),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1503 (
            .O(N__6146),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1502 (
            .O(N__6141),
            .I(N__6138));
    LocalMux I__1501 (
            .O(N__6138),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    CascadeMux I__1500 (
            .O(N__6135),
            .I(N__6132));
    InMux I__1499 (
            .O(N__6132),
            .I(N__6129));
    LocalMux I__1498 (
            .O(N__6129),
            .I(N__6124));
    InMux I__1497 (
            .O(N__6128),
            .I(N__6121));
    InMux I__1496 (
            .O(N__6127),
            .I(N__6118));
    Span4Mux_v I__1495 (
            .O(N__6124),
            .I(N__6115));
    LocalMux I__1494 (
            .O(N__6121),
            .I(N__6110));
    LocalMux I__1493 (
            .O(N__6118),
            .I(N__6110));
    Sp12to4 I__1492 (
            .O(N__6115),
            .I(N__6107));
    Span4Mux_v I__1491 (
            .O(N__6110),
            .I(N__6104));
    Span12Mux_h I__1490 (
            .O(N__6107),
            .I(N__6101));
    Sp12to4 I__1489 (
            .O(N__6104),
            .I(N__6098));
    Span12Mux_v I__1488 (
            .O(N__6101),
            .I(N__6093));
    Span12Mux_h I__1487 (
            .O(N__6098),
            .I(N__6093));
    Odrv12 I__1486 (
            .O(N__6093),
            .I(D_UM_AMIGA_in_1));
    InMux I__1485 (
            .O(N__6090),
            .I(N__6084));
    InMux I__1484 (
            .O(N__6089),
            .I(N__6081));
    InMux I__1483 (
            .O(N__6088),
            .I(N__6076));
    InMux I__1482 (
            .O(N__6087),
            .I(N__6076));
    LocalMux I__1481 (
            .O(N__6084),
            .I(N__6072));
    LocalMux I__1480 (
            .O(N__6081),
            .I(N__6069));
    LocalMux I__1479 (
            .O(N__6076),
            .I(N__6066));
    ClkMux I__1478 (
            .O(N__6075),
            .I(N__6057));
    Glb2LocalMux I__1477 (
            .O(N__6072),
            .I(N__6057));
    Glb2LocalMux I__1476 (
            .O(N__6069),
            .I(N__6057));
    Glb2LocalMux I__1475 (
            .O(N__6066),
            .I(N__6057));
    GlobalMux I__1474 (
            .O(N__6057),
            .I(CLK40));
    CascadeMux I__1473 (
            .O(N__6054),
            .I(\U111_CYCLE_SM.N_91_cascade_ ));
    InMux I__1472 (
            .O(N__6051),
            .I(N__6048));
    LocalMux I__1471 (
            .O(N__6048),
            .I(N__6045));
    Span4Mux_v I__1470 (
            .O(N__6045),
            .I(N__6042));
    Span4Mux_v I__1469 (
            .O(N__6042),
            .I(N__6037));
    InMux I__1468 (
            .O(N__6041),
            .I(N__6034));
    InMux I__1467 (
            .O(N__6040),
            .I(N__6031));
    Sp12to4 I__1466 (
            .O(N__6037),
            .I(N__6024));
    LocalMux I__1465 (
            .O(N__6034),
            .I(N__6024));
    LocalMux I__1464 (
            .O(N__6031),
            .I(N__6024));
    Span12Mux_h I__1463 (
            .O(N__6024),
            .I(N__6021));
    Span12Mux_v I__1462 (
            .O(N__6021),
            .I(N__6018));
    Odrv12 I__1461 (
            .O(N__6018),
            .I(D_UM_AMIGA_in_6));
    InMux I__1460 (
            .O(N__6015),
            .I(N__6012));
    LocalMux I__1459 (
            .O(N__6012),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    IoInMux I__1458 (
            .O(N__6009),
            .I(N__6006));
    LocalMux I__1457 (
            .O(N__6006),
            .I(N__6003));
    Span4Mux_s3_h I__1456 (
            .O(N__6003),
            .I(N__6000));
    Span4Mux_h I__1455 (
            .O(N__6000),
            .I(N__5997));
    Span4Mux_h I__1454 (
            .O(N__5997),
            .I(N__5994));
    Span4Mux_h I__1453 (
            .O(N__5994),
            .I(N__5991));
    Odrv4 I__1452 (
            .O(N__5991),
            .I(un1_D_UM_AMIGA_6));
    CascadeMux I__1451 (
            .O(N__5988),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ));
    IoInMux I__1450 (
            .O(N__5985),
            .I(N__5978));
    IoInMux I__1449 (
            .O(N__5984),
            .I(N__5975));
    IoInMux I__1448 (
            .O(N__5983),
            .I(N__5972));
    IoInMux I__1447 (
            .O(N__5982),
            .I(N__5969));
    InMux I__1446 (
            .O(N__5981),
            .I(N__5964));
    LocalMux I__1445 (
            .O(N__5978),
            .I(N__5955));
    LocalMux I__1444 (
            .O(N__5975),
            .I(N__5955));
    LocalMux I__1443 (
            .O(N__5972),
            .I(N__5955));
    LocalMux I__1442 (
            .O(N__5969),
            .I(N__5955));
    IoInMux I__1441 (
            .O(N__5968),
            .I(N__5952));
    IoInMux I__1440 (
            .O(N__5967),
            .I(N__5943));
    LocalMux I__1439 (
            .O(N__5964),
            .I(N__5940));
    IoSpan4Mux I__1438 (
            .O(N__5955),
            .I(N__5930));
    LocalMux I__1437 (
            .O(N__5952),
            .I(N__5930));
    IoInMux I__1436 (
            .O(N__5951),
            .I(N__5927));
    IoInMux I__1435 (
            .O(N__5950),
            .I(N__5924));
    IoInMux I__1434 (
            .O(N__5949),
            .I(N__5921));
    IoInMux I__1433 (
            .O(N__5948),
            .I(N__5918));
    IoInMux I__1432 (
            .O(N__5947),
            .I(N__5915));
    IoInMux I__1431 (
            .O(N__5946),
            .I(N__5912));
    LocalMux I__1430 (
            .O(N__5943),
            .I(N__5908));
    Span4Mux_h I__1429 (
            .O(N__5940),
            .I(N__5905));
    IoInMux I__1428 (
            .O(N__5939),
            .I(N__5901));
    IoInMux I__1427 (
            .O(N__5938),
            .I(N__5898));
    IoInMux I__1426 (
            .O(N__5937),
            .I(N__5895));
    IoInMux I__1425 (
            .O(N__5936),
            .I(N__5892));
    IoInMux I__1424 (
            .O(N__5935),
            .I(N__5889));
    IoSpan4Mux I__1423 (
            .O(N__5930),
            .I(N__5870));
    LocalMux I__1422 (
            .O(N__5927),
            .I(N__5870));
    LocalMux I__1421 (
            .O(N__5924),
            .I(N__5870));
    LocalMux I__1420 (
            .O(N__5921),
            .I(N__5870));
    LocalMux I__1419 (
            .O(N__5918),
            .I(N__5870));
    LocalMux I__1418 (
            .O(N__5915),
            .I(N__5870));
    LocalMux I__1417 (
            .O(N__5912),
            .I(N__5870));
    IoInMux I__1416 (
            .O(N__5911),
            .I(N__5867));
    Span4Mux_s3_v I__1415 (
            .O(N__5908),
            .I(N__5863));
    Span4Mux_v I__1414 (
            .O(N__5905),
            .I(N__5860));
    InMux I__1413 (
            .O(N__5904),
            .I(N__5857));
    LocalMux I__1412 (
            .O(N__5901),
            .I(N__5846));
    LocalMux I__1411 (
            .O(N__5898),
            .I(N__5846));
    LocalMux I__1410 (
            .O(N__5895),
            .I(N__5846));
    LocalMux I__1409 (
            .O(N__5892),
            .I(N__5846));
    LocalMux I__1408 (
            .O(N__5889),
            .I(N__5846));
    IoInMux I__1407 (
            .O(N__5888),
            .I(N__5843));
    IoInMux I__1406 (
            .O(N__5887),
            .I(N__5840));
    IoInMux I__1405 (
            .O(N__5886),
            .I(N__5837));
    IoInMux I__1404 (
            .O(N__5885),
            .I(N__5834));
    IoSpan4Mux I__1403 (
            .O(N__5870),
            .I(N__5825));
    LocalMux I__1402 (
            .O(N__5867),
            .I(N__5825));
    IoInMux I__1401 (
            .O(N__5866),
            .I(N__5822));
    Span4Mux_v I__1400 (
            .O(N__5863),
            .I(N__5817));
    Span4Mux_h I__1399 (
            .O(N__5860),
            .I(N__5812));
    LocalMux I__1398 (
            .O(N__5857),
            .I(N__5812));
    IoSpan4Mux I__1397 (
            .O(N__5846),
            .I(N__5801));
    LocalMux I__1396 (
            .O(N__5843),
            .I(N__5801));
    LocalMux I__1395 (
            .O(N__5840),
            .I(N__5801));
    LocalMux I__1394 (
            .O(N__5837),
            .I(N__5801));
    LocalMux I__1393 (
            .O(N__5834),
            .I(N__5801));
    IoInMux I__1392 (
            .O(N__5833),
            .I(N__5798));
    IoInMux I__1391 (
            .O(N__5832),
            .I(N__5795));
    IoInMux I__1390 (
            .O(N__5831),
            .I(N__5792));
    IoInMux I__1389 (
            .O(N__5830),
            .I(N__5789));
    IoSpan4Mux I__1388 (
            .O(N__5825),
            .I(N__5784));
    LocalMux I__1387 (
            .O(N__5822),
            .I(N__5784));
    IoInMux I__1386 (
            .O(N__5821),
            .I(N__5781));
    IoInMux I__1385 (
            .O(N__5820),
            .I(N__5778));
    Span4Mux_v I__1384 (
            .O(N__5817),
            .I(N__5774));
    Span4Mux_v I__1383 (
            .O(N__5812),
            .I(N__5771));
    IoSpan4Mux I__1382 (
            .O(N__5801),
            .I(N__5760));
    LocalMux I__1381 (
            .O(N__5798),
            .I(N__5760));
    LocalMux I__1380 (
            .O(N__5795),
            .I(N__5760));
    LocalMux I__1379 (
            .O(N__5792),
            .I(N__5760));
    LocalMux I__1378 (
            .O(N__5789),
            .I(N__5760));
    IoSpan4Mux I__1377 (
            .O(N__5784),
            .I(N__5753));
    LocalMux I__1376 (
            .O(N__5781),
            .I(N__5753));
    LocalMux I__1375 (
            .O(N__5778),
            .I(N__5753));
    IoInMux I__1374 (
            .O(N__5777),
            .I(N__5750));
    Sp12to4 I__1373 (
            .O(N__5774),
            .I(N__5745));
    Sp12to4 I__1372 (
            .O(N__5771),
            .I(N__5741));
    IoSpan4Mux I__1371 (
            .O(N__5760),
            .I(N__5738));
    IoSpan4Mux I__1370 (
            .O(N__5753),
            .I(N__5733));
    LocalMux I__1369 (
            .O(N__5750),
            .I(N__5733));
    IoInMux I__1368 (
            .O(N__5749),
            .I(N__5730));
    IoInMux I__1367 (
            .O(N__5748),
            .I(N__5727));
    Span12Mux_h I__1366 (
            .O(N__5745),
            .I(N__5724));
    IoInMux I__1365 (
            .O(N__5744),
            .I(N__5721));
    Span12Mux_h I__1364 (
            .O(N__5741),
            .I(N__5718));
    IoSpan4Mux I__1363 (
            .O(N__5738),
            .I(N__5713));
    IoSpan4Mux I__1362 (
            .O(N__5733),
            .I(N__5713));
    LocalMux I__1361 (
            .O(N__5730),
            .I(N__5710));
    LocalMux I__1360 (
            .O(N__5727),
            .I(N__5707));
    Span12Mux_h I__1359 (
            .O(N__5724),
            .I(N__5702));
    LocalMux I__1358 (
            .O(N__5721),
            .I(N__5702));
    Odrv12 I__1357 (
            .O(N__5718),
            .I(RnW_c));
    Odrv4 I__1356 (
            .O(N__5713),
            .I(RnW_c));
    Odrv4 I__1355 (
            .O(N__5710),
            .I(RnW_c));
    Odrv4 I__1354 (
            .O(N__5707),
            .I(RnW_c));
    Odrv12 I__1353 (
            .O(N__5702),
            .I(RnW_c));
    CascadeMux I__1352 (
            .O(N__5691),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ));
    InMux I__1351 (
            .O(N__5688),
            .I(N__5685));
    LocalMux I__1350 (
            .O(N__5685),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ));
    CascadeMux I__1349 (
            .O(N__5682),
            .I(N__5675));
    InMux I__1348 (
            .O(N__5681),
            .I(N__5672));
    InMux I__1347 (
            .O(N__5680),
            .I(N__5669));
    InMux I__1346 (
            .O(N__5679),
            .I(N__5666));
    InMux I__1345 (
            .O(N__5678),
            .I(N__5663));
    InMux I__1344 (
            .O(N__5675),
            .I(N__5660));
    LocalMux I__1343 (
            .O(N__5672),
            .I(N__5657));
    LocalMux I__1342 (
            .O(N__5669),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1341 (
            .O(N__5666),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1340 (
            .O(N__5663),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    LocalMux I__1339 (
            .O(N__5660),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    Odrv4 I__1338 (
            .O(N__5657),
            .I(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ));
    InMux I__1337 (
            .O(N__5646),
            .I(N__5640));
    InMux I__1336 (
            .O(N__5645),
            .I(N__5637));
    CascadeMux I__1335 (
            .O(N__5644),
            .I(N__5632));
    InMux I__1334 (
            .O(N__5643),
            .I(N__5628));
    LocalMux I__1333 (
            .O(N__5640),
            .I(N__5623));
    LocalMux I__1332 (
            .O(N__5637),
            .I(N__5623));
    InMux I__1331 (
            .O(N__5636),
            .I(N__5618));
    InMux I__1330 (
            .O(N__5635),
            .I(N__5618));
    InMux I__1329 (
            .O(N__5632),
            .I(N__5613));
    InMux I__1328 (
            .O(N__5631),
            .I(N__5613));
    LocalMux I__1327 (
            .O(N__5628),
            .I(N__5610));
    Span4Mux_v I__1326 (
            .O(N__5623),
            .I(N__5602));
    LocalMux I__1325 (
            .O(N__5618),
            .I(N__5602));
    LocalMux I__1324 (
            .O(N__5613),
            .I(N__5602));
    Span4Mux_v I__1323 (
            .O(N__5610),
            .I(N__5598));
    InMux I__1322 (
            .O(N__5609),
            .I(N__5595));
    Span4Mux_v I__1321 (
            .O(N__5602),
            .I(N__5592));
    InMux I__1320 (
            .O(N__5601),
            .I(N__5589));
    Sp12to4 I__1319 (
            .O(N__5598),
            .I(N__5584));
    LocalMux I__1318 (
            .O(N__5595),
            .I(N__5584));
    Span4Mux_h I__1317 (
            .O(N__5592),
            .I(N__5581));
    LocalMux I__1316 (
            .O(N__5589),
            .I(N__5578));
    Span12Mux_h I__1315 (
            .O(N__5584),
            .I(N__5575));
    Sp12to4 I__1314 (
            .O(N__5581),
            .I(N__5572));
    Span4Mux_v I__1313 (
            .O(N__5578),
            .I(N__5569));
    Span12Mux_v I__1312 (
            .O(N__5575),
            .I(N__5566));
    Span12Mux_v I__1311 (
            .O(N__5572),
            .I(N__5561));
    Sp12to4 I__1310 (
            .O(N__5569),
            .I(N__5561));
    Odrv12 I__1309 (
            .O(N__5566),
            .I(RESETn_c));
    Odrv12 I__1308 (
            .O(N__5561),
            .I(RESETn_c));
    InMux I__1307 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__1306 (
            .O(N__5553),
            .I(N__5550));
    Span4Mux_v I__1305 (
            .O(N__5550),
            .I(N__5547));
    Odrv4 I__1304 (
            .O(N__5547),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    CascadeMux I__1303 (
            .O(N__5544),
            .I(N__5541));
    InMux I__1302 (
            .O(N__5541),
            .I(N__5537));
    InMux I__1301 (
            .O(N__5540),
            .I(N__5534));
    LocalMux I__1300 (
            .O(N__5537),
            .I(N__5531));
    LocalMux I__1299 (
            .O(N__5534),
            .I(N__5528));
    Span4Mux_v I__1298 (
            .O(N__5531),
            .I(N__5524));
    Span4Mux_v I__1297 (
            .O(N__5528),
            .I(N__5521));
    InMux I__1296 (
            .O(N__5527),
            .I(N__5518));
    Span4Mux_v I__1295 (
            .O(N__5524),
            .I(N__5515));
    Span4Mux_v I__1294 (
            .O(N__5521),
            .I(N__5510));
    LocalMux I__1293 (
            .O(N__5518),
            .I(N__5510));
    Span4Mux_v I__1292 (
            .O(N__5515),
            .I(N__5507));
    Span4Mux_v I__1291 (
            .O(N__5510),
            .I(N__5504));
    Sp12to4 I__1290 (
            .O(N__5507),
            .I(N__5499));
    Sp12to4 I__1289 (
            .O(N__5504),
            .I(N__5499));
    Span12Mux_h I__1288 (
            .O(N__5499),
            .I(N__5496));
    Odrv12 I__1287 (
            .O(N__5496),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1286 (
            .O(N__5493),
            .I(N__5490));
    LocalMux I__1285 (
            .O(N__5490),
            .I(N__5487));
    Span12Mux_s11_v I__1284 (
            .O(N__5487),
            .I(N__5484));
    Span12Mux_h I__1283 (
            .O(N__5484),
            .I(N__5481));
    Odrv12 I__1282 (
            .O(N__5481),
            .I(un1_D_UU_AMIGA_2));
    IoInMux I__1281 (
            .O(N__5478),
            .I(N__5473));
    IoInMux I__1280 (
            .O(N__5477),
            .I(N__5470));
    IoInMux I__1279 (
            .O(N__5476),
            .I(N__5467));
    LocalMux I__1278 (
            .O(N__5473),
            .I(N__5464));
    LocalMux I__1277 (
            .O(N__5470),
            .I(N__5461));
    LocalMux I__1276 (
            .O(N__5467),
            .I(N__5458));
    Span12Mux_s4_v I__1275 (
            .O(N__5464),
            .I(N__5455));
    Span12Mux_s9_h I__1274 (
            .O(N__5461),
            .I(N__5450));
    Span12Mux_s10_h I__1273 (
            .O(N__5458),
            .I(N__5450));
    Odrv12 I__1272 (
            .O(N__5455),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__1271 (
            .O(N__5450),
            .I(GB_BUFFER_CLK40_THRU_CO));
    CascadeMux I__1270 (
            .O(N__5445),
            .I(N__5441));
    InMux I__1269 (
            .O(N__5444),
            .I(N__5438));
    InMux I__1268 (
            .O(N__5441),
            .I(N__5435));
    LocalMux I__1267 (
            .O(N__5438),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    LocalMux I__1266 (
            .O(N__5435),
            .I(\U111_CYCLE_SM.TA_ENZ0 ));
    IoInMux I__1265 (
            .O(N__5430),
            .I(N__5426));
    IoInMux I__1264 (
            .O(N__5429),
            .I(N__5423));
    LocalMux I__1263 (
            .O(N__5426),
            .I(N__5420));
    LocalMux I__1262 (
            .O(N__5423),
            .I(N__5417));
    Span4Mux_s3_v I__1261 (
            .O(N__5420),
            .I(N__5414));
    Span4Mux_s2_v I__1260 (
            .O(N__5417),
            .I(N__5411));
    Sp12to4 I__1259 (
            .O(N__5414),
            .I(N__5408));
    Span4Mux_h I__1258 (
            .O(N__5411),
            .I(N__5405));
    Span12Mux_s11_h I__1257 (
            .O(N__5408),
            .I(N__5402));
    Span4Mux_v I__1256 (
            .O(N__5405),
            .I(N__5399));
    Span12Mux_v I__1255 (
            .O(N__5402),
            .I(N__5396));
    Sp12to4 I__1254 (
            .O(N__5399),
            .I(N__5393));
    Odrv12 I__1253 (
            .O(N__5396),
            .I(U111_CYCLE_SM_TAn_0_i));
    Odrv12 I__1252 (
            .O(N__5393),
            .I(U111_CYCLE_SM_TAn_0_i));
    InMux I__1251 (
            .O(N__5388),
            .I(N__5381));
    InMux I__1250 (
            .O(N__5387),
            .I(N__5381));
    InMux I__1249 (
            .O(N__5386),
            .I(N__5375));
    LocalMux I__1248 (
            .O(N__5381),
            .I(N__5369));
    InMux I__1247 (
            .O(N__5380),
            .I(N__5363));
    InMux I__1246 (
            .O(N__5379),
            .I(N__5360));
    InMux I__1245 (
            .O(N__5378),
            .I(N__5357));
    LocalMux I__1244 (
            .O(N__5375),
            .I(N__5353));
    InMux I__1243 (
            .O(N__5374),
            .I(N__5349));
    InMux I__1242 (
            .O(N__5373),
            .I(N__5345));
    InMux I__1241 (
            .O(N__5372),
            .I(N__5334));
    Span4Mux_h I__1240 (
            .O(N__5369),
            .I(N__5331));
    InMux I__1239 (
            .O(N__5368),
            .I(N__5328));
    InMux I__1238 (
            .O(N__5367),
            .I(N__5323));
    InMux I__1237 (
            .O(N__5366),
            .I(N__5323));
    LocalMux I__1236 (
            .O(N__5363),
            .I(N__5318));
    LocalMux I__1235 (
            .O(N__5360),
            .I(N__5313));
    LocalMux I__1234 (
            .O(N__5357),
            .I(N__5313));
    InMux I__1233 (
            .O(N__5356),
            .I(N__5310));
    Span4Mux_h I__1232 (
            .O(N__5353),
            .I(N__5304));
    InMux I__1231 (
            .O(N__5352),
            .I(N__5301));
    LocalMux I__1230 (
            .O(N__5349),
            .I(N__5298));
    InMux I__1229 (
            .O(N__5348),
            .I(N__5295));
    LocalMux I__1228 (
            .O(N__5345),
            .I(N__5292));
    InMux I__1227 (
            .O(N__5344),
            .I(N__5289));
    InMux I__1226 (
            .O(N__5343),
            .I(N__5286));
    InMux I__1225 (
            .O(N__5342),
            .I(N__5281));
    InMux I__1224 (
            .O(N__5341),
            .I(N__5281));
    InMux I__1223 (
            .O(N__5340),
            .I(N__5276));
    InMux I__1222 (
            .O(N__5339),
            .I(N__5276));
    InMux I__1221 (
            .O(N__5338),
            .I(N__5272));
    InMux I__1220 (
            .O(N__5337),
            .I(N__5269));
    LocalMux I__1219 (
            .O(N__5334),
            .I(N__5265));
    Span4Mux_v I__1218 (
            .O(N__5331),
            .I(N__5262));
    LocalMux I__1217 (
            .O(N__5328),
            .I(N__5259));
    LocalMux I__1216 (
            .O(N__5323),
            .I(N__5256));
    InMux I__1215 (
            .O(N__5322),
            .I(N__5251));
    InMux I__1214 (
            .O(N__5321),
            .I(N__5251));
    Span4Mux_h I__1213 (
            .O(N__5318),
            .I(N__5246));
    Span4Mux_v I__1212 (
            .O(N__5313),
            .I(N__5246));
    LocalMux I__1211 (
            .O(N__5310),
            .I(N__5243));
    InMux I__1210 (
            .O(N__5309),
            .I(N__5240));
    InMux I__1209 (
            .O(N__5308),
            .I(N__5237));
    InMux I__1208 (
            .O(N__5307),
            .I(N__5234));
    Span4Mux_v I__1207 (
            .O(N__5304),
            .I(N__5229));
    LocalMux I__1206 (
            .O(N__5301),
            .I(N__5229));
    Span4Mux_v I__1205 (
            .O(N__5298),
            .I(N__5223));
    LocalMux I__1204 (
            .O(N__5295),
            .I(N__5223));
    Span4Mux_v I__1203 (
            .O(N__5292),
            .I(N__5216));
    LocalMux I__1202 (
            .O(N__5289),
            .I(N__5216));
    LocalMux I__1201 (
            .O(N__5286),
            .I(N__5216));
    LocalMux I__1200 (
            .O(N__5281),
            .I(N__5211));
    LocalMux I__1199 (
            .O(N__5276),
            .I(N__5211));
    InMux I__1198 (
            .O(N__5275),
            .I(N__5208));
    LocalMux I__1197 (
            .O(N__5272),
            .I(N__5205));
    LocalMux I__1196 (
            .O(N__5269),
            .I(N__5202));
    InMux I__1195 (
            .O(N__5268),
            .I(N__5199));
    Span4Mux_h I__1194 (
            .O(N__5265),
            .I(N__5195));
    Span4Mux_v I__1193 (
            .O(N__5262),
            .I(N__5190));
    Span4Mux_h I__1192 (
            .O(N__5259),
            .I(N__5190));
    Span4Mux_v I__1191 (
            .O(N__5256),
            .I(N__5185));
    LocalMux I__1190 (
            .O(N__5251),
            .I(N__5185));
    Span4Mux_v I__1189 (
            .O(N__5246),
            .I(N__5174));
    Span4Mux_h I__1188 (
            .O(N__5243),
            .I(N__5174));
    LocalMux I__1187 (
            .O(N__5240),
            .I(N__5174));
    LocalMux I__1186 (
            .O(N__5237),
            .I(N__5174));
    LocalMux I__1185 (
            .O(N__5234),
            .I(N__5174));
    Span4Mux_v I__1184 (
            .O(N__5229),
            .I(N__5171));
    InMux I__1183 (
            .O(N__5228),
            .I(N__5168));
    Span4Mux_h I__1182 (
            .O(N__5223),
            .I(N__5165));
    Span4Mux_h I__1181 (
            .O(N__5216),
            .I(N__5158));
    Span4Mux_v I__1180 (
            .O(N__5211),
            .I(N__5158));
    LocalMux I__1179 (
            .O(N__5208),
            .I(N__5158));
    Span4Mux_v I__1178 (
            .O(N__5205),
            .I(N__5151));
    Span4Mux_h I__1177 (
            .O(N__5202),
            .I(N__5151));
    LocalMux I__1176 (
            .O(N__5199),
            .I(N__5151));
    InMux I__1175 (
            .O(N__5198),
            .I(N__5148));
    Sp12to4 I__1174 (
            .O(N__5195),
            .I(N__5145));
    Span4Mux_h I__1173 (
            .O(N__5190),
            .I(N__5140));
    Span4Mux_v I__1172 (
            .O(N__5185),
            .I(N__5140));
    Span4Mux_v I__1171 (
            .O(N__5174),
            .I(N__5137));
    Sp12to4 I__1170 (
            .O(N__5171),
            .I(N__5132));
    LocalMux I__1169 (
            .O(N__5168),
            .I(N__5132));
    Span4Mux_v I__1168 (
            .O(N__5165),
            .I(N__5123));
    Span4Mux_v I__1167 (
            .O(N__5158),
            .I(N__5123));
    Span4Mux_h I__1166 (
            .O(N__5151),
            .I(N__5123));
    LocalMux I__1165 (
            .O(N__5148),
            .I(N__5123));
    Odrv12 I__1164 (
            .O(N__5145),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1163 (
            .O(N__5140),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1162 (
            .O(N__5137),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv12 I__1161 (
            .O(N__5132),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    Odrv4 I__1160 (
            .O(N__5123),
            .I(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ));
    InMux I__1159 (
            .O(N__5112),
            .I(N__5106));
    InMux I__1158 (
            .O(N__5111),
            .I(N__5106));
    LocalMux I__1157 (
            .O(N__5106),
            .I(N__5103));
    Span12Mux_h I__1156 (
            .O(N__5103),
            .I(N__5100));
    Span12Mux_v I__1155 (
            .O(N__5100),
            .I(N__5097));
    Odrv12 I__1154 (
            .O(N__5097),
            .I(PORTSIZE_c));
    InMux I__1153 (
            .O(N__5094),
            .I(N__5088));
    InMux I__1152 (
            .O(N__5093),
            .I(N__5088));
    LocalMux I__1151 (
            .O(N__5088),
            .I(N__5085));
    Span12Mux_h I__1150 (
            .O(N__5085),
            .I(N__5082));
    Span12Mux_v I__1149 (
            .O(N__5082),
            .I(N__5079));
    Odrv12 I__1148 (
            .O(N__5079),
            .I(SIZ_c_1));
    CascadeMux I__1147 (
            .O(N__5076),
            .I(N__5073));
    InMux I__1146 (
            .O(N__5073),
            .I(N__5067));
    InMux I__1145 (
            .O(N__5072),
            .I(N__5067));
    LocalMux I__1144 (
            .O(N__5067),
            .I(N__5064));
    Span12Mux_h I__1143 (
            .O(N__5064),
            .I(N__5061));
    Span12Mux_v I__1142 (
            .O(N__5061),
            .I(N__5058));
    Odrv12 I__1141 (
            .O(N__5058),
            .I(SIZ_c_0));
    InMux I__1140 (
            .O(N__5055),
            .I(N__5052));
    LocalMux I__1139 (
            .O(N__5052),
            .I(N__5049));
    Span4Mux_h I__1138 (
            .O(N__5049),
            .I(N__5044));
    InMux I__1137 (
            .O(N__5048),
            .I(N__5039));
    InMux I__1136 (
            .O(N__5047),
            .I(N__5039));
    Sp12to4 I__1135 (
            .O(N__5044),
            .I(N__5036));
    LocalMux I__1134 (
            .O(N__5039),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    Odrv12 I__1133 (
            .O(N__5036),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    CascadeMux I__1132 (
            .O(N__5031),
            .I(\U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ));
    InMux I__1131 (
            .O(N__5028),
            .I(N__5025));
    LocalMux I__1130 (
            .O(N__5025),
            .I(N__5022));
    Span4Mux_h I__1129 (
            .O(N__5022),
            .I(N__5019));
    Sp12to4 I__1128 (
            .O(N__5019),
            .I(N__5016));
    Span12Mux_v I__1127 (
            .O(N__5016),
            .I(N__5013));
    Odrv12 I__1126 (
            .O(N__5013),
            .I(TS_CPUn_c));
    InMux I__1125 (
            .O(N__5010),
            .I(N__5007));
    LocalMux I__1124 (
            .O(N__5007),
            .I(\U111_CYCLE_SM.TS_EN_5 ));
    InMux I__1123 (
            .O(N__5004),
            .I(N__5001));
    LocalMux I__1122 (
            .O(N__5001),
            .I(\U111_CYCLE_SM.N_69_0 ));
    IoInMux I__1121 (
            .O(N__4998),
            .I(N__4995));
    LocalMux I__1120 (
            .O(N__4995),
            .I(N__4991));
    IoInMux I__1119 (
            .O(N__4994),
            .I(N__4986));
    IoSpan4Mux I__1118 (
            .O(N__4991),
            .I(N__4983));
    IoInMux I__1117 (
            .O(N__4990),
            .I(N__4978));
    IoInMux I__1116 (
            .O(N__4989),
            .I(N__4978));
    LocalMux I__1115 (
            .O(N__4986),
            .I(N__4975));
    IoSpan4Mux I__1114 (
            .O(N__4983),
            .I(N__4972));
    LocalMux I__1113 (
            .O(N__4978),
            .I(N__4969));
    Span4Mux_s3_h I__1112 (
            .O(N__4975),
            .I(N__4966));
    IoSpan4Mux I__1111 (
            .O(N__4972),
            .I(N__4961));
    IoSpan4Mux I__1110 (
            .O(N__4969),
            .I(N__4961));
    Span4Mux_v I__1109 (
            .O(N__4966),
            .I(N__4958));
    Span4Mux_s2_v I__1108 (
            .O(N__4961),
            .I(N__4955));
    Sp12to4 I__1107 (
            .O(N__4958),
            .I(N__4952));
    Span4Mux_v I__1106 (
            .O(N__4955),
            .I(N__4949));
    Span12Mux_h I__1105 (
            .O(N__4952),
            .I(N__4946));
    Span4Mux_v I__1104 (
            .O(N__4949),
            .I(N__4943));
    Odrv12 I__1103 (
            .O(N__4946),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1102 (
            .O(N__4943),
            .I(CONSTANT_ONE_NET));
    InMux I__1101 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__1100 (
            .O(N__4935),
            .I(N__4932));
    Span4Mux_v I__1099 (
            .O(N__4932),
            .I(N__4929));
    Span4Mux_h I__1098 (
            .O(N__4929),
            .I(N__4926));
    Sp12to4 I__1097 (
            .O(N__4926),
            .I(N__4923));
    Odrv12 I__1096 (
            .O(N__4923),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__1095 (
            .O(N__4920),
            .I(N__4917));
    LocalMux I__1094 (
            .O(N__4917),
            .I(N__4914));
    IoSpan4Mux I__1093 (
            .O(N__4914),
            .I(N__4911));
    Span4Mux_s2_h I__1092 (
            .O(N__4911),
            .I(N__4908));
    Span4Mux_h I__1091 (
            .O(N__4908),
            .I(N__4905));
    Sp12to4 I__1090 (
            .O(N__4905),
            .I(N__4902));
    Odrv12 I__1089 (
            .O(N__4902),
            .I(un1_D_LM_AMIGA_7));
    CascadeMux I__1088 (
            .O(N__4899),
            .I(N__4896));
    InMux I__1087 (
            .O(N__4896),
            .I(N__4893));
    LocalMux I__1086 (
            .O(N__4893),
            .I(N__4890));
    Span4Mux_v I__1085 (
            .O(N__4890),
            .I(N__4887));
    Span4Mux_v I__1084 (
            .O(N__4887),
            .I(N__4884));
    Sp12to4 I__1083 (
            .O(N__4884),
            .I(N__4881));
    Span12Mux_h I__1082 (
            .O(N__4881),
            .I(N__4878));
    Odrv12 I__1081 (
            .O(N__4878),
            .I(D_UM_040_in_7));
    IoInMux I__1080 (
            .O(N__4875),
            .I(N__4872));
    LocalMux I__1079 (
            .O(N__4872),
            .I(N__4869));
    IoSpan4Mux I__1078 (
            .O(N__4869),
            .I(N__4865));
    InMux I__1077 (
            .O(N__4868),
            .I(N__4862));
    Span4Mux_s3_h I__1076 (
            .O(N__4865),
            .I(N__4859));
    LocalMux I__1075 (
            .O(N__4862),
            .I(N__4856));
    Sp12to4 I__1074 (
            .O(N__4859),
            .I(N__4853));
    Sp12to4 I__1073 (
            .O(N__4856),
            .I(N__4850));
    Span12Mux_v I__1072 (
            .O(N__4853),
            .I(N__4847));
    Span12Mux_v I__1071 (
            .O(N__4850),
            .I(N__4844));
    Span12Mux_h I__1070 (
            .O(N__4847),
            .I(N__4841));
    Span12Mux_h I__1069 (
            .O(N__4844),
            .I(N__4838));
    Span12Mux_h I__1068 (
            .O(N__4841),
            .I(N__4833));
    Span12Mux_v I__1067 (
            .O(N__4838),
            .I(N__4833));
    Odrv12 I__1066 (
            .O(N__4833),
            .I(D_LL_040_in_7));
    IoInMux I__1065 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__1064 (
            .O(N__4827),
            .I(N__4824));
    Span12Mux_s2_h I__1063 (
            .O(N__4824),
            .I(N__4821));
    Span12Mux_h I__1062 (
            .O(N__4821),
            .I(N__4818));
    Odrv12 I__1061 (
            .O(N__4818),
            .I(un1_D_UM_040_7));
    InMux I__1060 (
            .O(N__4815),
            .I(N__4812));
    LocalMux I__1059 (
            .O(N__4812),
            .I(N__4809));
    Sp12to4 I__1058 (
            .O(N__4809),
            .I(N__4806));
    Span12Mux_v I__1057 (
            .O(N__4806),
            .I(N__4803));
    Span12Mux_h I__1056 (
            .O(N__4803),
            .I(N__4800));
    Odrv12 I__1055 (
            .O(N__4800),
            .I(D_UU_040_in_0));
    IoInMux I__1054 (
            .O(N__4797),
            .I(N__4793));
    CascadeMux I__1053 (
            .O(N__4796),
            .I(N__4790));
    LocalMux I__1052 (
            .O(N__4793),
            .I(N__4787));
    InMux I__1051 (
            .O(N__4790),
            .I(N__4784));
    IoSpan4Mux I__1050 (
            .O(N__4787),
            .I(N__4781));
    LocalMux I__1049 (
            .O(N__4784),
            .I(N__4778));
    IoSpan4Mux I__1048 (
            .O(N__4781),
            .I(N__4775));
    Span4Mux_h I__1047 (
            .O(N__4778),
            .I(N__4772));
    Span4Mux_s2_h I__1046 (
            .O(N__4775),
            .I(N__4769));
    Sp12to4 I__1045 (
            .O(N__4772),
            .I(N__4766));
    Sp12to4 I__1044 (
            .O(N__4769),
            .I(N__4763));
    Span12Mux_v I__1043 (
            .O(N__4766),
            .I(N__4760));
    Span12Mux_h I__1042 (
            .O(N__4763),
            .I(N__4757));
    Span12Mux_v I__1041 (
            .O(N__4760),
            .I(N__4754));
    Span12Mux_h I__1040 (
            .O(N__4757),
            .I(N__4751));
    Span12Mux_h I__1039 (
            .O(N__4754),
            .I(N__4748));
    Odrv12 I__1038 (
            .O(N__4751),
            .I(D_LM_040_in_0));
    Odrv12 I__1037 (
            .O(N__4748),
            .I(D_LM_040_in_0));
    IoInMux I__1036 (
            .O(N__4743),
            .I(N__4740));
    LocalMux I__1035 (
            .O(N__4740),
            .I(N__4737));
    Span4Mux_s3_v I__1034 (
            .O(N__4737),
            .I(N__4734));
    Sp12to4 I__1033 (
            .O(N__4734),
            .I(N__4731));
    Span12Mux_h I__1032 (
            .O(N__4731),
            .I(N__4728));
    Odrv12 I__1031 (
            .O(N__4728),
            .I(un1_D_UU_040_0));
    IoInMux I__1030 (
            .O(N__4725),
            .I(N__4721));
    CascadeMux I__1029 (
            .O(N__4724),
            .I(N__4718));
    LocalMux I__1028 (
            .O(N__4721),
            .I(N__4715));
    InMux I__1027 (
            .O(N__4718),
            .I(N__4712));
    IoSpan4Mux I__1026 (
            .O(N__4715),
            .I(N__4709));
    LocalMux I__1025 (
            .O(N__4712),
            .I(N__4706));
    Span4Mux_s3_h I__1024 (
            .O(N__4709),
            .I(N__4703));
    Sp12to4 I__1023 (
            .O(N__4706),
            .I(N__4700));
    Sp12to4 I__1022 (
            .O(N__4703),
            .I(N__4697));
    Span12Mux_v I__1021 (
            .O(N__4700),
            .I(N__4694));
    Span12Mux_v I__1020 (
            .O(N__4697),
            .I(N__4691));
    Span12Mux_v I__1019 (
            .O(N__4694),
            .I(N__4686));
    Span12Mux_h I__1018 (
            .O(N__4691),
            .I(N__4686));
    Span12Mux_h I__1017 (
            .O(N__4686),
            .I(N__4683));
    Odrv12 I__1016 (
            .O(N__4683),
            .I(D_LL_040_in_5));
    InMux I__1015 (
            .O(N__4680),
            .I(N__4677));
    LocalMux I__1014 (
            .O(N__4677),
            .I(N__4674));
    Span4Mux_v I__1013 (
            .O(N__4674),
            .I(N__4671));
    Span4Mux_h I__1012 (
            .O(N__4671),
            .I(N__4668));
    Sp12to4 I__1011 (
            .O(N__4668),
            .I(N__4665));
    Span12Mux_h I__1010 (
            .O(N__4665),
            .I(N__4662));
    Odrv12 I__1009 (
            .O(N__4662),
            .I(D_UM_040_in_5));
    IoInMux I__1008 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__1007 (
            .O(N__4656),
            .I(N__4653));
    IoSpan4Mux I__1006 (
            .O(N__4653),
            .I(N__4650));
    IoSpan4Mux I__1005 (
            .O(N__4650),
            .I(N__4647));
    Span4Mux_s2_v I__1004 (
            .O(N__4647),
            .I(N__4644));
    Span4Mux_v I__1003 (
            .O(N__4644),
            .I(N__4641));
    Odrv4 I__1002 (
            .O(N__4641),
            .I(un1_D_UM_040_5));
    InMux I__1001 (
            .O(N__4638),
            .I(N__4635));
    LocalMux I__1000 (
            .O(N__4635),
            .I(N__4632));
    Span4Mux_v I__999 (
            .O(N__4632),
            .I(N__4629));
    Span4Mux_h I__998 (
            .O(N__4629),
            .I(N__4626));
    Sp12to4 I__997 (
            .O(N__4626),
            .I(N__4623));
    Span12Mux_h I__996 (
            .O(N__4623),
            .I(N__4620));
    Odrv12 I__995 (
            .O(N__4620),
            .I(D_UU_040_in_5));
    IoInMux I__994 (
            .O(N__4617),
            .I(N__4614));
    LocalMux I__993 (
            .O(N__4614),
            .I(N__4610));
    CascadeMux I__992 (
            .O(N__4613),
            .I(N__4607));
    IoSpan4Mux I__991 (
            .O(N__4610),
            .I(N__4604));
    InMux I__990 (
            .O(N__4607),
            .I(N__4601));
    Span4Mux_s2_h I__989 (
            .O(N__4604),
            .I(N__4598));
    LocalMux I__988 (
            .O(N__4601),
            .I(N__4595));
    Span4Mux_v I__987 (
            .O(N__4598),
            .I(N__4592));
    Span4Mux_v I__986 (
            .O(N__4595),
            .I(N__4589));
    Sp12to4 I__985 (
            .O(N__4592),
            .I(N__4586));
    Sp12to4 I__984 (
            .O(N__4589),
            .I(N__4583));
    Span12Mux_s9_h I__983 (
            .O(N__4586),
            .I(N__4580));
    Span12Mux_h I__982 (
            .O(N__4583),
            .I(N__4577));
    Span12Mux_h I__981 (
            .O(N__4580),
            .I(N__4574));
    Span12Mux_v I__980 (
            .O(N__4577),
            .I(N__4571));
    Odrv12 I__979 (
            .O(N__4574),
            .I(D_LM_040_in_5));
    Odrv12 I__978 (
            .O(N__4571),
            .I(D_LM_040_in_5));
    CascadeMux I__977 (
            .O(N__4566),
            .I(N__4555));
    InMux I__976 (
            .O(N__4565),
            .I(N__4549));
    InMux I__975 (
            .O(N__4564),
            .I(N__4549));
    CascadeMux I__974 (
            .O(N__4563),
            .I(N__4546));
    InMux I__973 (
            .O(N__4562),
            .I(N__4543));
    InMux I__972 (
            .O(N__4561),
            .I(N__4540));
    CascadeMux I__971 (
            .O(N__4560),
            .I(N__4536));
    InMux I__970 (
            .O(N__4559),
            .I(N__4533));
    InMux I__969 (
            .O(N__4558),
            .I(N__4530));
    InMux I__968 (
            .O(N__4555),
            .I(N__4527));
    CascadeMux I__967 (
            .O(N__4554),
            .I(N__4522));
    LocalMux I__966 (
            .O(N__4549),
            .I(N__4519));
    InMux I__965 (
            .O(N__4546),
            .I(N__4516));
    LocalMux I__964 (
            .O(N__4543),
            .I(N__4511));
    LocalMux I__963 (
            .O(N__4540),
            .I(N__4511));
    InMux I__962 (
            .O(N__4539),
            .I(N__4508));
    InMux I__961 (
            .O(N__4536),
            .I(N__4505));
    LocalMux I__960 (
            .O(N__4533),
            .I(N__4496));
    LocalMux I__959 (
            .O(N__4530),
            .I(N__4496));
    LocalMux I__958 (
            .O(N__4527),
            .I(N__4496));
    InMux I__957 (
            .O(N__4526),
            .I(N__4493));
    InMux I__956 (
            .O(N__4525),
            .I(N__4487));
    InMux I__955 (
            .O(N__4522),
            .I(N__4487));
    Span4Mux_v I__954 (
            .O(N__4519),
            .I(N__4482));
    LocalMux I__953 (
            .O(N__4516),
            .I(N__4482));
    Span4Mux_v I__952 (
            .O(N__4511),
            .I(N__4473));
    LocalMux I__951 (
            .O(N__4508),
            .I(N__4473));
    LocalMux I__950 (
            .O(N__4505),
            .I(N__4473));
    InMux I__949 (
            .O(N__4504),
            .I(N__4470));
    InMux I__948 (
            .O(N__4503),
            .I(N__4467));
    Span4Mux_v I__947 (
            .O(N__4496),
            .I(N__4461));
    LocalMux I__946 (
            .O(N__4493),
            .I(N__4461));
    InMux I__945 (
            .O(N__4492),
            .I(N__4458));
    LocalMux I__944 (
            .O(N__4487),
            .I(N__4454));
    Span4Mux_v I__943 (
            .O(N__4482),
            .I(N__4445));
    InMux I__942 (
            .O(N__4481),
            .I(N__4440));
    InMux I__941 (
            .O(N__4480),
            .I(N__4440));
    Span4Mux_v I__940 (
            .O(N__4473),
            .I(N__4431));
    LocalMux I__939 (
            .O(N__4470),
            .I(N__4431));
    LocalMux I__938 (
            .O(N__4467),
            .I(N__4431));
    InMux I__937 (
            .O(N__4466),
            .I(N__4428));
    Span4Mux_v I__936 (
            .O(N__4461),
            .I(N__4422));
    LocalMux I__935 (
            .O(N__4458),
            .I(N__4422));
    InMux I__934 (
            .O(N__4457),
            .I(N__4419));
    Span4Mux_v I__933 (
            .O(N__4454),
            .I(N__4416));
    InMux I__932 (
            .O(N__4453),
            .I(N__4413));
    InMux I__931 (
            .O(N__4452),
            .I(N__4410));
    InMux I__930 (
            .O(N__4451),
            .I(N__4404));
    InMux I__929 (
            .O(N__4450),
            .I(N__4404));
    InMux I__928 (
            .O(N__4449),
            .I(N__4401));
    InMux I__927 (
            .O(N__4448),
            .I(N__4397));
    Span4Mux_v I__926 (
            .O(N__4445),
            .I(N__4392));
    LocalMux I__925 (
            .O(N__4440),
            .I(N__4392));
    InMux I__924 (
            .O(N__4439),
            .I(N__4387));
    InMux I__923 (
            .O(N__4438),
            .I(N__4387));
    Span4Mux_v I__922 (
            .O(N__4431),
            .I(N__4382));
    LocalMux I__921 (
            .O(N__4428),
            .I(N__4382));
    InMux I__920 (
            .O(N__4427),
            .I(N__4379));
    Span4Mux_v I__919 (
            .O(N__4422),
            .I(N__4374));
    LocalMux I__918 (
            .O(N__4419),
            .I(N__4374));
    Span4Mux_v I__917 (
            .O(N__4416),
            .I(N__4367));
    LocalMux I__916 (
            .O(N__4413),
            .I(N__4367));
    LocalMux I__915 (
            .O(N__4410),
            .I(N__4367));
    InMux I__914 (
            .O(N__4409),
            .I(N__4364));
    LocalMux I__913 (
            .O(N__4404),
            .I(N__4358));
    LocalMux I__912 (
            .O(N__4401),
            .I(N__4358));
    IoInMux I__911 (
            .O(N__4400),
            .I(N__4355));
    LocalMux I__910 (
            .O(N__4397),
            .I(N__4352));
    Span4Mux_v I__909 (
            .O(N__4392),
            .I(N__4347));
    LocalMux I__908 (
            .O(N__4387),
            .I(N__4347));
    Span4Mux_v I__907 (
            .O(N__4382),
            .I(N__4342));
    LocalMux I__906 (
            .O(N__4379),
            .I(N__4342));
    Span4Mux_v I__905 (
            .O(N__4374),
            .I(N__4338));
    Span4Mux_v I__904 (
            .O(N__4367),
            .I(N__4333));
    LocalMux I__903 (
            .O(N__4364),
            .I(N__4333));
    InMux I__902 (
            .O(N__4363),
            .I(N__4330));
    Span12Mux_h I__901 (
            .O(N__4358),
            .I(N__4327));
    LocalMux I__900 (
            .O(N__4355),
            .I(N__4324));
    Span12Mux_h I__899 (
            .O(N__4352),
            .I(N__4321));
    Span4Mux_v I__898 (
            .O(N__4347),
            .I(N__4318));
    Span4Mux_v I__897 (
            .O(N__4342),
            .I(N__4315));
    InMux I__896 (
            .O(N__4341),
            .I(N__4312));
    Span4Mux_h I__895 (
            .O(N__4338),
            .I(N__4305));
    Span4Mux_v I__894 (
            .O(N__4333),
            .I(N__4305));
    LocalMux I__893 (
            .O(N__4330),
            .I(N__4305));
    Span12Mux_v I__892 (
            .O(N__4327),
            .I(N__4302));
    Span4Mux_s3_v I__891 (
            .O(N__4324),
            .I(N__4299));
    Span12Mux_v I__890 (
            .O(N__4321),
            .I(N__4290));
    Sp12to4 I__889 (
            .O(N__4318),
            .I(N__4290));
    Sp12to4 I__888 (
            .O(N__4315),
            .I(N__4290));
    LocalMux I__887 (
            .O(N__4312),
            .I(N__4290));
    Span4Mux_v I__886 (
            .O(N__4305),
            .I(N__4287));
    Odrv12 I__885 (
            .O(N__4302),
            .I(A_AMIGA_c_1));
    Odrv4 I__884 (
            .O(N__4299),
            .I(A_AMIGA_c_1));
    Odrv12 I__883 (
            .O(N__4290),
            .I(A_AMIGA_c_1));
    Odrv4 I__882 (
            .O(N__4287),
            .I(A_AMIGA_c_1));
    IoInMux I__881 (
            .O(N__4278),
            .I(N__4275));
    LocalMux I__880 (
            .O(N__4275),
            .I(N__4272));
    Span12Mux_s2_h I__879 (
            .O(N__4272),
            .I(N__4269));
    Span12Mux_h I__878 (
            .O(N__4269),
            .I(N__4266));
    Odrv12 I__877 (
            .O(N__4266),
            .I(un1_D_UU_040_5));
    InMux I__876 (
            .O(N__4263),
            .I(N__4260));
    LocalMux I__875 (
            .O(N__4260),
            .I(N__4257));
    Span4Mux_v I__874 (
            .O(N__4257),
            .I(N__4254));
    Odrv4 I__873 (
            .O(N__4254),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    CascadeMux I__872 (
            .O(N__4251),
            .I(N__4248));
    InMux I__871 (
            .O(N__4248),
            .I(N__4244));
    InMux I__870 (
            .O(N__4247),
            .I(N__4241));
    LocalMux I__869 (
            .O(N__4244),
            .I(N__4237));
    LocalMux I__868 (
            .O(N__4241),
            .I(N__4234));
    InMux I__867 (
            .O(N__4240),
            .I(N__4231));
    Span4Mux_v I__866 (
            .O(N__4237),
            .I(N__4228));
    Span4Mux_v I__865 (
            .O(N__4234),
            .I(N__4223));
    LocalMux I__864 (
            .O(N__4231),
            .I(N__4223));
    Span4Mux_v I__863 (
            .O(N__4228),
            .I(N__4220));
    Span4Mux_v I__862 (
            .O(N__4223),
            .I(N__4217));
    Sp12to4 I__861 (
            .O(N__4220),
            .I(N__4212));
    Sp12to4 I__860 (
            .O(N__4217),
            .I(N__4212));
    Span12Mux_h I__859 (
            .O(N__4212),
            .I(N__4209));
    Odrv12 I__858 (
            .O(N__4209),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__857 (
            .O(N__4206),
            .I(N__4203));
    LocalMux I__856 (
            .O(N__4203),
            .I(N__4200));
    IoSpan4Mux I__855 (
            .O(N__4200),
            .I(N__4197));
    Sp12to4 I__854 (
            .O(N__4197),
            .I(N__4194));
    Span12Mux_s6_v I__853 (
            .O(N__4194),
            .I(N__4191));
    Odrv12 I__852 (
            .O(N__4191),
            .I(un1_D_UU_AMIGA_6));
    InMux I__851 (
            .O(N__4188),
            .I(N__4185));
    LocalMux I__850 (
            .O(N__4185),
            .I(N__4182));
    Span12Mux_h I__849 (
            .O(N__4182),
            .I(N__4179));
    Odrv12 I__848 (
            .O(N__4179),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__847 (
            .O(N__4176),
            .I(N__4173));
    LocalMux I__846 (
            .O(N__4173),
            .I(N__4170));
    IoSpan4Mux I__845 (
            .O(N__4170),
            .I(N__4167));
    IoSpan4Mux I__844 (
            .O(N__4167),
            .I(N__4164));
    Sp12to4 I__843 (
            .O(N__4164),
            .I(N__4161));
    Span12Mux_s7_h I__842 (
            .O(N__4161),
            .I(N__4158));
    Odrv12 I__841 (
            .O(N__4158),
            .I(un1_D_LM_AMIGA_0));
    IoInMux I__840 (
            .O(N__4155),
            .I(N__4152));
    LocalMux I__839 (
            .O(N__4152),
            .I(N__4149));
    Span12Mux_s9_h I__838 (
            .O(N__4149),
            .I(N__4146));
    Odrv12 I__837 (
            .O(N__4146),
            .I(un1_D_UM_AMIGA_0));
    SRMux I__836 (
            .O(N__4143),
            .I(N__4140));
    LocalMux I__835 (
            .O(N__4140),
            .I(N__4137));
    Odrv4 I__834 (
            .O(N__4137),
            .I(\U111_CYCLE_SM.RESETn_c_i ));
    InMux I__833 (
            .O(N__4134),
            .I(N__4131));
    LocalMux I__832 (
            .O(N__4131),
            .I(N__4128));
    Span4Mux_h I__831 (
            .O(N__4128),
            .I(N__4125));
    Sp12to4 I__830 (
            .O(N__4125),
            .I(N__4122));
    Span12Mux_v I__829 (
            .O(N__4122),
            .I(N__4118));
    InMux I__828 (
            .O(N__4121),
            .I(N__4115));
    Odrv12 I__827 (
            .O(N__4118),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    LocalMux I__826 (
            .O(N__4115),
            .I(\U111_CYCLE_SM.A_OUTZ0 ));
    InMux I__825 (
            .O(N__4110),
            .I(N__4107));
    LocalMux I__824 (
            .O(N__4107),
            .I(\U111_CYCLE_SM.A_OUT_0 ));
    CascadeMux I__823 (
            .O(N__4104),
            .I(N__4101));
    InMux I__822 (
            .O(N__4101),
            .I(N__4098));
    LocalMux I__821 (
            .O(N__4098),
            .I(N__4095));
    Span4Mux_v I__820 (
            .O(N__4095),
            .I(N__4091));
    InMux I__819 (
            .O(N__4094),
            .I(N__4088));
    Span4Mux_v I__818 (
            .O(N__4091),
            .I(N__4085));
    LocalMux I__817 (
            .O(N__4088),
            .I(N__4082));
    Span4Mux_v I__816 (
            .O(N__4085),
            .I(N__4078));
    Span4Mux_v I__815 (
            .O(N__4082),
            .I(N__4075));
    InMux I__814 (
            .O(N__4081),
            .I(N__4072));
    Sp12to4 I__813 (
            .O(N__4078),
            .I(N__4065));
    Sp12to4 I__812 (
            .O(N__4075),
            .I(N__4065));
    LocalMux I__811 (
            .O(N__4072),
            .I(N__4065));
    Span12Mux_h I__810 (
            .O(N__4065),
            .I(N__4062));
    Odrv12 I__809 (
            .O(N__4062),
            .I(D_UM_AMIGA_in_0));
    InMux I__808 (
            .O(N__4059),
            .I(N__4056));
    LocalMux I__807 (
            .O(N__4056),
            .I(N__4053));
    Odrv12 I__806 (
            .O(N__4053),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__805 (
            .O(N__4050),
            .I(N__4047));
    LocalMux I__804 (
            .O(N__4047),
            .I(N__4044));
    Span4Mux_v I__803 (
            .O(N__4044),
            .I(N__4041));
    Sp12to4 I__802 (
            .O(N__4041),
            .I(N__4038));
    Span12Mux_h I__801 (
            .O(N__4038),
            .I(N__4035));
    Odrv12 I__800 (
            .O(N__4035),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__799 (
            .O(N__4032),
            .I(N__4029));
    LocalMux I__798 (
            .O(N__4029),
            .I(N__4026));
    IoSpan4Mux I__797 (
            .O(N__4026),
            .I(N__4023));
    IoSpan4Mux I__796 (
            .O(N__4023),
            .I(N__4020));
    Span4Mux_s2_h I__795 (
            .O(N__4020),
            .I(N__4017));
    Sp12to4 I__794 (
            .O(N__4017),
            .I(N__4014));
    Span12Mux_s10_h I__793 (
            .O(N__4014),
            .I(N__4011));
    Odrv12 I__792 (
            .O(N__4011),
            .I(un1_D_LM_AMIGA_4));
    InMux I__791 (
            .O(N__4008),
            .I(N__4005));
    LocalMux I__790 (
            .O(N__4005),
            .I(N__4002));
    Span4Mux_v I__789 (
            .O(N__4002),
            .I(N__3999));
    Span4Mux_v I__788 (
            .O(N__3999),
            .I(N__3996));
    Sp12to4 I__787 (
            .O(N__3996),
            .I(N__3993));
    Span12Mux_h I__786 (
            .O(N__3993),
            .I(N__3990));
    Odrv12 I__785 (
            .O(N__3990),
            .I(D_UU_040_in_1));
    IoInMux I__784 (
            .O(N__3987),
            .I(N__3983));
    InMux I__783 (
            .O(N__3986),
            .I(N__3980));
    LocalMux I__782 (
            .O(N__3983),
            .I(N__3977));
    LocalMux I__781 (
            .O(N__3980),
            .I(N__3974));
    Span4Mux_s3_h I__780 (
            .O(N__3977),
            .I(N__3971));
    Span4Mux_h I__779 (
            .O(N__3974),
            .I(N__3968));
    Sp12to4 I__778 (
            .O(N__3971),
            .I(N__3965));
    Sp12to4 I__777 (
            .O(N__3968),
            .I(N__3962));
    Span12Mux_v I__776 (
            .O(N__3965),
            .I(N__3959));
    Span12Mux_v I__775 (
            .O(N__3962),
            .I(N__3956));
    Span12Mux_h I__774 (
            .O(N__3959),
            .I(N__3951));
    Span12Mux_v I__773 (
            .O(N__3956),
            .I(N__3951));
    Span12Mux_h I__772 (
            .O(N__3951),
            .I(N__3948));
    Odrv12 I__771 (
            .O(N__3948),
            .I(D_LM_040_in_1));
    IoInMux I__770 (
            .O(N__3945),
            .I(N__3942));
    LocalMux I__769 (
            .O(N__3942),
            .I(N__3939));
    IoSpan4Mux I__768 (
            .O(N__3939),
            .I(N__3936));
    Sp12to4 I__767 (
            .O(N__3936),
            .I(N__3933));
    Span12Mux_s6_h I__766 (
            .O(N__3933),
            .I(N__3930));
    Odrv12 I__765 (
            .O(N__3930),
            .I(un1_D_UU_040_1));
    CascadeMux I__764 (
            .O(N__3927),
            .I(N__3924));
    InMux I__763 (
            .O(N__3924),
            .I(N__3921));
    LocalMux I__762 (
            .O(N__3921),
            .I(N__3918));
    Span4Mux_v I__761 (
            .O(N__3918),
            .I(N__3915));
    Sp12to4 I__760 (
            .O(N__3915),
            .I(N__3912));
    Span12Mux_h I__759 (
            .O(N__3912),
            .I(N__3909));
    Odrv12 I__758 (
            .O(N__3909),
            .I(D_UU_040_in_2));
    InMux I__757 (
            .O(N__3906),
            .I(N__3902));
    IoInMux I__756 (
            .O(N__3905),
            .I(N__3899));
    LocalMux I__755 (
            .O(N__3902),
            .I(N__3896));
    LocalMux I__754 (
            .O(N__3899),
            .I(N__3893));
    Sp12to4 I__753 (
            .O(N__3896),
            .I(N__3890));
    Span12Mux_s9_h I__752 (
            .O(N__3893),
            .I(N__3887));
    Span12Mux_v I__751 (
            .O(N__3890),
            .I(N__3884));
    Span12Mux_v I__750 (
            .O(N__3887),
            .I(N__3881));
    Span12Mux_v I__749 (
            .O(N__3884),
            .I(N__3878));
    Span12Mux_h I__748 (
            .O(N__3881),
            .I(N__3875));
    Span12Mux_h I__747 (
            .O(N__3878),
            .I(N__3872));
    Odrv12 I__746 (
            .O(N__3875),
            .I(D_LM_040_in_2));
    Odrv12 I__745 (
            .O(N__3872),
            .I(D_LM_040_in_2));
    IoInMux I__744 (
            .O(N__3867),
            .I(N__3864));
    LocalMux I__743 (
            .O(N__3864),
            .I(N__3861));
    IoSpan4Mux I__742 (
            .O(N__3861),
            .I(N__3858));
    IoSpan4Mux I__741 (
            .O(N__3858),
            .I(N__3855));
    Span4Mux_s2_v I__740 (
            .O(N__3855),
            .I(N__3852));
    Span4Mux_v I__739 (
            .O(N__3852),
            .I(N__3849));
    Odrv4 I__738 (
            .O(N__3849),
            .I(un1_D_UU_040_2));
    CascadeMux I__737 (
            .O(N__3846),
            .I(N__3843));
    InMux I__736 (
            .O(N__3843),
            .I(N__3840));
    LocalMux I__735 (
            .O(N__3840),
            .I(N__3837));
    Span4Mux_v I__734 (
            .O(N__3837),
            .I(N__3834));
    Span4Mux_h I__733 (
            .O(N__3834),
            .I(N__3831));
    Sp12to4 I__732 (
            .O(N__3831),
            .I(N__3828));
    Odrv12 I__731 (
            .O(N__3828),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__730 (
            .O(N__3825),
            .I(N__3822));
    LocalMux I__729 (
            .O(N__3822),
            .I(N__3819));
    Span4Mux_s3_h I__728 (
            .O(N__3819),
            .I(N__3816));
    Span4Mux_v I__727 (
            .O(N__3816),
            .I(N__3813));
    Span4Mux_v I__726 (
            .O(N__3813),
            .I(N__3810));
    Span4Mux_h I__725 (
            .O(N__3810),
            .I(N__3807));
    Sp12to4 I__724 (
            .O(N__3807),
            .I(N__3804));
    Odrv12 I__723 (
            .O(N__3804),
            .I(un1_D_LL_AMIGA_6));
    InMux I__722 (
            .O(N__3801),
            .I(N__3797));
    IoInMux I__721 (
            .O(N__3800),
            .I(N__3794));
    LocalMux I__720 (
            .O(N__3797),
            .I(N__3791));
    LocalMux I__719 (
            .O(N__3794),
            .I(N__3788));
    Span4Mux_v I__718 (
            .O(N__3791),
            .I(N__3785));
    Span4Mux_s3_h I__717 (
            .O(N__3788),
            .I(N__3782));
    Sp12to4 I__716 (
            .O(N__3785),
            .I(N__3779));
    Sp12to4 I__715 (
            .O(N__3782),
            .I(N__3776));
    Span12Mux_h I__714 (
            .O(N__3779),
            .I(N__3773));
    Span12Mux_v I__713 (
            .O(N__3776),
            .I(N__3770));
    Span12Mux_v I__712 (
            .O(N__3773),
            .I(N__3767));
    Span12Mux_h I__711 (
            .O(N__3770),
            .I(N__3764));
    Span12Mux_v I__710 (
            .O(N__3767),
            .I(N__3759));
    Span12Mux_h I__709 (
            .O(N__3764),
            .I(N__3759));
    Odrv12 I__708 (
            .O(N__3759),
            .I(D_LL_040_in_3));
    CascadeMux I__707 (
            .O(N__3756),
            .I(N__3753));
    InMux I__706 (
            .O(N__3753),
            .I(N__3750));
    LocalMux I__705 (
            .O(N__3750),
            .I(N__3747));
    Span4Mux_h I__704 (
            .O(N__3747),
            .I(N__3744));
    Sp12to4 I__703 (
            .O(N__3744),
            .I(N__3741));
    Span12Mux_v I__702 (
            .O(N__3741),
            .I(N__3738));
    Span12Mux_h I__701 (
            .O(N__3738),
            .I(N__3735));
    Odrv12 I__700 (
            .O(N__3735),
            .I(D_UM_040_in_3));
    IoInMux I__699 (
            .O(N__3732),
            .I(N__3729));
    LocalMux I__698 (
            .O(N__3729),
            .I(N__3726));
    IoSpan4Mux I__697 (
            .O(N__3726),
            .I(N__3723));
    Span4Mux_s3_h I__696 (
            .O(N__3723),
            .I(N__3720));
    Span4Mux_h I__695 (
            .O(N__3720),
            .I(N__3717));
    Span4Mux_h I__694 (
            .O(N__3717),
            .I(N__3714));
    Odrv4 I__693 (
            .O(N__3714),
            .I(un1_D_UM_040_3));
    InMux I__692 (
            .O(N__3711),
            .I(N__3708));
    LocalMux I__691 (
            .O(N__3708),
            .I(N__3705));
    Span4Mux_v I__690 (
            .O(N__3705),
            .I(N__3702));
    Span4Mux_h I__689 (
            .O(N__3702),
            .I(N__3699));
    Sp12to4 I__688 (
            .O(N__3699),
            .I(N__3696));
    Odrv12 I__687 (
            .O(N__3696),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__686 (
            .O(N__3693),
            .I(N__3690));
    LocalMux I__685 (
            .O(N__3690),
            .I(N__3687));
    IoSpan4Mux I__684 (
            .O(N__3687),
            .I(N__3684));
    Sp12to4 I__683 (
            .O(N__3684),
            .I(N__3681));
    Span12Mux_s7_v I__682 (
            .O(N__3681),
            .I(N__3678));
    Span12Mux_h I__681 (
            .O(N__3678),
            .I(N__3675));
    Odrv12 I__680 (
            .O(N__3675),
            .I(un1_D_LL_AMIGA_3));
    InMux I__679 (
            .O(N__3672),
            .I(N__3669));
    LocalMux I__678 (
            .O(N__3669),
            .I(N__3666));
    Span4Mux_v I__677 (
            .O(N__3666),
            .I(N__3663));
    Sp12to4 I__676 (
            .O(N__3663),
            .I(N__3660));
    Span12Mux_h I__675 (
            .O(N__3660),
            .I(N__3657));
    Odrv12 I__674 (
            .O(N__3657),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__673 (
            .O(N__3654),
            .I(N__3651));
    LocalMux I__672 (
            .O(N__3651),
            .I(N__3648));
    IoSpan4Mux I__671 (
            .O(N__3648),
            .I(N__3645));
    Span4Mux_s3_h I__670 (
            .O(N__3645),
            .I(N__3642));
    Sp12to4 I__669 (
            .O(N__3642),
            .I(N__3639));
    Span12Mux_h I__668 (
            .O(N__3639),
            .I(N__3636));
    Odrv12 I__667 (
            .O(N__3636),
            .I(un1_D_LL_AMIGA_1));
    CascadeMux I__666 (
            .O(N__3633),
            .I(N__3630));
    InMux I__665 (
            .O(N__3630),
            .I(N__3627));
    LocalMux I__664 (
            .O(N__3627),
            .I(N__3624));
    Span4Mux_v I__663 (
            .O(N__3624),
            .I(N__3621));
    Sp12to4 I__662 (
            .O(N__3621),
            .I(N__3618));
    Span12Mux_h I__661 (
            .O(N__3618),
            .I(N__3615));
    Odrv12 I__660 (
            .O(N__3615),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__659 (
            .O(N__3612),
            .I(N__3609));
    LocalMux I__658 (
            .O(N__3609),
            .I(N__3606));
    Span4Mux_s1_h I__657 (
            .O(N__3606),
            .I(N__3603));
    Span4Mux_h I__656 (
            .O(N__3603),
            .I(N__3600));
    Sp12to4 I__655 (
            .O(N__3600),
            .I(N__3597));
    Span12Mux_s9_v I__654 (
            .O(N__3597),
            .I(N__3594));
    Span12Mux_h I__653 (
            .O(N__3594),
            .I(N__3591));
    Odrv12 I__652 (
            .O(N__3591),
            .I(un1_D_LL_AMIGA_5));
    CascadeMux I__651 (
            .O(N__3588),
            .I(N__3585));
    InMux I__650 (
            .O(N__3585),
            .I(N__3582));
    LocalMux I__649 (
            .O(N__3582),
            .I(N__3579));
    Span12Mux_v I__648 (
            .O(N__3579),
            .I(N__3576));
    Odrv12 I__647 (
            .O(N__3576),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__646 (
            .O(N__3573),
            .I(N__3570));
    LocalMux I__645 (
            .O(N__3570),
            .I(N__3567));
    IoSpan4Mux I__644 (
            .O(N__3567),
            .I(N__3564));
    Span4Mux_s0_h I__643 (
            .O(N__3564),
            .I(N__3561));
    Sp12to4 I__642 (
            .O(N__3561),
            .I(N__3558));
    Span12Mux_s8_v I__641 (
            .O(N__3558),
            .I(N__3555));
    Span12Mux_h I__640 (
            .O(N__3555),
            .I(N__3552));
    Odrv12 I__639 (
            .O(N__3552),
            .I(un1_D_LL_AMIGA_4));
    CascadeMux I__638 (
            .O(N__3549),
            .I(N__3546));
    InMux I__637 (
            .O(N__3546),
            .I(N__3543));
    LocalMux I__636 (
            .O(N__3543),
            .I(N__3540));
    Span12Mux_h I__635 (
            .O(N__3540),
            .I(N__3537));
    Odrv12 I__634 (
            .O(N__3537),
            .I(D_UM_040_in_2));
    IoInMux I__633 (
            .O(N__3534),
            .I(N__3531));
    LocalMux I__632 (
            .O(N__3531),
            .I(N__3527));
    InMux I__631 (
            .O(N__3530),
            .I(N__3524));
    IoSpan4Mux I__630 (
            .O(N__3527),
            .I(N__3521));
    LocalMux I__629 (
            .O(N__3524),
            .I(N__3518));
    Span4Mux_s2_h I__628 (
            .O(N__3521),
            .I(N__3515));
    Span4Mux_v I__627 (
            .O(N__3518),
            .I(N__3512));
    Sp12to4 I__626 (
            .O(N__3515),
            .I(N__3509));
    Sp12to4 I__625 (
            .O(N__3512),
            .I(N__3506));
    Span12Mux_h I__624 (
            .O(N__3509),
            .I(N__3503));
    Span12Mux_h I__623 (
            .O(N__3506),
            .I(N__3500));
    Span12Mux_h I__622 (
            .O(N__3503),
            .I(N__3495));
    Span12Mux_v I__621 (
            .O(N__3500),
            .I(N__3495));
    Odrv12 I__620 (
            .O(N__3495),
            .I(D_LL_040_in_2));
    IoInMux I__619 (
            .O(N__3492),
            .I(N__3489));
    LocalMux I__618 (
            .O(N__3489),
            .I(N__3486));
    Span4Mux_s2_h I__617 (
            .O(N__3486),
            .I(N__3483));
    Span4Mux_h I__616 (
            .O(N__3483),
            .I(N__3480));
    Span4Mux_h I__615 (
            .O(N__3480),
            .I(N__3477));
    Span4Mux_v I__614 (
            .O(N__3477),
            .I(N__3474));
    Odrv4 I__613 (
            .O(N__3474),
            .I(un1_D_UM_040_2));
    InMux I__612 (
            .O(N__3471),
            .I(N__3468));
    LocalMux I__611 (
            .O(N__3468),
            .I(N__3465));
    Span12Mux_h I__610 (
            .O(N__3465),
            .I(N__3462));
    Odrv12 I__609 (
            .O(N__3462),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__608 (
            .O(N__3459),
            .I(N__3456));
    LocalMux I__607 (
            .O(N__3456),
            .I(N__3453));
    Span4Mux_s1_h I__606 (
            .O(N__3453),
            .I(N__3450));
    Sp12to4 I__605 (
            .O(N__3450),
            .I(N__3447));
    Span12Mux_v I__604 (
            .O(N__3447),
            .I(N__3444));
    Span12Mux_h I__603 (
            .O(N__3444),
            .I(N__3441));
    Odrv12 I__602 (
            .O(N__3441),
            .I(un1_D_LM_AMIGA_3));
    InMux I__601 (
            .O(N__3438),
            .I(N__3435));
    LocalMux I__600 (
            .O(N__3435),
            .I(N__3432));
    Span12Mux_v I__599 (
            .O(N__3432),
            .I(N__3429));
    Odrv12 I__598 (
            .O(N__3429),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__597 (
            .O(N__3426),
            .I(N__3423));
    LocalMux I__596 (
            .O(N__3423),
            .I(N__3420));
    Span4Mux_s2_h I__595 (
            .O(N__3420),
            .I(N__3417));
    Sp12to4 I__594 (
            .O(N__3417),
            .I(N__3414));
    Span12Mux_v I__593 (
            .O(N__3414),
            .I(N__3411));
    Span12Mux_h I__592 (
            .O(N__3411),
            .I(N__3408));
    Odrv12 I__591 (
            .O(N__3408),
            .I(un1_D_LM_AMIGA_5));
    CascadeMux I__590 (
            .O(N__3405),
            .I(N__3402));
    InMux I__589 (
            .O(N__3402),
            .I(N__3399));
    LocalMux I__588 (
            .O(N__3399),
            .I(N__3396));
    Span4Mux_v I__587 (
            .O(N__3396),
            .I(N__3393));
    Span4Mux_v I__586 (
            .O(N__3393),
            .I(N__3390));
    Sp12to4 I__585 (
            .O(N__3390),
            .I(N__3387));
    Span12Mux_h I__584 (
            .O(N__3387),
            .I(N__3384));
    Odrv12 I__583 (
            .O(N__3384),
            .I(D_UU_040_in_4));
    IoInMux I__582 (
            .O(N__3381),
            .I(N__3378));
    LocalMux I__581 (
            .O(N__3378),
            .I(N__3375));
    Span4Mux_s1_h I__580 (
            .O(N__3375),
            .I(N__3372));
    Sp12to4 I__579 (
            .O(N__3372),
            .I(N__3368));
    InMux I__578 (
            .O(N__3371),
            .I(N__3365));
    Span12Mux_v I__577 (
            .O(N__3368),
            .I(N__3362));
    LocalMux I__576 (
            .O(N__3365),
            .I(N__3359));
    Span12Mux_h I__575 (
            .O(N__3362),
            .I(N__3356));
    Span12Mux_h I__574 (
            .O(N__3359),
            .I(N__3353));
    Span12Mux_h I__573 (
            .O(N__3356),
            .I(N__3350));
    Span12Mux_v I__572 (
            .O(N__3353),
            .I(N__3347));
    Odrv12 I__571 (
            .O(N__3350),
            .I(D_LM_040_in_4));
    Odrv12 I__570 (
            .O(N__3347),
            .I(D_LM_040_in_4));
    IoInMux I__569 (
            .O(N__3342),
            .I(N__3339));
    LocalMux I__568 (
            .O(N__3339),
            .I(N__3336));
    Span12Mux_s6_v I__567 (
            .O(N__3336),
            .I(N__3333));
    Odrv12 I__566 (
            .O(N__3333),
            .I(un1_D_UU_040_4));
    InMux I__565 (
            .O(N__3330),
            .I(N__3327));
    LocalMux I__564 (
            .O(N__3327),
            .I(N__3324));
    Span4Mux_v I__563 (
            .O(N__3324),
            .I(N__3321));
    Span4Mux_h I__562 (
            .O(N__3321),
            .I(N__3318));
    Sp12to4 I__561 (
            .O(N__3318),
            .I(N__3315));
    Odrv12 I__560 (
            .O(N__3315),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__559 (
            .O(N__3312),
            .I(N__3309));
    LocalMux I__558 (
            .O(N__3309),
            .I(N__3306));
    IoSpan4Mux I__557 (
            .O(N__3306),
            .I(N__3303));
    Sp12to4 I__556 (
            .O(N__3303),
            .I(N__3300));
    Span12Mux_s7_h I__555 (
            .O(N__3300),
            .I(N__3297));
    Span12Mux_h I__554 (
            .O(N__3297),
            .I(N__3294));
    Odrv12 I__553 (
            .O(N__3294),
            .I(un1_D_LL_AMIGA_0));
    IoInMux I__552 (
            .O(N__3291),
            .I(N__3288));
    LocalMux I__551 (
            .O(N__3288),
            .I(N__3285));
    IoSpan4Mux I__550 (
            .O(N__3285),
            .I(N__3282));
    Span4Mux_s2_v I__549 (
            .O(N__3282),
            .I(N__3279));
    Odrv4 I__548 (
            .O(N__3279),
            .I(TSn_c));
    InMux I__547 (
            .O(N__3276),
            .I(N__3273));
    LocalMux I__546 (
            .O(N__3273),
            .I(N__3270));
    Span12Mux_h I__545 (
            .O(N__3270),
            .I(N__3267));
    Odrv12 I__544 (
            .O(N__3267),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__543 (
            .O(N__3264),
            .I(N__3261));
    LocalMux I__542 (
            .O(N__3261),
            .I(N__3258));
    Span12Mux_s2_h I__541 (
            .O(N__3258),
            .I(N__3255));
    Span12Mux_h I__540 (
            .O(N__3255),
            .I(N__3252));
    Span12Mux_v I__539 (
            .O(N__3252),
            .I(N__3249));
    Odrv12 I__538 (
            .O(N__3249),
            .I(un1_D_LM_AMIGA_2));
    InMux I__537 (
            .O(N__3246),
            .I(N__3243));
    LocalMux I__536 (
            .O(N__3243),
            .I(N__3240));
    Sp12to4 I__535 (
            .O(N__3240),
            .I(N__3237));
    Span12Mux_v I__534 (
            .O(N__3237),
            .I(N__3234));
    Span12Mux_h I__533 (
            .O(N__3234),
            .I(N__3231));
    Odrv12 I__532 (
            .O(N__3231),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__531 (
            .O(N__3228),
            .I(N__3225));
    LocalMux I__530 (
            .O(N__3225),
            .I(N__3222));
    IoSpan4Mux I__529 (
            .O(N__3222),
            .I(N__3219));
    Span4Mux_s0_h I__528 (
            .O(N__3219),
            .I(N__3216));
    Sp12to4 I__527 (
            .O(N__3216),
            .I(N__3213));
    Span12Mux_s8_h I__526 (
            .O(N__3213),
            .I(N__3210));
    Odrv12 I__525 (
            .O(N__3210),
            .I(un1_D_LM_AMIGA_6));
    CascadeMux I__524 (
            .O(N__3207),
            .I(N__3204));
    InMux I__523 (
            .O(N__3204),
            .I(N__3201));
    LocalMux I__522 (
            .O(N__3201),
            .I(N__3198));
    Odrv12 I__521 (
            .O(N__3198),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__520 (
            .O(N__3195),
            .I(N__3192));
    LocalMux I__519 (
            .O(N__3192),
            .I(N__3189));
    Span4Mux_s2_h I__518 (
            .O(N__3189),
            .I(N__3186));
    Span4Mux_h I__517 (
            .O(N__3186),
            .I(N__3183));
    Sp12to4 I__516 (
            .O(N__3183),
            .I(N__3180));
    Span12Mux_v I__515 (
            .O(N__3180),
            .I(N__3177));
    Span12Mux_h I__514 (
            .O(N__3177),
            .I(N__3174));
    Odrv12 I__513 (
            .O(N__3174),
            .I(un1_D_LM_AMIGA_1));
    InMux I__512 (
            .O(N__3171),
            .I(N__3168));
    LocalMux I__511 (
            .O(N__3168),
            .I(N__3165));
    Span12Mux_v I__510 (
            .O(N__3165),
            .I(N__3162));
    Span12Mux_h I__509 (
            .O(N__3162),
            .I(N__3159));
    Odrv12 I__508 (
            .O(N__3159),
            .I(D_UM_040_in_6));
    IoInMux I__507 (
            .O(N__3156),
            .I(N__3153));
    LocalMux I__506 (
            .O(N__3153),
            .I(N__3150));
    IoSpan4Mux I__505 (
            .O(N__3150),
            .I(N__3146));
    CascadeMux I__504 (
            .O(N__3149),
            .I(N__3143));
    IoSpan4Mux I__503 (
            .O(N__3146),
            .I(N__3140));
    InMux I__502 (
            .O(N__3143),
            .I(N__3137));
    Span4Mux_s2_h I__501 (
            .O(N__3140),
            .I(N__3134));
    LocalMux I__500 (
            .O(N__3137),
            .I(N__3131));
    Sp12to4 I__499 (
            .O(N__3134),
            .I(N__3128));
    Span12Mux_v I__498 (
            .O(N__3131),
            .I(N__3125));
    Span12Mux_h I__497 (
            .O(N__3128),
            .I(N__3122));
    Span12Mux_v I__496 (
            .O(N__3125),
            .I(N__3119));
    Span12Mux_h I__495 (
            .O(N__3122),
            .I(N__3116));
    Span12Mux_h I__494 (
            .O(N__3119),
            .I(N__3113));
    Odrv12 I__493 (
            .O(N__3116),
            .I(D_LL_040_in_6));
    Odrv12 I__492 (
            .O(N__3113),
            .I(D_LL_040_in_6));
    IoInMux I__491 (
            .O(N__3108),
            .I(N__3105));
    LocalMux I__490 (
            .O(N__3105),
            .I(N__3102));
    Span12Mux_s2_h I__489 (
            .O(N__3102),
            .I(N__3099));
    Span12Mux_v I__488 (
            .O(N__3099),
            .I(N__3096));
    Odrv12 I__487 (
            .O(N__3096),
            .I(un1_D_UM_040_6));
    CascadeMux I__486 (
            .O(N__3093),
            .I(N__3090));
    InMux I__485 (
            .O(N__3090),
            .I(N__3087));
    LocalMux I__484 (
            .O(N__3087),
            .I(N__3084));
    Span4Mux_v I__483 (
            .O(N__3084),
            .I(N__3081));
    Sp12to4 I__482 (
            .O(N__3081),
            .I(N__3078));
    Span12Mux_h I__481 (
            .O(N__3078),
            .I(N__3075));
    Span12Mux_h I__480 (
            .O(N__3075),
            .I(N__3072));
    Odrv12 I__479 (
            .O(N__3072),
            .I(D_UM_040_in_4));
    IoInMux I__478 (
            .O(N__3069),
            .I(N__3066));
    LocalMux I__477 (
            .O(N__3066),
            .I(N__3062));
    InMux I__476 (
            .O(N__3065),
            .I(N__3059));
    Span4Mux_s2_h I__475 (
            .O(N__3062),
            .I(N__3056));
    LocalMux I__474 (
            .O(N__3059),
            .I(N__3053));
    Span4Mux_v I__473 (
            .O(N__3056),
            .I(N__3050));
    Span12Mux_v I__472 (
            .O(N__3053),
            .I(N__3047));
    Sp12to4 I__471 (
            .O(N__3050),
            .I(N__3044));
    Span12Mux_v I__470 (
            .O(N__3047),
            .I(N__3041));
    Span12Mux_h I__469 (
            .O(N__3044),
            .I(N__3038));
    Span12Mux_h I__468 (
            .O(N__3041),
            .I(N__3035));
    Span12Mux_h I__467 (
            .O(N__3038),
            .I(N__3032));
    Odrv12 I__466 (
            .O(N__3035),
            .I(D_LL_040_in_4));
    Odrv12 I__465 (
            .O(N__3032),
            .I(D_LL_040_in_4));
    IoInMux I__464 (
            .O(N__3027),
            .I(N__3024));
    LocalMux I__463 (
            .O(N__3024),
            .I(N__3021));
    Span4Mux_s1_h I__462 (
            .O(N__3021),
            .I(N__3018));
    Span4Mux_h I__461 (
            .O(N__3018),
            .I(N__3015));
    Span4Mux_h I__460 (
            .O(N__3015),
            .I(N__3012));
    Odrv4 I__459 (
            .O(N__3012),
            .I(un1_D_UM_040_4));
    InMux I__458 (
            .O(N__3009),
            .I(N__3006));
    LocalMux I__457 (
            .O(N__3006),
            .I(N__3003));
    Span4Mux_v I__456 (
            .O(N__3003),
            .I(N__3000));
    Span4Mux_h I__455 (
            .O(N__3000),
            .I(N__2997));
    Span4Mux_h I__454 (
            .O(N__2997),
            .I(N__2994));
    Sp12to4 I__453 (
            .O(N__2994),
            .I(N__2991));
    Span12Mux_h I__452 (
            .O(N__2991),
            .I(N__2988));
    Odrv12 I__451 (
            .O(N__2988),
            .I(D_UU_040_in_3));
    IoInMux I__450 (
            .O(N__2985),
            .I(N__2982));
    LocalMux I__449 (
            .O(N__2982),
            .I(N__2979));
    IoSpan4Mux I__448 (
            .O(N__2979),
            .I(N__2976));
    IoSpan4Mux I__447 (
            .O(N__2976),
            .I(N__2972));
    InMux I__446 (
            .O(N__2975),
            .I(N__2969));
    Span4Mux_s2_h I__445 (
            .O(N__2972),
            .I(N__2966));
    LocalMux I__444 (
            .O(N__2969),
            .I(N__2963));
    Sp12to4 I__443 (
            .O(N__2966),
            .I(N__2960));
    Span12Mux_s10_v I__442 (
            .O(N__2963),
            .I(N__2957));
    Span12Mux_h I__441 (
            .O(N__2960),
            .I(N__2954));
    Span12Mux_v I__440 (
            .O(N__2957),
            .I(N__2951));
    Span12Mux_h I__439 (
            .O(N__2954),
            .I(N__2948));
    Span12Mux_h I__438 (
            .O(N__2951),
            .I(N__2945));
    Odrv12 I__437 (
            .O(N__2948),
            .I(D_LM_040_in_3));
    Odrv12 I__436 (
            .O(N__2945),
            .I(D_LM_040_in_3));
    IoInMux I__435 (
            .O(N__2940),
            .I(N__2937));
    LocalMux I__434 (
            .O(N__2937),
            .I(N__2934));
    IoSpan4Mux I__433 (
            .O(N__2934),
            .I(N__2931));
    IoSpan4Mux I__432 (
            .O(N__2931),
            .I(N__2928));
    Span4Mux_s2_v I__431 (
            .O(N__2928),
            .I(N__2925));
    Span4Mux_v I__430 (
            .O(N__2925),
            .I(N__2922));
    Odrv4 I__429 (
            .O(N__2922),
            .I(un1_D_UU_040_3));
    IoInMux I__428 (
            .O(N__2919),
            .I(N__2916));
    LocalMux I__427 (
            .O(N__2916),
            .I(N__2913));
    Span4Mux_s2_h I__426 (
            .O(N__2913),
            .I(N__2910));
    Span4Mux_v I__425 (
            .O(N__2910),
            .I(N__2906));
    InMux I__424 (
            .O(N__2909),
            .I(N__2903));
    Sp12to4 I__423 (
            .O(N__2906),
            .I(N__2900));
    LocalMux I__422 (
            .O(N__2903),
            .I(N__2897));
    Span12Mux_h I__421 (
            .O(N__2900),
            .I(N__2894));
    Span12Mux_s11_v I__420 (
            .O(N__2897),
            .I(N__2891));
    Span12Mux_h I__419 (
            .O(N__2894),
            .I(N__2888));
    Span12Mux_h I__418 (
            .O(N__2891),
            .I(N__2885));
    Odrv12 I__417 (
            .O(N__2888),
            .I(D_LM_040_in_6));
    Odrv12 I__416 (
            .O(N__2885),
            .I(D_LM_040_in_6));
    CascadeMux I__415 (
            .O(N__2880),
            .I(N__2877));
    InMux I__414 (
            .O(N__2877),
            .I(N__2874));
    LocalMux I__413 (
            .O(N__2874),
            .I(N__2871));
    Span4Mux_v I__412 (
            .O(N__2871),
            .I(N__2868));
    Sp12to4 I__411 (
            .O(N__2868),
            .I(N__2865));
    Span12Mux_h I__410 (
            .O(N__2865),
            .I(N__2862));
    Span12Mux_h I__409 (
            .O(N__2862),
            .I(N__2859));
    Odrv12 I__408 (
            .O(N__2859),
            .I(D_UU_040_in_6));
    IoInMux I__407 (
            .O(N__2856),
            .I(N__2853));
    LocalMux I__406 (
            .O(N__2853),
            .I(N__2850));
    IoSpan4Mux I__405 (
            .O(N__2850),
            .I(N__2847));
    Span4Mux_s2_v I__404 (
            .O(N__2847),
            .I(N__2844));
    Span4Mux_v I__403 (
            .O(N__2844),
            .I(N__2841));
    Odrv4 I__402 (
            .O(N__2841),
            .I(un1_D_UU_040_6));
    InMux I__401 (
            .O(N__2838),
            .I(N__2835));
    LocalMux I__400 (
            .O(N__2835),
            .I(N__2832));
    Span4Mux_v I__399 (
            .O(N__2832),
            .I(N__2829));
    Sp12to4 I__398 (
            .O(N__2829),
            .I(N__2826));
    Odrv12 I__397 (
            .O(N__2826),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__396 (
            .O(N__2823),
            .I(N__2820));
    LocalMux I__395 (
            .O(N__2820),
            .I(N__2817));
    IoSpan4Mux I__394 (
            .O(N__2817),
            .I(N__2814));
    Sp12to4 I__393 (
            .O(N__2814),
            .I(N__2811));
    Span12Mux_s9_h I__392 (
            .O(N__2811),
            .I(N__2808));
    Span12Mux_h I__391 (
            .O(N__2808),
            .I(N__2805));
    Odrv12 I__390 (
            .O(N__2805),
            .I(un1_D_LL_AMIGA_7));
    IoInMux I__389 (
            .O(N__2802),
            .I(N__2798));
    InMux I__388 (
            .O(N__2801),
            .I(N__2795));
    LocalMux I__387 (
            .O(N__2798),
            .I(N__2792));
    LocalMux I__386 (
            .O(N__2795),
            .I(N__2789));
    Span4Mux_s3_h I__385 (
            .O(N__2792),
            .I(N__2786));
    Sp12to4 I__384 (
            .O(N__2789),
            .I(N__2783));
    Sp12to4 I__383 (
            .O(N__2786),
            .I(N__2780));
    Span12Mux_v I__382 (
            .O(N__2783),
            .I(N__2777));
    Span12Mux_v I__381 (
            .O(N__2780),
            .I(N__2774));
    Span12Mux_v I__380 (
            .O(N__2777),
            .I(N__2771));
    Span12Mux_h I__379 (
            .O(N__2774),
            .I(N__2768));
    Span12Mux_h I__378 (
            .O(N__2771),
            .I(N__2765));
    Span12Mux_h I__377 (
            .O(N__2768),
            .I(N__2762));
    Odrv12 I__376 (
            .O(N__2765),
            .I(D_LL_040_in_1));
    Odrv12 I__375 (
            .O(N__2762),
            .I(D_LL_040_in_1));
    InMux I__374 (
            .O(N__2757),
            .I(N__2754));
    LocalMux I__373 (
            .O(N__2754),
            .I(N__2751));
    Span4Mux_h I__372 (
            .O(N__2751),
            .I(N__2748));
    Sp12to4 I__371 (
            .O(N__2748),
            .I(N__2745));
    Span12Mux_v I__370 (
            .O(N__2745),
            .I(N__2742));
    Span12Mux_h I__369 (
            .O(N__2742),
            .I(N__2739));
    Odrv12 I__368 (
            .O(N__2739),
            .I(D_UM_040_in_1));
    IoInMux I__367 (
            .O(N__2736),
            .I(N__2733));
    LocalMux I__366 (
            .O(N__2733),
            .I(N__2730));
    IoSpan4Mux I__365 (
            .O(N__2730),
            .I(N__2727));
    Sp12to4 I__364 (
            .O(N__2727),
            .I(N__2724));
    Odrv12 I__363 (
            .O(N__2724),
            .I(un1_D_UM_040_1));
    InMux I__362 (
            .O(N__2721),
            .I(N__2718));
    LocalMux I__361 (
            .O(N__2718),
            .I(N__2715));
    Span4Mux_v I__360 (
            .O(N__2715),
            .I(N__2712));
    Span4Mux_h I__359 (
            .O(N__2712),
            .I(N__2709));
    Sp12to4 I__358 (
            .O(N__2709),
            .I(N__2706));
    Span12Mux_h I__357 (
            .O(N__2706),
            .I(N__2703));
    Odrv12 I__356 (
            .O(N__2703),
            .I(D_UU_040_in_7));
    IoInMux I__355 (
            .O(N__2700),
            .I(N__2697));
    LocalMux I__354 (
            .O(N__2697),
            .I(N__2693));
    CascadeMux I__353 (
            .O(N__2696),
            .I(N__2690));
    IoSpan4Mux I__352 (
            .O(N__2693),
            .I(N__2687));
    InMux I__351 (
            .O(N__2690),
            .I(N__2684));
    Span4Mux_s2_h I__350 (
            .O(N__2687),
            .I(N__2681));
    LocalMux I__349 (
            .O(N__2684),
            .I(N__2678));
    Sp12to4 I__348 (
            .O(N__2681),
            .I(N__2675));
    Span4Mux_v I__347 (
            .O(N__2678),
            .I(N__2672));
    Span12Mux_h I__346 (
            .O(N__2675),
            .I(N__2669));
    Sp12to4 I__345 (
            .O(N__2672),
            .I(N__2666));
    Span12Mux_h I__344 (
            .O(N__2669),
            .I(N__2663));
    Span12Mux_h I__343 (
            .O(N__2666),
            .I(N__2660));
    Odrv12 I__342 (
            .O(N__2663),
            .I(D_LM_040_in_7));
    Odrv12 I__341 (
            .O(N__2660),
            .I(D_LM_040_in_7));
    IoInMux I__340 (
            .O(N__2655),
            .I(N__2652));
    LocalMux I__339 (
            .O(N__2652),
            .I(N__2649));
    IoSpan4Mux I__338 (
            .O(N__2649),
            .I(N__2646));
    Sp12to4 I__337 (
            .O(N__2646),
            .I(N__2643));
    Span12Mux_s6_v I__336 (
            .O(N__2643),
            .I(N__2640));
    Odrv12 I__335 (
            .O(N__2640),
            .I(un1_D_UU_040_7));
    InMux I__334 (
            .O(N__2637),
            .I(N__2634));
    LocalMux I__333 (
            .O(N__2634),
            .I(N__2631));
    Span4Mux_h I__332 (
            .O(N__2631),
            .I(N__2628));
    Span4Mux_v I__331 (
            .O(N__2628),
            .I(N__2625));
    Odrv4 I__330 (
            .O(N__2625),
            .I(A_040_c_0));
    IoInMux I__329 (
            .O(N__2622),
            .I(N__2619));
    LocalMux I__328 (
            .O(N__2619),
            .I(N__2616));
    Span4Mux_s2_v I__327 (
            .O(N__2616),
            .I(N__2613));
    Span4Mux_v I__326 (
            .O(N__2613),
            .I(N__2610));
    Odrv4 I__325 (
            .O(N__2610),
            .I(A_AMIGA_c_0));
    InMux I__324 (
            .O(N__2607),
            .I(N__2604));
    LocalMux I__323 (
            .O(N__2604),
            .I(N__2601));
    Span12Mux_h I__322 (
            .O(N__2601),
            .I(N__2598));
    Odrv12 I__321 (
            .O(N__2598),
            .I(A_040_c_1));
    InMux I__320 (
            .O(N__2595),
            .I(N__2592));
    LocalMux I__319 (
            .O(N__2592),
            .I(N__2589));
    Span12Mux_v I__318 (
            .O(N__2589),
            .I(N__2586));
    Odrv12 I__317 (
            .O(N__2586),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__316 (
            .O(N__2583),
            .I(N__2580));
    LocalMux I__315 (
            .O(N__2580),
            .I(N__2577));
    IoSpan4Mux I__314 (
            .O(N__2577),
            .I(N__2574));
    IoSpan4Mux I__313 (
            .O(N__2574),
            .I(N__2571));
    Span4Mux_s3_h I__312 (
            .O(N__2571),
            .I(N__2568));
    Sp12to4 I__311 (
            .O(N__2568),
            .I(N__2565));
    Span12Mux_s11_h I__310 (
            .O(N__2565),
            .I(N__2562));
    Odrv12 I__309 (
            .O(N__2562),
            .I(un1_D_LL_AMIGA_2));
    IoInMux I__308 (
            .O(N__2559),
            .I(N__2552));
    IoInMux I__307 (
            .O(N__2558),
            .I(N__2549));
    IoInMux I__306 (
            .O(N__2557),
            .I(N__2546));
    IoInMux I__305 (
            .O(N__2556),
            .I(N__2539));
    IoInMux I__304 (
            .O(N__2555),
            .I(N__2536));
    LocalMux I__303 (
            .O(N__2552),
            .I(N__2527));
    LocalMux I__302 (
            .O(N__2549),
            .I(N__2527));
    LocalMux I__301 (
            .O(N__2546),
            .I(N__2527));
    IoInMux I__300 (
            .O(N__2545),
            .I(N__2524));
    IoInMux I__299 (
            .O(N__2544),
            .I(N__2521));
    IoInMux I__298 (
            .O(N__2543),
            .I(N__2518));
    IoInMux I__297 (
            .O(N__2542),
            .I(N__2515));
    LocalMux I__296 (
            .O(N__2539),
            .I(N__2503));
    LocalMux I__295 (
            .O(N__2536),
            .I(N__2503));
    IoInMux I__294 (
            .O(N__2535),
            .I(N__2500));
    IoInMux I__293 (
            .O(N__2534),
            .I(N__2497));
    IoSpan4Mux I__292 (
            .O(N__2527),
            .I(N__2486));
    LocalMux I__291 (
            .O(N__2524),
            .I(N__2486));
    LocalMux I__290 (
            .O(N__2521),
            .I(N__2486));
    LocalMux I__289 (
            .O(N__2518),
            .I(N__2486));
    LocalMux I__288 (
            .O(N__2515),
            .I(N__2486));
    IoInMux I__287 (
            .O(N__2514),
            .I(N__2483));
    IoInMux I__286 (
            .O(N__2513),
            .I(N__2480));
    IoInMux I__285 (
            .O(N__2512),
            .I(N__2477));
    IoInMux I__284 (
            .O(N__2511),
            .I(N__2474));
    IoInMux I__283 (
            .O(N__2510),
            .I(N__2467));
    IoInMux I__282 (
            .O(N__2509),
            .I(N__2464));
    IoInMux I__281 (
            .O(N__2508),
            .I(N__2461));
    IoSpan4Mux I__280 (
            .O(N__2503),
            .I(N__2454));
    LocalMux I__279 (
            .O(N__2500),
            .I(N__2454));
    LocalMux I__278 (
            .O(N__2497),
            .I(N__2451));
    IoSpan4Mux I__277 (
            .O(N__2486),
            .I(N__2440));
    LocalMux I__276 (
            .O(N__2483),
            .I(N__2440));
    LocalMux I__275 (
            .O(N__2480),
            .I(N__2440));
    LocalMux I__274 (
            .O(N__2477),
            .I(N__2440));
    LocalMux I__273 (
            .O(N__2474),
            .I(N__2440));
    IoInMux I__272 (
            .O(N__2473),
            .I(N__2437));
    IoInMux I__271 (
            .O(N__2472),
            .I(N__2434));
    IoInMux I__270 (
            .O(N__2471),
            .I(N__2431));
    IoInMux I__269 (
            .O(N__2470),
            .I(N__2428));
    LocalMux I__268 (
            .O(N__2467),
            .I(N__2423));
    LocalMux I__267 (
            .O(N__2464),
            .I(N__2418));
    LocalMux I__266 (
            .O(N__2461),
            .I(N__2418));
    IoInMux I__265 (
            .O(N__2460),
            .I(N__2415));
    IoInMux I__264 (
            .O(N__2459),
            .I(N__2412));
    Span4Mux_s3_v I__263 (
            .O(N__2454),
            .I(N__2403));
    Span4Mux_s3_v I__262 (
            .O(N__2451),
            .I(N__2400));
    IoSpan4Mux I__261 (
            .O(N__2440),
            .I(N__2389));
    LocalMux I__260 (
            .O(N__2437),
            .I(N__2389));
    LocalMux I__259 (
            .O(N__2434),
            .I(N__2389));
    LocalMux I__258 (
            .O(N__2431),
            .I(N__2389));
    LocalMux I__257 (
            .O(N__2428),
            .I(N__2389));
    IoInMux I__256 (
            .O(N__2427),
            .I(N__2386));
    IoInMux I__255 (
            .O(N__2426),
            .I(N__2383));
    IoSpan4Mux I__254 (
            .O(N__2423),
            .I(N__2374));
    IoSpan4Mux I__253 (
            .O(N__2418),
            .I(N__2374));
    LocalMux I__252 (
            .O(N__2415),
            .I(N__2374));
    LocalMux I__251 (
            .O(N__2412),
            .I(N__2374));
    IoInMux I__250 (
            .O(N__2411),
            .I(N__2371));
    IoInMux I__249 (
            .O(N__2410),
            .I(N__2368));
    IoInMux I__248 (
            .O(N__2409),
            .I(N__2365));
    IoInMux I__247 (
            .O(N__2408),
            .I(N__2362));
    IoInMux I__246 (
            .O(N__2407),
            .I(N__2359));
    IoInMux I__245 (
            .O(N__2406),
            .I(N__2356));
    Span4Mux_v I__244 (
            .O(N__2403),
            .I(N__2353));
    Span4Mux_v I__243 (
            .O(N__2400),
            .I(N__2350));
    IoSpan4Mux I__242 (
            .O(N__2389),
            .I(N__2343));
    LocalMux I__241 (
            .O(N__2386),
            .I(N__2343));
    LocalMux I__240 (
            .O(N__2383),
            .I(N__2343));
    IoSpan4Mux I__239 (
            .O(N__2374),
            .I(N__2332));
    LocalMux I__238 (
            .O(N__2371),
            .I(N__2332));
    LocalMux I__237 (
            .O(N__2368),
            .I(N__2332));
    LocalMux I__236 (
            .O(N__2365),
            .I(N__2332));
    LocalMux I__235 (
            .O(N__2362),
            .I(N__2332));
    LocalMux I__234 (
            .O(N__2359),
            .I(N__2327));
    LocalMux I__233 (
            .O(N__2356),
            .I(N__2327));
    Sp12to4 I__232 (
            .O(N__2353),
            .I(N__2322));
    Sp12to4 I__231 (
            .O(N__2350),
            .I(N__2322));
    IoSpan4Mux I__230 (
            .O(N__2343),
            .I(N__2317));
    IoSpan4Mux I__229 (
            .O(N__2332),
            .I(N__2317));
    Span12Mux_s7_v I__228 (
            .O(N__2327),
            .I(N__2312));
    Span12Mux_h I__227 (
            .O(N__2322),
            .I(N__2312));
    Span4Mux_s3_h I__226 (
            .O(N__2317),
            .I(N__2309));
    Span12Mux_v I__225 (
            .O(N__2312),
            .I(N__2306));
    Span4Mux_h I__224 (
            .O(N__2309),
            .I(N__2303));
    Odrv12 I__223 (
            .O(N__2306),
            .I(RnW_c_i_0));
    Odrv4 I__222 (
            .O(N__2303),
            .I(RnW_c_i_0));
    InMux I__221 (
            .O(N__2298),
            .I(N__2295));
    LocalMux I__220 (
            .O(N__2295),
            .I(N__2292));
    Span12Mux_h I__219 (
            .O(N__2292),
            .I(N__2289));
    Span12Mux_h I__218 (
            .O(N__2289),
            .I(N__2286));
    Odrv12 I__217 (
            .O(N__2286),
            .I(D_UM_040_in_0));
    IoInMux I__216 (
            .O(N__2283),
            .I(N__2279));
    CascadeMux I__215 (
            .O(N__2282),
            .I(N__2276));
    LocalMux I__214 (
            .O(N__2279),
            .I(N__2273));
    InMux I__213 (
            .O(N__2276),
            .I(N__2270));
    IoSpan4Mux I__212 (
            .O(N__2273),
            .I(N__2267));
    LocalMux I__211 (
            .O(N__2270),
            .I(N__2264));
    Span4Mux_s2_h I__210 (
            .O(N__2267),
            .I(N__2261));
    Span12Mux_v I__209 (
            .O(N__2264),
            .I(N__2258));
    Sp12to4 I__208 (
            .O(N__2261),
            .I(N__2255));
    Span12Mux_v I__207 (
            .O(N__2258),
            .I(N__2252));
    Span12Mux_h I__206 (
            .O(N__2255),
            .I(N__2249));
    Span12Mux_h I__205 (
            .O(N__2252),
            .I(N__2246));
    Span12Mux_h I__204 (
            .O(N__2249),
            .I(N__2243));
    Odrv12 I__203 (
            .O(N__2246),
            .I(D_LL_040_in_0));
    Odrv12 I__202 (
            .O(N__2243),
            .I(D_LL_040_in_0));
    IoInMux I__201 (
            .O(N__2238),
            .I(N__2235));
    LocalMux I__200 (
            .O(N__2235),
            .I(N__2232));
    Span4Mux_s1_h I__199 (
            .O(N__2232),
            .I(N__2229));
    Span4Mux_h I__198 (
            .O(N__2229),
            .I(N__2226));
    Span4Mux_h I__197 (
            .O(N__2226),
            .I(N__2223));
    Odrv4 I__196 (
            .O(N__2223),
            .I(un1_D_UM_040_0));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .I(N__6227));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ),
            .I(N__6231));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .I(N__6224));
    INV \INVU111_CYCLE_SM.LW_CYCLEC  (
            .O(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .I(N__6225));
    INV \INVU111_CYCLE_SM.CYCLE_STATE_0C  (
            .O(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .I(N__6228));
    INV \INVU111_CYCLE_SM.TS_ENC  (
            .O(\INVU111_CYCLE_SM.TS_ENC_net ),
            .I(N__6229));
    INV \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C  (
            .O(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .I(N__6226));
    INV \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C  (
            .O(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .I(N__6230));
    INV \INVU111_CYCLE_SM.A_OUTC  (
            .O(\INVU111_CYCLE_SM.A_OUTC_net ),
            .I(N__6232));
    INV \INVU111_CYCLE_SM.TA_ENC  (
            .O(\INVU111_CYCLE_SM.TA_ENC_net ),
            .I(N__6233));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__6075));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_2 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_2  (
            .in0(N__2637),
            .in1(N__7479),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_6  (
            .in0(N__2607),
            .in1(N__7478),
            .in2(_gnd_net_),
            .in3(N__4134),
            .lcout(A_AMIGA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_6_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_6_3_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_6_3_5  (
            .in0(N__4363),
            .in1(N__5386),
            .in2(N__6445),
            .in3(N__2595),
            .lcout(un1_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RnW_c_sbtinv_LC_6_7_0.C_ON=1'b0;
    defparam RnW_c_sbtinv_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam RnW_c_sbtinv_LC_6_7_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RnW_c_sbtinv_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5981),
            .lcout(RnW_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_6_9_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_6_9_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_6_9_2  (
            .in0(N__2298),
            .in1(N__5352),
            .in2(N__2282),
            .in3(N__4409),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_6_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_6_10_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_6_10_4  (
            .in0(N__5337),
            .in1(N__7113),
            .in2(N__3207),
            .in3(N__4452),
            .lcout(un1_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_6_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_6_12_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_6_12_3  (
            .in0(N__5368),
            .in1(N__3171),
            .in2(N__3149),
            .in3(N__4453),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_6_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_6_19_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_6_19_2  (
            .in0(N__4449),
            .in1(N__5380),
            .in2(N__3093),
            .in3(N__3065),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_0  (
            .in0(N__5387),
            .in1(N__3009),
            .in2(N__4554),
            .in3(N__2975),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_6_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_6_20_7 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_6_20_7  (
            .in0(N__2909),
            .in1(N__5388),
            .in2(N__2880),
            .in3(N__4525),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_5 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_5  (
            .in0(N__2838),
            .in1(N__5338),
            .in2(N__6776),
            .in3(N__4466),
            .lcout(un1_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_7_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_7_15_6 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_7_15_6  (
            .in0(N__2801),
            .in1(N__5356),
            .in2(N__4560),
            .in3(N__2757),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_7_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_7_20_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_7_20_1  (
            .in0(N__5373),
            .in1(N__2721),
            .in2(N__2696),
            .in3(N__4561),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_0  (
            .in0(N__5374),
            .in1(N__6684),
            .in2(N__3588),
            .in3(N__4427),
            .lcout(un1_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_1  (
            .in0(N__4503),
            .in1(N__5268),
            .in2(N__3549),
            .in3(N__3530),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_8_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_8_11_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_8_11_1  (
            .in0(N__4504),
            .in1(N__5228),
            .in2(N__6540),
            .in3(N__3471),
            .lcout(un1_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_8_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_8_15_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_8_15_2  (
            .in0(N__3438),
            .in1(N__5309),
            .in2(N__6609),
            .in3(N__4539),
            .lcout(un1_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_1 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_1  (
            .in0(N__4562),
            .in1(N__5379),
            .in2(N__3405),
            .in3(N__3371),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_9_1_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_9_1_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_9_1_1  (
            .in0(N__4341),
            .in1(N__5372),
            .in2(N__4104),
            .in3(N__3330),
            .lcout(un1_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_9_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_9_1_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__5601),
            .in2(_gnd_net_),
            .in3(N__5055),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_9_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_9_12_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_9_12_3  (
            .in0(N__5307),
            .in1(N__3276),
            .in2(N__5544),
            .in3(N__4492),
            .lcout(un1_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_14_5 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_14_5  (
            .in0(N__3246),
            .in1(N__5308),
            .in2(N__4251),
            .in3(N__4526),
            .lcout(un1_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_2 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_2  (
            .in0(N__5344),
            .in1(N__4008),
            .in2(N__4566),
            .in3(N__3986),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_0  (
            .in0(N__4559),
            .in1(N__5378),
            .in2(N__3927),
            .in3(N__3906),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_10_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_10_6_6 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_10_6_6  (
            .in0(N__6051),
            .in1(N__5348),
            .in2(N__3846),
            .in3(N__4457),
            .lcout(un1_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_10_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNO_0_LC_10_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNO_0_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5609),
            .lcout(\U111_CYCLE_SM.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_18_1 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_18_1  (
            .in0(N__5343),
            .in1(N__3801),
            .in2(N__3756),
            .in3(N__4558),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_11_2_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_11_2_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_11_2_4  (
            .in0(N__5367),
            .in1(N__3711),
            .in2(N__6861),
            .in3(N__4439),
            .lcout(un1_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_2_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_2_5 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_2_5  (
            .in0(N__4438),
            .in1(N__5366),
            .in2(N__6135),
            .in3(N__3672),
            .lcout(un1_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_2 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_2  (
            .in0(N__5322),
            .in1(N__7038),
            .in2(N__3633),
            .in3(N__4481),
            .lcout(un1_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_11_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_11_6_6 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_11_6_6  (
            .in0(N__5321),
            .in1(N__4188),
            .in2(N__7185),
            .in3(N__4480),
            .lcout(un1_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_11_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_11_9_0  (
            .in0(N__7461),
            .in1(N__4059),
            .in2(_gnd_net_),
            .in3(N__4094),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_LC_11_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_LC_11_10_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TA_EN_LC_11_10_1 .LUT_INIT=16'b1111000011011100;
    LogicCell40 \U111_CYCLE_SM.TA_EN_LC_11_10_1  (
            .in0(N__5680),
            .in1(N__6399),
            .in2(N__5445),
            .in3(N__6291),
            .lcout(\U111_CYCLE_SM.TA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TA_ENC_net ),
            .ce(),
            .sr(N__4143));
    defparam \U111_CYCLE_SM.A_OUT_LC_11_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A_OUT_LC_11_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.A_OUT_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__5643),
            .in2(_gnd_net_),
            .in3(N__4110),
            .lcout(\U111_CYCLE_SM.A_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.A_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_11_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A_OUT_RNO_0_LC_11_11_7 .LUT_INIT=16'b1010101011001110;
    LogicCell40 \U111_CYCLE_SM.A_OUT_RNO_0_LC_11_11_7  (
            .in0(N__4121),
            .in1(N__6392),
            .in2(N__5682),
            .in3(N__6284),
            .lcout(\U111_CYCLE_SM.A_OUT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_4  (
            .in0(N__6040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__7272),
            .sr(N__7243));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_11_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4081),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net ),
            .ce(N__7272),
            .sr(N__7243));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_1 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_1  (
            .in0(N__4050),
            .in1(N__5198),
            .in2(N__6951),
            .in3(N__4448),
            .lcout(un1_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_2  (
            .in0(N__5540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7273),
            .sr(N__7236));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_4  (
            .in0(N__4247),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net ),
            .ce(N__7273),
            .sr(N__7236));
    defparam CONSTANT_ONE_LUT4_LC_11_16_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_16_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_11_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_11_16_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_11_16_4  (
            .in0(N__5275),
            .in1(N__7335),
            .in2(N__4563),
            .in3(N__4938),
            .lcout(un1_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_11_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_11_19_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_11_19_3  (
            .in0(N__4450),
            .in1(N__5339),
            .in2(N__4899),
            .in3(N__4868),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_19_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_19_4  (
            .in0(N__5340),
            .in1(N__4815),
            .in2(N__4796),
            .in3(N__4451),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_1  (
            .in0(N__4565),
            .in1(N__5342),
            .in2(N__4724),
            .in3(N__4680),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_11_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_11_20_4 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_11_20_4  (
            .in0(N__5341),
            .in1(N__4638),
            .in2(N__4613),
            .in3(N__4564),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_5  (
            .in0(N__4263),
            .in1(N__4240),
            .in2(_gnd_net_),
            .in3(N__7467),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_7  (
            .in0(N__5556),
            .in1(N__5527),
            .in2(_gnd_net_),
            .in3(N__7466),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_1.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6090),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_10_3 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_10_3  (
            .in0(N__5444),
            .in1(N__6341),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(U111_CYCLE_SM_TAn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_12_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_12_11_0 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_12_11_0  (
            .in0(N__5010),
            .in1(N__5004),
            .in2(N__5644),
            .in3(N__5048),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TS_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_12_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_12_11_3 .LUT_INIT=16'b0000101100000111;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_12_11_3  (
            .in0(N__5093),
            .in1(N__5111),
            .in2(N__7460),
            .in3(N__5072),
            .lcout(\U111_CYCLE_SM.un1_LW_TRANS_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_12_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_12_11_4 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_12_11_4  (
            .in0(N__5112),
            .in1(N__5094),
            .in2(N__5076),
            .in3(N__5047),
            .lcout(),
            .ltout(\U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_12_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_START_LC_12_11_5 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_START_LC_12_11_5  (
            .in0(N__7419),
            .in1(N__5631),
            .in2(N__5031),
            .in3(N__5679),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TS_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_11_6 .LUT_INIT=16'b0101001101010000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_11_6  (
            .in0(N__6283),
            .in1(N__5028),
            .in2(N__6398),
            .in3(N__6088),
            .lcout(\U111_CYCLE_SM.TS_EN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_11_7 .LUT_INIT=16'b1100110010111011;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_11_7  (
            .in0(N__6087),
            .in1(N__6388),
            .in2(_gnd_net_),
            .in3(N__6282),
            .lcout(\U111_CYCLE_SM.N_69_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_12_0  (
            .in0(N__5678),
            .in1(N__6089),
            .in2(_gnd_net_),
            .in3(N__6393),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_12_1 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_12_1  (
            .in0(N__5635),
            .in1(N__6342),
            .in2(N__6054),
            .in3(N__6288),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_12_2 .LUT_INIT=16'b1100010000001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_12_2  (
            .in0(N__6289),
            .in1(N__5636),
            .in2(N__6350),
            .in3(N__6394),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.CYCLE_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_3 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_3  (
            .in0(N__6041),
            .in1(N__6015),
            .in2(N__7424),
            .in3(_gnd_net_),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_0 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__6346),
            .in2(N__6290),
            .in3(N__6385),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_1 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_1  (
            .in0(N__5645),
            .in1(_gnd_net_),
            .in2(N__5988),
            .in3(N__5904),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0 ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5691),
            .in3(N__5688),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_13_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__5681),
            .in2(_gnd_net_),
            .in3(N__6280),
            .lcout(),
            .ltout(\U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_CYCLE_LC_12_13_4 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_LC_12_13_4  (
            .in0(N__5646),
            .in1(N__6243),
            .in2(N__6402),
            .in3(N__6387),
            .lcout(\U111_CYCLE_SM.LW_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.LW_CYCLEC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_13_5 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_13_5  (
            .in0(N__6386),
            .in1(N__7383),
            .in2(N__6351),
            .in3(N__6281),
            .lcout(\U111_CYCLE_SM.LW_CYCLE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_12_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_12_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6854),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_1  (
            .in0(N__6674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_12_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_12_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_12_14_3  (
            .in0(N__6533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_14_4  (
            .in0(N__6128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_14_5  (
            .in0(N__6777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6608),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net ),
            .ce(N__7271),
            .sr(N__7232));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_1.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_1 (
            .in0(N__6237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_12_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_12_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_12_15_3  (
            .in0(N__7425),
            .in1(N__6141),
            .in2(_gnd_net_),
            .in3(N__6127),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_12_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_12_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_12_16_3  (
            .in0(N__6853),
            .in1(N__6810),
            .in2(_gnd_net_),
            .in3(N__7426),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_19_2  (
            .in0(N__6766),
            .in1(N__6726),
            .in2(_gnd_net_),
            .in3(N__7463),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_4  (
            .in0(N__6693),
            .in1(N__6662),
            .in2(_gnd_net_),
            .in3(N__7462),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_20_1  (
            .in0(N__7465),
            .in1(N__6618),
            .in2(_gnd_net_),
            .in3(N__6595),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_12_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_12_20_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_12_20_4  (
            .in0(N__6526),
            .in1(N__7464),
            .in2(_gnd_net_),
            .in3(N__6495),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_11_4  (
            .in0(N__6447),
            .in1(N__6408),
            .in2(_gnd_net_),
            .in3(N__7423),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_3  (
            .in0(N__6446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net ),
            .ce(N__7274),
            .sr(N__7244));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_0  (
            .in0(N__7034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .ce(N__7275),
            .sr(N__7245));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1  (
            .in0(N__7109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .ce(N__7275),
            .sr(N__7245));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_13_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_13_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_13_14_3  (
            .in0(N__6950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .ce(N__7275),
            .sr(N__7245));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7334),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .ce(N__7275),
            .sr(N__7245));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_13_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7178),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net ),
            .ce(N__7275),
            .sr(N__7245));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_13_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_13_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_13_18_1  (
            .in0(N__7469),
            .in1(N__7194),
            .in2(_gnd_net_),
            .in3(N__7171),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4  (
            .in0(N__7102),
            .in1(N__7068),
            .in2(_gnd_net_),
            .in3(N__7468),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_0  (
            .in0(N__7030),
            .in1(N__6990),
            .in2(_gnd_net_),
            .in3(N__7470),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_13_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_13_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_13_20_3  (
            .in0(N__7471),
            .in1(N__6960),
            .in2(_gnd_net_),
            .in3(N__6946),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7  (
            .in0(N__7472),
            .in1(N__7344),
            .in2(_gnd_net_),
            .in3(N__7327),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

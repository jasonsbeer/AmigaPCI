// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 13 2025 21:12:32

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    TBIn,
    RAMSPACEn,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    PRnW,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    BLSn,
    TCIn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    output TBIn;
    input RAMSPACEn;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output PRnW;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output BLSn;
    output TCIn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12850;
    wire N__12849;
    wire N__12848;
    wire N__12841;
    wire N__12840;
    wire N__12839;
    wire N__12832;
    wire N__12831;
    wire N__12830;
    wire N__12823;
    wire N__12822;
    wire N__12821;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12787;
    wire N__12786;
    wire N__12785;
    wire N__12778;
    wire N__12777;
    wire N__12776;
    wire N__12769;
    wire N__12768;
    wire N__12767;
    wire N__12760;
    wire N__12759;
    wire N__12758;
    wire N__12751;
    wire N__12750;
    wire N__12749;
    wire N__12742;
    wire N__12741;
    wire N__12740;
    wire N__12733;
    wire N__12732;
    wire N__12731;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12715;
    wire N__12714;
    wire N__12713;
    wire N__12706;
    wire N__12705;
    wire N__12704;
    wire N__12697;
    wire N__12696;
    wire N__12695;
    wire N__12688;
    wire N__12687;
    wire N__12686;
    wire N__12679;
    wire N__12678;
    wire N__12677;
    wire N__12670;
    wire N__12669;
    wire N__12668;
    wire N__12661;
    wire N__12660;
    wire N__12659;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12634;
    wire N__12633;
    wire N__12632;
    wire N__12625;
    wire N__12624;
    wire N__12623;
    wire N__12616;
    wire N__12615;
    wire N__12614;
    wire N__12607;
    wire N__12606;
    wire N__12605;
    wire N__12598;
    wire N__12597;
    wire N__12596;
    wire N__12589;
    wire N__12588;
    wire N__12587;
    wire N__12580;
    wire N__12579;
    wire N__12578;
    wire N__12571;
    wire N__12570;
    wire N__12569;
    wire N__12562;
    wire N__12561;
    wire N__12560;
    wire N__12553;
    wire N__12552;
    wire N__12551;
    wire N__12544;
    wire N__12543;
    wire N__12542;
    wire N__12535;
    wire N__12534;
    wire N__12533;
    wire N__12526;
    wire N__12525;
    wire N__12524;
    wire N__12517;
    wire N__12516;
    wire N__12515;
    wire N__12508;
    wire N__12507;
    wire N__12506;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12490;
    wire N__12489;
    wire N__12488;
    wire N__12481;
    wire N__12480;
    wire N__12479;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12463;
    wire N__12462;
    wire N__12461;
    wire N__12454;
    wire N__12453;
    wire N__12452;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12436;
    wire N__12435;
    wire N__12434;
    wire N__12427;
    wire N__12426;
    wire N__12425;
    wire N__12418;
    wire N__12417;
    wire N__12416;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12400;
    wire N__12399;
    wire N__12398;
    wire N__12391;
    wire N__12390;
    wire N__12389;
    wire N__12382;
    wire N__12381;
    wire N__12380;
    wire N__12373;
    wire N__12372;
    wire N__12371;
    wire N__12364;
    wire N__12363;
    wire N__12362;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12346;
    wire N__12345;
    wire N__12344;
    wire N__12337;
    wire N__12336;
    wire N__12335;
    wire N__12328;
    wire N__12327;
    wire N__12326;
    wire N__12319;
    wire N__12318;
    wire N__12317;
    wire N__12310;
    wire N__12309;
    wire N__12308;
    wire N__12301;
    wire N__12300;
    wire N__12299;
    wire N__12292;
    wire N__12291;
    wire N__12290;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12274;
    wire N__12273;
    wire N__12272;
    wire N__12265;
    wire N__12264;
    wire N__12263;
    wire N__12256;
    wire N__12255;
    wire N__12254;
    wire N__12247;
    wire N__12246;
    wire N__12245;
    wire N__12238;
    wire N__12237;
    wire N__12236;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12220;
    wire N__12219;
    wire N__12218;
    wire N__12211;
    wire N__12210;
    wire N__12209;
    wire N__12202;
    wire N__12201;
    wire N__12200;
    wire N__12193;
    wire N__12192;
    wire N__12191;
    wire N__12184;
    wire N__12183;
    wire N__12182;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12157;
    wire N__12156;
    wire N__12155;
    wire N__12148;
    wire N__12147;
    wire N__12146;
    wire N__12139;
    wire N__12138;
    wire N__12137;
    wire N__12130;
    wire N__12129;
    wire N__12128;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12076;
    wire N__12075;
    wire N__12074;
    wire N__12067;
    wire N__12066;
    wire N__12065;
    wire N__12058;
    wire N__12057;
    wire N__12056;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12040;
    wire N__12039;
    wire N__12038;
    wire N__12031;
    wire N__12030;
    wire N__12029;
    wire N__12022;
    wire N__12021;
    wire N__12020;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11986;
    wire N__11985;
    wire N__11984;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11907;
    wire N__11906;
    wire N__11905;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11894;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11860;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11848;
    wire N__11845;
    wire N__11840;
    wire N__11839;
    wire N__11832;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11814;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11799;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11779;
    wire N__11776;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11724;
    wire N__11721;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11706;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11690;
    wire N__11689;
    wire N__11684;
    wire N__11681;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11669;
    wire N__11666;
    wire N__11665;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11650;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11638;
    wire N__11633;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11621;
    wire N__11616;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11592;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11575;
    wire N__11570;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11537;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11511;
    wire N__11508;
    wire N__11503;
    wire N__11500;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11481;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11465;
    wire N__11462;
    wire N__11457;
    wire N__11454;
    wire N__11453;
    wire N__11448;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11357;
    wire N__11352;
    wire N__11351;
    wire N__11350;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11328;
    wire N__11323;
    wire N__11318;
    wire N__11315;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11260;
    wire N__11255;
    wire N__11252;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11209;
    wire N__11202;
    wire N__11199;
    wire N__11198;
    wire N__11195;
    wire N__11194;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11142;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11126;
    wire N__11123;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11111;
    wire N__11108;
    wire N__11101;
    wire N__11098;
    wire N__11097;
    wire N__11094;
    wire N__11089;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11042;
    wire N__11039;
    wire N__11038;
    wire N__11037;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11020;
    wire N__11019;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__11011;
    wire N__11010;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11002;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10994;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10963;
    wire N__10960;
    wire N__10955;
    wire N__10950;
    wire N__10947;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10919;
    wire N__10918;
    wire N__10915;
    wire N__10904;
    wire N__10899;
    wire N__10896;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10868;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10831;
    wire N__10828;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10786;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10759;
    wire N__10758;
    wire N__10757;
    wire N__10756;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10722;
    wire N__10721;
    wire N__10720;
    wire N__10719;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10704;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10681;
    wire N__10678;
    wire N__10677;
    wire N__10676;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10657;
    wire N__10656;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10493;
    wire N__10488;
    wire N__10485;
    wire N__10480;
    wire N__10479;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10472;
    wire N__10471;
    wire N__10468;
    wire N__10461;
    wire N__10456;
    wire N__10455;
    wire N__10454;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10436;
    wire N__10431;
    wire N__10426;
    wire N__10425;
    wire N__10422;
    wire N__10417;
    wire N__10414;
    wire N__10409;
    wire N__10398;
    wire N__10395;
    wire N__10394;
    wire N__10391;
    wire N__10386;
    wire N__10379;
    wire N__10376;
    wire N__10375;
    wire N__10374;
    wire N__10373;
    wire N__10366;
    wire N__10365;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10348;
    wire N__10347;
    wire N__10346;
    wire N__10341;
    wire N__10336;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10315;
    wire N__10310;
    wire N__10297;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10285;
    wire N__10282;
    wire N__10273;
    wire N__10266;
    wire N__10263;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10229;
    wire N__10228;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10220;
    wire N__10219;
    wire N__10218;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10213;
    wire N__10212;
    wire N__10211;
    wire N__10210;
    wire N__10209;
    wire N__10208;
    wire N__10207;
    wire N__10206;
    wire N__10205;
    wire N__10204;
    wire N__10203;
    wire N__10202;
    wire N__10201;
    wire N__10200;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10195;
    wire N__10194;
    wire N__10193;
    wire N__10192;
    wire N__10191;
    wire N__10188;
    wire N__10187;
    wire N__10186;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10038;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10010;
    wire N__10009;
    wire N__10008;
    wire N__10005;
    wire N__10000;
    wire N__9997;
    wire N__9996;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9948;
    wire N__9945;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9880;
    wire N__9875;
    wire N__9872;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9820;
    wire N__9815;
    wire N__9812;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9788;
    wire N__9787;
    wire N__9784;
    wire N__9779;
    wire N__9774;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9737;
    wire N__9734;
    wire N__9729;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9564;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9549;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9510;
    wire N__9507;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9486;
    wire N__9477;
    wire N__9474;
    wire N__9473;
    wire N__9472;
    wire N__9469;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9447;
    wire N__9446;
    wire N__9445;
    wire N__9444;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9396;
    wire N__9391;
    wire N__9386;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9338;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9301;
    wire N__9300;
    wire N__9295;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9254;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9188;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9168;
    wire N__9165;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9110;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9090;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8980;
    wire N__8975;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8960;
    wire N__8957;
    wire N__8946;
    wire N__8945;
    wire N__8942;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8932;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8913;
    wire N__8910;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8823;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8699;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8680;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8525;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8514;
    wire N__8513;
    wire N__8510;
    wire N__8505;
    wire N__8498;
    wire N__8493;
    wire N__8484;
    wire N__8483;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8460;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8427;
    wire N__8424;
    wire N__8419;
    wire N__8416;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8382;
    wire N__8381;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8375;
    wire N__8370;
    wire N__8369;
    wire N__8366;
    wire N__8365;
    wire N__8364;
    wire N__8361;
    wire N__8360;
    wire N__8359;
    wire N__8358;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8346;
    wire N__8343;
    wire N__8342;
    wire N__8341;
    wire N__8340;
    wire N__8339;
    wire N__8338;
    wire N__8337;
    wire N__8336;
    wire N__8335;
    wire N__8334;
    wire N__8333;
    wire N__8330;
    wire N__8325;
    wire N__8318;
    wire N__8311;
    wire N__8308;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8282;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8223;
    wire N__8220;
    wire N__8219;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8202;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8178;
    wire N__8169;
    wire N__8166;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8151;
    wire N__8150;
    wire N__8149;
    wire N__8142;
    wire N__8139;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8091;
    wire N__8088;
    wire N__8087;
    wire N__8086;
    wire N__8083;
    wire N__8078;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8003;
    wire N__8002;
    wire N__8001;
    wire N__8000;
    wire N__7999;
    wire N__7998;
    wire N__7995;
    wire N__7990;
    wire N__7989;
    wire N__7986;
    wire N__7985;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7974;
    wire N__7969;
    wire N__7968;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7963;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7957;
    wire N__7956;
    wire N__7955;
    wire N__7954;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7931;
    wire N__7926;
    wire N__7921;
    wire N__7910;
    wire N__7899;
    wire N__7892;
    wire N__7889;
    wire N__7884;
    wire N__7879;
    wire N__7874;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7790;
    wire N__7789;
    wire N__7786;
    wire N__7781;
    wire N__7776;
    wire N__7773;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7758;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7737;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7729;
    wire N__7724;
    wire N__7723;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7611;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7593;
    wire N__7592;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7527;
    wire N__7524;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7423;
    wire N__7418;
    wire N__7415;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7400;
    wire N__7399;
    wire N__7396;
    wire N__7391;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7376;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7362;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7350;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7326;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7304;
    wire N__7303;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7275;
    wire N__7274;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7260;
    wire N__7259;
    wire N__7256;
    wire N__7255;
    wire N__7254;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7246;
    wire N__7241;
    wire N__7238;
    wire N__7233;
    wire N__7226;
    wire N__7215;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7172;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7164;
    wire N__7163;
    wire N__7160;
    wire N__7159;
    wire N__7158;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7138;
    wire N__7135;
    wire N__7134;
    wire N__7131;
    wire N__7130;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7090;
    wire N__7087;
    wire N__7068;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7058;
    wire N__7055;
    wire N__7050;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7035;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7004;
    wire N__7001;
    wire N__6984;
    wire N__6983;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6958;
    wire N__6953;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6942;
    wire N__6939;
    wire N__6934;
    wire N__6931;
    wire N__6926;
    wire N__6923;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6902;
    wire N__6901;
    wire N__6898;
    wire N__6893;
    wire N__6888;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6873;
    wire N__6870;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6855;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6824;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6816;
    wire N__6813;
    wire N__6812;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6794;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6767;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6561;
    wire N__6560;
    wire N__6559;
    wire N__6558;
    wire N__6557;
    wire N__6556;
    wire N__6555;
    wire N__6554;
    wire N__6553;
    wire N__6552;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6548;
    wire N__6547;
    wire N__6544;
    wire N__6539;
    wire N__6532;
    wire N__6527;
    wire N__6520;
    wire N__6513;
    wire N__6510;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6480;
    wire N__6477;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6473;
    wire N__6472;
    wire N__6471;
    wire N__6468;
    wire N__6467;
    wire N__6466;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6456;
    wire N__6455;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6435;
    wire N__6432;
    wire N__6427;
    wire N__6422;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6349;
    wire N__6348;
    wire N__6347;
    wire N__6346;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6328;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6307;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6289;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6132;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6059;
    wire N__6058;
    wire N__6057;
    wire N__6054;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6033;
    wire N__6028;
    wire N__6023;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5858;
    wire N__5857;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5798;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5774;
    wire N__5771;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5715;
    wire N__5714;
    wire N__5713;
    wire N__5712;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5654;
    wire N__5651;
    wire N__5646;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5628;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5598;
    wire N__5595;
    wire N__5594;
    wire N__5593;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5546;
    wire N__5543;
    wire N__5542;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5532;
    wire N__5531;
    wire N__5528;
    wire N__5527;
    wire N__5526;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5507;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5485;
    wire N__5478;
    wire N__5475;
    wire N__5470;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5400;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5390;
    wire N__5389;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5360;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5298;
    wire N__5295;
    wire N__5294;
    wire N__5289;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5163;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5118;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5103;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4988;
    wire N__4987;
    wire N__4986;
    wire N__4983;
    wire N__4976;
    wire N__4969;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4685;
    wire N__4684;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4584;
    wire N__4581;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_iso_i;
    wire \INVU712_CYCLE_TERM.TACK_STATE_3C_net ;
    wire CLK40_PLL_i_i;
    wire \U712_CHIP_RAM.N_592_cascade_ ;
    wire \U712_CHIP_RAM.N_482_cascade_ ;
    wire bfn_7_12_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_483 ;
    wire \U712_CHIP_RAM.N_335_cascade_ ;
    wire \U712_CHIP_RAM.N_507_cascade_ ;
    wire \U712_CHIP_RAM.N_477 ;
    wire \U712_CHIP_RAM.N_477_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.N_406_cascade_ ;
    wire TACK_OUT;
    wire \INVU712_CYCLE_TERM.TACK_OUTC_net ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0 ;
    wire \U712_CHIP_RAM.N_478 ;
    wire A_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire VBENn_c;
    wire CMA_c_10;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.SDRAM_COUNTER19_cascade_ ;
    wire \U712_CHIP_RAM.N_349_cascade_ ;
    wire \U712_CHIP_RAM.N_349 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.N_509 ;
    wire \U712_CHIP_RAM.N_509_cascade_ ;
    wire \U712_CHIP_RAM.N_504 ;
    wire \U712_CHIP_RAM.N_583_cascade_ ;
    wire \U712_CHIP_RAM.N_591 ;
    wire \U712_CHIP_RAM.N_402_cascade_ ;
    wire \U712_CHIP_RAM.N_375_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0 ;
    wire \U712_CHIP_RAM.N_375_0_i_cascade_ ;
    wire \U712_CHIP_RAM.N_402 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_426 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_586 ;
    wire \U712_CHIP_RAM.N_359 ;
    wire \U712_CHIP_RAM.N_586_cascade_ ;
    wire \U712_CHIP_RAM.N_419_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_332_cascade_ ;
    wire \U712_CHIP_RAM.N_510_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire CMA_c_1;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.N_389 ;
    wire \U712_CHIP_RAM.N_343_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.N_334 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1 ;
    wire \U712_CHIP_RAM.N_366_cascade_ ;
    wire \U712_CHIP_RAM.N_335 ;
    wire \U712_CHIP_RAM.DBENn_8_1_cascade_ ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_ ;
    wire AWEn_c;
    wire DMA_LATCH_EN_c;
    wire DMA_WRITE_CYCLE;
    wire DRDDIR_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_503_cascade_ ;
    wire \U712_CHIP_RAM.N_420 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_590 ;
    wire \U712_CHIP_RAM.N_476 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_248_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_358_i_cascade_ ;
    wire TACK_EN;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \INVU712_CYCLE_TERM.TACK_STATE_1C_net ;
    wire DBRn_c;
    wire \U712_REG_SM.N_352_cascade_ ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire UDSn_c;
    wire \U712_REG_SM.N_429 ;
    wire LDSn_c;
    wire \U712_REG_SM.N_493 ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ;
    wire A_c_14;
    wire \U712_CHIP_RAM.N_383 ;
    wire CMA_c_3;
    wire CMA_c_4;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.N_343 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire A_c_2;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire A_c_4;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_7;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire A_c_8;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_514_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_350 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ;
    wire \U712_CHIP_RAM.N_501 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.N_481_cascade_ ;
    wire \U712_REG_SM.N_428_cascade_ ;
    wire REGSPACEn_c;
    wire \U712_CHIP_RAM.N_500 ;
    wire \U712_CHIP_RAM.N_503 ;
    wire \U712_CHIP_RAM.N_500_cascade_ ;
    wire \U712_CHIP_RAM.N_514 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.N_337 ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_332 ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.N_248_0 ;
    wire RnW_c;
    wire DBR_SYNCZ0Z_0;
    wire REG_TACK;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire C3_c;
    wire BLSn_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_345_cascade_ ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_396 ;
    wire \U712_REG_SM.N_435_cascade_ ;
    wire \U712_REG_SM.N_352 ;
    wire \U712_REG_SM.N_357 ;
    wire \U712_REG_SM.N_353 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire \U712_CHIP_RAM.N_450 ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_510 ;
    wire \U712_CHIP_RAM.N_461 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ;
    wire LATCH_CLK_c;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire PRnW_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_351_cascade_ ;
    wire \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire TSn_c;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.N_448_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.N_365 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_4 ;
    wire \U712_REG_SM.N_588 ;
    wire \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_8 ;
    wire \U712_REG_SM.N_395_cascade_ ;
    wire \U712_REG_SM.N_439_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_5_iv_0_0 ;
    wire \U712_REG_SM.N_395 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_131 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_7 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ;
    wire REG_CYCLEm;
    wire N_196_i;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.N_492 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire DBR_SYNC_i_1;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire bfn_12_13_0_;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire \U712_REG_SM.N_351 ;
    wire \U712_REG_SM.N_435 ;
    wire \U712_REG_SM.N_345 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_131_0 ;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_8;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire DRA_c_0;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_13_12_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_6;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DRA_c_3;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire N_412_i;
    wire AGNUS_REV_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RAS0n_c;
    wire RAS1n_c;
    wire RESETn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire CLK80_PLL;
    wire \U712_BYTE_ENABLE.N_467 ;
    wire \U712_BYTE_ENABLE.N_455_cascade_ ;
    wire N_38_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_455 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_ ;
    wire N_209_i;
    wire \U712_BYTE_ENABLE.N_331_i ;
    wire CPU_CYCLEm;
    wire N_205;
    wire N_411_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire N_213;
    wire \U712_BYTE_ENABLE.N_464 ;
    wire N_40_i;
    wire \U712_BYTE_ENABLE.N_452 ;
    wire CASUn_c;
    wire N_208_i;
    wire CASLn_c;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_BYTE_ENABLE.N_456 ;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4521),
            .RESETB(N__8409),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12850),
            .DIN(N__12849),
            .DOUT(N__12848),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12850),
            .PADOUT(N__12849),
            .PADIN(N__12848),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11202),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12841),
            .DIN(N__12840),
            .DOUT(N__12839),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12841),
            .PADOUT(N__12840),
            .PADIN(N__12839),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12832),
            .DIN(N__12831),
            .DOUT(N__12830),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12832),
            .PADOUT(N__12831),
            .PADIN(N__12830),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7635),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12823),
            .DIN(N__12822),
            .DOUT(N__12821),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12823),
            .PADOUT(N__12822),
            .PADIN(N__12821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12814),
            .DIN(N__12813),
            .DOUT(N__12812),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12814),
            .PADOUT(N__12813),
            .PADIN(N__12812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12805),
            .DIN(N__12804),
            .DOUT(N__12803),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12805),
            .PADOUT(N__12804),
            .PADIN(N__12803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12796),
            .DIN(N__12795),
            .DOUT(N__12794),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12796),
            .PADOUT(N__12795),
            .PADIN(N__12794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12787),
            .DIN(N__12786),
            .DOUT(N__12785),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12787),
            .PADOUT(N__12786),
            .PADIN(N__12785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12778),
            .DIN(N__12777),
            .DOUT(N__12776),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12778),
            .PADOUT(N__12777),
            .PADIN(N__12776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12769),
            .DIN(N__12768),
            .DOUT(N__12767),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12769),
            .PADOUT(N__12768),
            .PADIN(N__12767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12760),
            .DIN(N__12759),
            .DOUT(N__12758),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12760),
            .PADOUT(N__12759),
            .PADIN(N__12758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12751),
            .DIN(N__12750),
            .DOUT(N__12749),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12751),
            .PADOUT(N__12750),
            .PADIN(N__12749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6084),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12742),
            .DIN(N__12741),
            .DOUT(N__12740),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12742),
            .PADOUT(N__12741),
            .PADIN(N__12740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11058),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12733),
            .DIN(N__12732),
            .DOUT(N__12731),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12733),
            .PADOUT(N__12732),
            .PADIN(N__12731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12724),
            .DIN(N__12723),
            .DOUT(N__12722),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12724),
            .PADOUT(N__12723),
            .PADIN(N__12722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8114),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12715),
            .DIN(N__12714),
            .DOUT(N__12713),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12715),
            .PADOUT(N__12714),
            .PADIN(N__12713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12706),
            .DIN(N__12705),
            .DOUT(N__12704),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12706),
            .PADOUT(N__12705),
            .PADIN(N__12704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12697),
            .DIN(N__12696),
            .DOUT(N__12695),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12697),
            .PADOUT(N__12696),
            .PADIN(N__12695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12688),
            .DIN(N__12687),
            .DOUT(N__12686),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12688),
            .PADOUT(N__12687),
            .PADIN(N__12686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12679),
            .DIN(N__12678),
            .DOUT(N__12677),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12679),
            .PADOUT(N__12678),
            .PADIN(N__12677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12670),
            .DIN(N__12669),
            .DOUT(N__12668),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12670),
            .PADOUT(N__12669),
            .PADIN(N__12668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5079),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12661),
            .DIN(N__12660),
            .DOUT(N__12659),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12661),
            .PADOUT(N__12660),
            .PADIN(N__12659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12652),
            .DIN(N__12651),
            .DOUT(N__12650),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12652),
            .PADOUT(N__12651),
            .PADIN(N__12650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12643),
            .DIN(N__12642),
            .DOUT(N__12641),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12643),
            .PADOUT(N__12642),
            .PADIN(N__12641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12634),
            .DIN(N__12633),
            .DOUT(N__12632),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12634),
            .PADOUT(N__12633),
            .PADIN(N__12632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12625),
            .DIN(N__12624),
            .DOUT(N__12623),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12625),
            .PADOUT(N__12624),
            .PADIN(N__12623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5775),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12616),
            .DIN(N__12615),
            .DOUT(N__12614),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12616),
            .PADOUT(N__12615),
            .PADIN(N__12614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12607),
            .DIN(N__12606),
            .DOUT(N__12605),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12607),
            .PADOUT(N__12606),
            .PADIN(N__12605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12598),
            .DIN(N__12597),
            .DOUT(N__12596),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12598),
            .PADOUT(N__12597),
            .PADIN(N__12596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12589),
            .DIN(N__12588),
            .DOUT(N__12587),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12589),
            .PADOUT(N__12588),
            .PADIN(N__12587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12580),
            .DIN(N__12579),
            .DOUT(N__12578),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12580),
            .PADOUT(N__12579),
            .PADIN(N__12578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12571),
            .DIN(N__12570),
            .DOUT(N__12569),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12571),
            .PADOUT(N__12570),
            .PADIN(N__12569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5265),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12562),
            .DIN(N__12561),
            .DOUT(N__12560),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12562),
            .PADOUT(N__12561),
            .PADIN(N__12560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12553),
            .DIN(N__12552),
            .DOUT(N__12551),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12553),
            .PADOUT(N__12552),
            .PADIN(N__12551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12544),
            .DIN(N__12543),
            .DOUT(N__12542),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12544),
            .PADOUT(N__12543),
            .PADIN(N__12542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12535),
            .DIN(N__12534),
            .DOUT(N__12533),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12535),
            .PADOUT(N__12534),
            .PADIN(N__12533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12526),
            .DIN(N__12525),
            .DOUT(N__12524),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12526),
            .PADOUT(N__12525),
            .PADIN(N__12524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12517),
            .DIN(N__12516),
            .DOUT(N__12515),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12517),
            .PADOUT(N__12516),
            .PADIN(N__12515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7572),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12508),
            .DIN(N__12507),
            .DOUT(N__12506),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12508),
            .PADOUT(N__12507),
            .PADIN(N__12506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12499),
            .DIN(N__12498),
            .DOUT(N__12497),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12499),
            .PADOUT(N__12498),
            .PADIN(N__12497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12490),
            .DIN(N__12489),
            .DOUT(N__12488),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12490),
            .PADOUT(N__12489),
            .PADIN(N__12488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9375),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12481),
            .DIN(N__12480),
            .DOUT(N__12479),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12481),
            .PADOUT(N__12480),
            .PADIN(N__12479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4833),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12472),
            .DIN(N__12471),
            .DOUT(N__12470),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12472),
            .PADOUT(N__12471),
            .PADIN(N__12470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12463),
            .DIN(N__12462),
            .DOUT(N__12461),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12463),
            .PADOUT(N__12462),
            .PADIN(N__12461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12454),
            .DIN(N__12453),
            .DOUT(N__12452),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12454),
            .PADOUT(N__12453),
            .PADIN(N__12452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6132),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12445),
            .DIN(N__12444),
            .DOUT(N__12443),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12445),
            .PADOUT(N__12444),
            .PADIN(N__12443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12436),
            .DIN(N__12435),
            .DOUT(N__12434),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12436),
            .PADOUT(N__12435),
            .PADIN(N__12434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11382),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12427),
            .DIN(N__12426),
            .DOUT(N__12425),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12427),
            .PADOUT(N__12426),
            .PADIN(N__12425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9978),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12418),
            .DIN(N__12417),
            .DOUT(N__12416),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12418),
            .PADOUT(N__12417),
            .PADIN(N__12416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5325),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12409),
            .DIN(N__12408),
            .DOUT(N__12407),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12409),
            .PADOUT(N__12408),
            .PADIN(N__12407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11943),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12400),
            .DIN(N__12399),
            .DOUT(N__12398),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12400),
            .PADOUT(N__12399),
            .PADIN(N__12398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12391),
            .DIN(N__12390),
            .DOUT(N__12389),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12391),
            .PADOUT(N__12390),
            .PADIN(N__12389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12382),
            .DIN(N__12381),
            .DOUT(N__12380),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12382),
            .PADOUT(N__12381),
            .PADIN(N__12380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4770),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12373),
            .DIN(N__12372),
            .DOUT(N__12371),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12373),
            .PADOUT(N__12372),
            .PADIN(N__12371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12364),
            .DIN(N__12363),
            .DOUT(N__12362),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12364),
            .PADOUT(N__12363),
            .PADIN(N__12362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12355),
            .DIN(N__12354),
            .DOUT(N__12353),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12355),
            .PADOUT(N__12354),
            .PADIN(N__12353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5058),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12346),
            .DIN(N__12345),
            .DOUT(N__12344),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12346),
            .PADOUT(N__12345),
            .PADIN(N__12344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11739),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12337),
            .DIN(N__12336),
            .DOUT(N__12335),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12337),
            .PADOUT(N__12336),
            .PADIN(N__12335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12328),
            .DIN(N__12327),
            .DOUT(N__12326),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12328),
            .PADOUT(N__12327),
            .PADIN(N__12326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11298),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12319),
            .DIN(N__12318),
            .DOUT(N__12317),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12319),
            .PADOUT(N__12318),
            .PADIN(N__12317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5770),
            .DIN0(),
            .DOUT0(N__4665),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12310),
            .DIN(N__12309),
            .DOUT(N__12308),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12310),
            .PADOUT(N__12309),
            .PADIN(N__12308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12301),
            .DIN(N__12300),
            .DOUT(N__12299),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12301),
            .PADOUT(N__12300),
            .PADIN(N__12299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12292),
            .DIN(N__12291),
            .DOUT(N__12290),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12292),
            .PADOUT(N__12291),
            .PADIN(N__12290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12283),
            .DIN(N__12282),
            .DOUT(N__12281),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12283),
            .PADOUT(N__12282),
            .PADIN(N__12281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5991),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12274),
            .DIN(N__12273),
            .DOUT(N__12272),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12274),
            .PADOUT(N__12273),
            .PADIN(N__12272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12265),
            .DIN(N__12264),
            .DOUT(N__12263),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12265),
            .PADOUT(N__12264),
            .PADIN(N__12263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12256),
            .DIN(N__12255),
            .DOUT(N__12254),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12256),
            .PADOUT(N__12255),
            .PADIN(N__12254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12247),
            .DIN(N__12246),
            .DOUT(N__12245),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12247),
            .PADOUT(N__12246),
            .PADIN(N__12245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12238),
            .DIN(N__12237),
            .DOUT(N__12236),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12238),
            .PADOUT(N__12237),
            .PADIN(N__12236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12229),
            .DIN(N__12228),
            .DOUT(N__12227),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12229),
            .PADOUT(N__12228),
            .PADIN(N__12227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5040),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12220),
            .DIN(N__12219),
            .DOUT(N__12218),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12220),
            .PADOUT(N__12219),
            .PADIN(N__12218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5928),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12211),
            .DIN(N__12210),
            .DOUT(N__12209),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12211),
            .PADOUT(N__12210),
            .PADIN(N__12209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12202),
            .DIN(N__12201),
            .DOUT(N__12200),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12202),
            .PADOUT(N__12201),
            .PADIN(N__12200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4929),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12193),
            .DIN(N__12192),
            .DOUT(N__12191),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12193),
            .PADOUT(N__12192),
            .PADIN(N__12191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12184),
            .DIN(N__12183),
            .DOUT(N__12182),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12184),
            .PADOUT(N__12183),
            .PADIN(N__12182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12175),
            .DIN(N__12174),
            .DOUT(N__12173),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12175),
            .PADOUT(N__12174),
            .PADIN(N__12173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6117),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12166),
            .DIN(N__12165),
            .DOUT(N__12164),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12166),
            .PADOUT(N__12165),
            .PADIN(N__12164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12157),
            .DIN(N__12156),
            .DOUT(N__12155),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12157),
            .PADOUT(N__12156),
            .PADIN(N__12155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12148),
            .DIN(N__12147),
            .DOUT(N__12146),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12148),
            .PADOUT(N__12147),
            .PADIN(N__12146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7680),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12139),
            .DIN(N__12138),
            .DOUT(N__12137),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12139),
            .PADOUT(N__12138),
            .PADIN(N__12137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5895),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12130),
            .DIN(N__12129),
            .DOUT(N__12128),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12130),
            .PADOUT(N__12129),
            .PADIN(N__12128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4602),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PRnW_obuf_iopad (
            .OE(N__12121),
            .DIN(N__12120),
            .DOUT(N__12119),
            .PACKAGEPIN(PRnW));
    defparam PRnW_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PRnW_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PRnW_obuf_preio (
            .PADOEN(N__12121),
            .PADOUT(N__12120),
            .PADIN(N__12119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8250),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12112),
            .DIN(N__12111),
            .DOUT(N__12110),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12112),
            .PADOUT(N__12111),
            .PADIN(N__12110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12103),
            .DIN(N__12102),
            .DOUT(N__12101),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12103),
            .PADOUT(N__12102),
            .PADIN(N__12101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4601),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12094),
            .DIN(N__12093),
            .DOUT(N__12092),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12094),
            .PADOUT(N__12093),
            .PADIN(N__12092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4539),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12085),
            .DIN(N__12084),
            .DOUT(N__12083),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12085),
            .PADOUT(N__12084),
            .PADIN(N__12083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12076),
            .DIN(N__12075),
            .DOUT(N__12074),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12076),
            .PADOUT(N__12075),
            .PADIN(N__12074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12067),
            .DIN(N__12066),
            .DOUT(N__12065),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12067),
            .PADOUT(N__12066),
            .PADIN(N__12065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12058),
            .DIN(N__12057),
            .DOUT(N__12056),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12058),
            .PADOUT(N__12057),
            .PADIN(N__12056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BLSn_obuf_iopad (
            .OE(N__12049),
            .DIN(N__12048),
            .DOUT(N__12047),
            .PACKAGEPIN(BLSn));
    defparam BLSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BLSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BLSn_obuf_preio (
            .PADOEN(N__12049),
            .PADOUT(N__12048),
            .PADIN(N__12047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7458),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12040),
            .DIN(N__12039),
            .DOUT(N__12038),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12040),
            .PADOUT(N__12039),
            .PADIN(N__12038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12031),
            .DIN(N__12030),
            .DOUT(N__12029),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12031),
            .PADOUT(N__12030),
            .PADIN(N__12029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4580),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12022),
            .DIN(N__12021),
            .DOUT(N__12020),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12022),
            .PADOUT(N__12021),
            .PADIN(N__12020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8805),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12013),
            .DIN(N__12012),
            .DOUT(N__12011),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12013),
            .PADOUT(N__12012),
            .PADIN(N__12011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10083),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12004),
            .DIN(N__12003),
            .DOUT(N__12002),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12004),
            .PADOUT(N__12003),
            .PADIN(N__12002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6378),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11995),
            .DIN(N__11994),
            .DOUT(N__11993),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11995),
            .PADOUT(N__11994),
            .PADIN(N__11993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11986),
            .DIN(N__11985),
            .DOUT(N__11984),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11986),
            .PADOUT(N__11985),
            .PADIN(N__11984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11977),
            .DIN(N__11976),
            .DOUT(N__11975),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11977),
            .PADOUT(N__11976),
            .PADIN(N__11975),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5774),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2876 (
            .O(N__11958),
            .I(N__11955));
    LocalMux I__2875 (
            .O(N__11955),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ));
    InMux I__2874 (
            .O(N__11952),
            .I(N__11949));
    LocalMux I__2873 (
            .O(N__11949),
            .I(\U712_BYTE_ENABLE.N_455 ));
    CascadeMux I__2872 (
            .O(N__11946),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_ ));
    IoInMux I__2871 (
            .O(N__11943),
            .I(N__11940));
    LocalMux I__2870 (
            .O(N__11940),
            .I(N__11937));
    Span4Mux_s1_h I__2869 (
            .O(N__11937),
            .I(N__11934));
    Sp12to4 I__2868 (
            .O(N__11934),
            .I(N__11931));
    Span12Mux_s11_v I__2867 (
            .O(N__11931),
            .I(N__11928));
    Span12Mux_h I__2866 (
            .O(N__11928),
            .I(N__11925));
    Odrv12 I__2865 (
            .O(N__11925),
            .I(N_209_i));
    CascadeMux I__2864 (
            .O(N__11922),
            .I(N__11918));
    InMux I__2863 (
            .O(N__11921),
            .I(N__11915));
    InMux I__2862 (
            .O(N__11918),
            .I(N__11912));
    LocalMux I__2861 (
            .O(N__11915),
            .I(\U712_BYTE_ENABLE.N_331_i ));
    LocalMux I__2860 (
            .O(N__11912),
            .I(\U712_BYTE_ENABLE.N_331_i ));
    InMux I__2859 (
            .O(N__11907),
            .I(N__11894));
    InMux I__2858 (
            .O(N__11906),
            .I(N__11894));
    InMux I__2857 (
            .O(N__11905),
            .I(N__11894));
    CascadeMux I__2856 (
            .O(N__11904),
            .I(N__11890));
    CascadeMux I__2855 (
            .O(N__11903),
            .I(N__11887));
    InMux I__2854 (
            .O(N__11902),
            .I(N__11883));
    InMux I__2853 (
            .O(N__11901),
            .I(N__11880));
    LocalMux I__2852 (
            .O(N__11894),
            .I(N__11877));
    InMux I__2851 (
            .O(N__11893),
            .I(N__11865));
    InMux I__2850 (
            .O(N__11890),
            .I(N__11860));
    InMux I__2849 (
            .O(N__11887),
            .I(N__11856));
    InMux I__2848 (
            .O(N__11886),
            .I(N__11853));
    LocalMux I__2847 (
            .O(N__11883),
            .I(N__11848));
    LocalMux I__2846 (
            .O(N__11880),
            .I(N__11848));
    Span4Mux_h I__2845 (
            .O(N__11877),
            .I(N__11845));
    InMux I__2844 (
            .O(N__11876),
            .I(N__11840));
    InMux I__2843 (
            .O(N__11875),
            .I(N__11840));
    InMux I__2842 (
            .O(N__11874),
            .I(N__11832));
    InMux I__2841 (
            .O(N__11873),
            .I(N__11832));
    InMux I__2840 (
            .O(N__11872),
            .I(N__11832));
    InMux I__2839 (
            .O(N__11871),
            .I(N__11825));
    InMux I__2838 (
            .O(N__11870),
            .I(N__11825));
    InMux I__2837 (
            .O(N__11869),
            .I(N__11825));
    InMux I__2836 (
            .O(N__11868),
            .I(N__11822));
    LocalMux I__2835 (
            .O(N__11865),
            .I(N__11819));
    InMux I__2834 (
            .O(N__11864),
            .I(N__11814));
    InMux I__2833 (
            .O(N__11863),
            .I(N__11814));
    LocalMux I__2832 (
            .O(N__11860),
            .I(N__11810));
    InMux I__2831 (
            .O(N__11859),
            .I(N__11807));
    LocalMux I__2830 (
            .O(N__11856),
            .I(N__11804));
    LocalMux I__2829 (
            .O(N__11853),
            .I(N__11799));
    Span4Mux_v I__2828 (
            .O(N__11848),
            .I(N__11799));
    Span4Mux_h I__2827 (
            .O(N__11845),
            .I(N__11794));
    LocalMux I__2826 (
            .O(N__11840),
            .I(N__11794));
    InMux I__2825 (
            .O(N__11839),
            .I(N__11791));
    LocalMux I__2824 (
            .O(N__11832),
            .I(N__11788));
    LocalMux I__2823 (
            .O(N__11825),
            .I(N__11779));
    LocalMux I__2822 (
            .O(N__11822),
            .I(N__11779));
    Span4Mux_h I__2821 (
            .O(N__11819),
            .I(N__11779));
    LocalMux I__2820 (
            .O(N__11814),
            .I(N__11779));
    InMux I__2819 (
            .O(N__11813),
            .I(N__11776));
    Odrv12 I__2818 (
            .O(N__11810),
            .I(CPU_CYCLEm));
    LocalMux I__2817 (
            .O(N__11807),
            .I(CPU_CYCLEm));
    Odrv4 I__2816 (
            .O(N__11804),
            .I(CPU_CYCLEm));
    Odrv4 I__2815 (
            .O(N__11799),
            .I(CPU_CYCLEm));
    Odrv4 I__2814 (
            .O(N__11794),
            .I(CPU_CYCLEm));
    LocalMux I__2813 (
            .O(N__11791),
            .I(CPU_CYCLEm));
    Odrv12 I__2812 (
            .O(N__11788),
            .I(CPU_CYCLEm));
    Odrv4 I__2811 (
            .O(N__11779),
            .I(CPU_CYCLEm));
    LocalMux I__2810 (
            .O(N__11776),
            .I(CPU_CYCLEm));
    IoInMux I__2809 (
            .O(N__11757),
            .I(N__11754));
    LocalMux I__2808 (
            .O(N__11754),
            .I(N__11751));
    IoSpan4Mux I__2807 (
            .O(N__11751),
            .I(N__11748));
    Span4Mux_s3_v I__2806 (
            .O(N__11748),
            .I(N__11745));
    Span4Mux_v I__2805 (
            .O(N__11745),
            .I(N__11742));
    Odrv4 I__2804 (
            .O(N__11742),
            .I(N_205));
    IoInMux I__2803 (
            .O(N__11739),
            .I(N__11736));
    LocalMux I__2802 (
            .O(N__11736),
            .I(N__11733));
    Span4Mux_s3_v I__2801 (
            .O(N__11733),
            .I(N__11730));
    Odrv4 I__2800 (
            .O(N__11730),
            .I(N_411_i));
    InMux I__2799 (
            .O(N__11727),
            .I(N__11721));
    InMux I__2798 (
            .O(N__11726),
            .I(N__11714));
    InMux I__2797 (
            .O(N__11725),
            .I(N__11714));
    InMux I__2796 (
            .O(N__11724),
            .I(N__11714));
    LocalMux I__2795 (
            .O(N__11721),
            .I(N__11706));
    LocalMux I__2794 (
            .O(N__11714),
            .I(N__11706));
    InMux I__2793 (
            .O(N__11713),
            .I(N__11701));
    InMux I__2792 (
            .O(N__11712),
            .I(N__11701));
    InMux I__2791 (
            .O(N__11711),
            .I(N__11698));
    Span4Mux_v I__2790 (
            .O(N__11706),
            .I(N__11695));
    LocalMux I__2789 (
            .O(N__11701),
            .I(N__11690));
    LocalMux I__2788 (
            .O(N__11698),
            .I(N__11690));
    Span4Mux_v I__2787 (
            .O(N__11695),
            .I(N__11684));
    Span4Mux_v I__2786 (
            .O(N__11690),
            .I(N__11684));
    InMux I__2785 (
            .O(N__11689),
            .I(N__11681));
    Sp12to4 I__2784 (
            .O(N__11684),
            .I(N__11676));
    LocalMux I__2783 (
            .O(N__11681),
            .I(N__11676));
    Span12Mux_h I__2782 (
            .O(N__11676),
            .I(N__11673));
    Odrv12 I__2781 (
            .O(N__11673),
            .I(A_c_1));
    InMux I__2780 (
            .O(N__11670),
            .I(N__11666));
    InMux I__2779 (
            .O(N__11669),
            .I(N__11658));
    LocalMux I__2778 (
            .O(N__11666),
            .I(N__11655));
    InMux I__2777 (
            .O(N__11665),
            .I(N__11650));
    InMux I__2776 (
            .O(N__11664),
            .I(N__11650));
    InMux I__2775 (
            .O(N__11663),
            .I(N__11645));
    InMux I__2774 (
            .O(N__11662),
            .I(N__11645));
    InMux I__2773 (
            .O(N__11661),
            .I(N__11642));
    LocalMux I__2772 (
            .O(N__11658),
            .I(N__11639));
    Span4Mux_h I__2771 (
            .O(N__11655),
            .I(N__11633));
    LocalMux I__2770 (
            .O(N__11650),
            .I(N__11633));
    LocalMux I__2769 (
            .O(N__11645),
            .I(N__11628));
    LocalMux I__2768 (
            .O(N__11642),
            .I(N__11628));
    Span4Mux_h I__2767 (
            .O(N__11639),
            .I(N__11625));
    InMux I__2766 (
            .O(N__11638),
            .I(N__11622));
    Span4Mux_v I__2765 (
            .O(N__11633),
            .I(N__11616));
    Span4Mux_v I__2764 (
            .O(N__11628),
            .I(N__11616));
    Span4Mux_h I__2763 (
            .O(N__11625),
            .I(N__11611));
    LocalMux I__2762 (
            .O(N__11622),
            .I(N__11611));
    InMux I__2761 (
            .O(N__11621),
            .I(N__11608));
    Sp12to4 I__2760 (
            .O(N__11616),
            .I(N__11605));
    Span4Mux_v I__2759 (
            .O(N__11611),
            .I(N__11602));
    LocalMux I__2758 (
            .O(N__11608),
            .I(N__11599));
    Span12Mux_h I__2757 (
            .O(N__11605),
            .I(N__11592));
    Sp12to4 I__2756 (
            .O(N__11602),
            .I(N__11592));
    Span12Mux_s10_v I__2755 (
            .O(N__11599),
            .I(N__11592));
    Odrv12 I__2754 (
            .O(N__11592),
            .I(A_c_0));
    CascadeMux I__2753 (
            .O(N__11589),
            .I(N__11584));
    CascadeMux I__2752 (
            .O(N__11588),
            .I(N__11579));
    CascadeMux I__2751 (
            .O(N__11587),
            .I(N__11576));
    InMux I__2750 (
            .O(N__11584),
            .I(N__11570));
    InMux I__2749 (
            .O(N__11583),
            .I(N__11570));
    CascadeMux I__2748 (
            .O(N__11582),
            .I(N__11567));
    InMux I__2747 (
            .O(N__11579),
            .I(N__11562));
    InMux I__2746 (
            .O(N__11576),
            .I(N__11562));
    CascadeMux I__2745 (
            .O(N__11575),
            .I(N__11559));
    LocalMux I__2744 (
            .O(N__11570),
            .I(N__11555));
    InMux I__2743 (
            .O(N__11567),
            .I(N__11552));
    LocalMux I__2742 (
            .O(N__11562),
            .I(N__11548));
    InMux I__2741 (
            .O(N__11559),
            .I(N__11545));
    InMux I__2740 (
            .O(N__11558),
            .I(N__11542));
    Span4Mux_v I__2739 (
            .O(N__11555),
            .I(N__11537));
    LocalMux I__2738 (
            .O(N__11552),
            .I(N__11537));
    CascadeMux I__2737 (
            .O(N__11551),
            .I(N__11533));
    Span4Mux_h I__2736 (
            .O(N__11548),
            .I(N__11530));
    LocalMux I__2735 (
            .O(N__11545),
            .I(N__11525));
    LocalMux I__2734 (
            .O(N__11542),
            .I(N__11525));
    Span4Mux_v I__2733 (
            .O(N__11537),
            .I(N__11522));
    InMux I__2732 (
            .O(N__11536),
            .I(N__11519));
    InMux I__2731 (
            .O(N__11533),
            .I(N__11516));
    Span4Mux_h I__2730 (
            .O(N__11530),
            .I(N__11511));
    Span4Mux_v I__2729 (
            .O(N__11525),
            .I(N__11511));
    Span4Mux_v I__2728 (
            .O(N__11522),
            .I(N__11508));
    LocalMux I__2727 (
            .O(N__11519),
            .I(N__11503));
    LocalMux I__2726 (
            .O(N__11516),
            .I(N__11503));
    Span4Mux_v I__2725 (
            .O(N__11511),
            .I(N__11500));
    Sp12to4 I__2724 (
            .O(N__11508),
            .I(N__11495));
    Span12Mux_v I__2723 (
            .O(N__11503),
            .I(N__11495));
    Sp12to4 I__2722 (
            .O(N__11500),
            .I(N__11492));
    Span12Mux_h I__2721 (
            .O(N__11495),
            .I(N__11489));
    Span12Mux_h I__2720 (
            .O(N__11492),
            .I(N__11486));
    Odrv12 I__2719 (
            .O(N__11489),
            .I(SIZ_c_1));
    Odrv12 I__2718 (
            .O(N__11486),
            .I(SIZ_c_1));
    InMux I__2717 (
            .O(N__11481),
            .I(N__11477));
    InMux I__2716 (
            .O(N__11480),
            .I(N__11474));
    LocalMux I__2715 (
            .O(N__11477),
            .I(N__11465));
    LocalMux I__2714 (
            .O(N__11474),
            .I(N__11465));
    InMux I__2713 (
            .O(N__11473),
            .I(N__11462));
    InMux I__2712 (
            .O(N__11472),
            .I(N__11457));
    InMux I__2711 (
            .O(N__11471),
            .I(N__11457));
    InMux I__2710 (
            .O(N__11470),
            .I(N__11454));
    Span4Mux_v I__2709 (
            .O(N__11465),
            .I(N__11448));
    LocalMux I__2708 (
            .O(N__11462),
            .I(N__11448));
    LocalMux I__2707 (
            .O(N__11457),
            .I(N__11443));
    LocalMux I__2706 (
            .O(N__11454),
            .I(N__11443));
    InMux I__2705 (
            .O(N__11453),
            .I(N__11440));
    Span4Mux_v I__2704 (
            .O(N__11448),
            .I(N__11437));
    Span4Mux_h I__2703 (
            .O(N__11443),
            .I(N__11434));
    LocalMux I__2702 (
            .O(N__11440),
            .I(N__11431));
    Span4Mux_v I__2701 (
            .O(N__11437),
            .I(N__11427));
    Span4Mux_h I__2700 (
            .O(N__11434),
            .I(N__11422));
    Span4Mux_v I__2699 (
            .O(N__11431),
            .I(N__11422));
    InMux I__2698 (
            .O(N__11430),
            .I(N__11419));
    Sp12to4 I__2697 (
            .O(N__11427),
            .I(N__11416));
    Span4Mux_v I__2696 (
            .O(N__11422),
            .I(N__11413));
    LocalMux I__2695 (
            .O(N__11419),
            .I(N__11410));
    Span12Mux_h I__2694 (
            .O(N__11416),
            .I(N__11403));
    Sp12to4 I__2693 (
            .O(N__11413),
            .I(N__11403));
    Span12Mux_v I__2692 (
            .O(N__11410),
            .I(N__11403));
    Odrv12 I__2691 (
            .O(N__11403),
            .I(SIZ_c_0));
    IoInMux I__2690 (
            .O(N__11400),
            .I(N__11397));
    LocalMux I__2689 (
            .O(N__11397),
            .I(N__11394));
    Span4Mux_s3_v I__2688 (
            .O(N__11394),
            .I(N__11391));
    Odrv4 I__2687 (
            .O(N__11391),
            .I(N_213));
    InMux I__2686 (
            .O(N__11388),
            .I(N__11385));
    LocalMux I__2685 (
            .O(N__11385),
            .I(\U712_BYTE_ENABLE.N_464 ));
    IoInMux I__2684 (
            .O(N__11382),
            .I(N__11379));
    LocalMux I__2683 (
            .O(N__11379),
            .I(N__11376));
    Sp12to4 I__2682 (
            .O(N__11376),
            .I(N__11373));
    Span12Mux_h I__2681 (
            .O(N__11373),
            .I(N__11370));
    Span12Mux_v I__2680 (
            .O(N__11370),
            .I(N__11367));
    Odrv12 I__2679 (
            .O(N__11367),
            .I(N_40_i));
    InMux I__2678 (
            .O(N__11364),
            .I(N__11361));
    LocalMux I__2677 (
            .O(N__11361),
            .I(\U712_BYTE_ENABLE.N_452 ));
    InMux I__2676 (
            .O(N__11358),
            .I(N__11352));
    InMux I__2675 (
            .O(N__11357),
            .I(N__11352));
    LocalMux I__2674 (
            .O(N__11352),
            .I(N__11346));
    InMux I__2673 (
            .O(N__11351),
            .I(N__11343));
    InMux I__2672 (
            .O(N__11350),
            .I(N__11340));
    CascadeMux I__2671 (
            .O(N__11349),
            .I(N__11336));
    Span4Mux_v I__2670 (
            .O(N__11346),
            .I(N__11333));
    LocalMux I__2669 (
            .O(N__11343),
            .I(N__11328));
    LocalMux I__2668 (
            .O(N__11340),
            .I(N__11328));
    InMux I__2667 (
            .O(N__11339),
            .I(N__11323));
    InMux I__2666 (
            .O(N__11336),
            .I(N__11323));
    Span4Mux_h I__2665 (
            .O(N__11333),
            .I(N__11318));
    Span4Mux_v I__2664 (
            .O(N__11328),
            .I(N__11318));
    LocalMux I__2663 (
            .O(N__11323),
            .I(N__11315));
    Span4Mux_h I__2662 (
            .O(N__11318),
            .I(N__11310));
    Span4Mux_v I__2661 (
            .O(N__11315),
            .I(N__11310));
    Sp12to4 I__2660 (
            .O(N__11310),
            .I(N__11307));
    Span12Mux_h I__2659 (
            .O(N__11307),
            .I(N__11304));
    Span12Mux_v I__2658 (
            .O(N__11304),
            .I(N__11301));
    Odrv12 I__2657 (
            .O(N__11301),
            .I(CASUn_c));
    IoInMux I__2656 (
            .O(N__11298),
            .I(N__11295));
    LocalMux I__2655 (
            .O(N__11295),
            .I(N__11292));
    Span4Mux_s3_h I__2654 (
            .O(N__11292),
            .I(N__11289));
    Span4Mux_v I__2653 (
            .O(N__11289),
            .I(N__11286));
    Span4Mux_h I__2652 (
            .O(N__11286),
            .I(N__11283));
    Span4Mux_h I__2651 (
            .O(N__11283),
            .I(N__11280));
    Odrv4 I__2650 (
            .O(N__11280),
            .I(N_208_i));
    InMux I__2649 (
            .O(N__11277),
            .I(N__11273));
    CascadeMux I__2648 (
            .O(N__11276),
            .I(N__11269));
    LocalMux I__2647 (
            .O(N__11273),
            .I(N__11264));
    InMux I__2646 (
            .O(N__11272),
            .I(N__11261));
    InMux I__2645 (
            .O(N__11269),
            .I(N__11255));
    InMux I__2644 (
            .O(N__11268),
            .I(N__11255));
    InMux I__2643 (
            .O(N__11267),
            .I(N__11252));
    Span4Mux_h I__2642 (
            .O(N__11264),
            .I(N__11247));
    LocalMux I__2641 (
            .O(N__11261),
            .I(N__11247));
    InMux I__2640 (
            .O(N__11260),
            .I(N__11244));
    LocalMux I__2639 (
            .O(N__11255),
            .I(N__11241));
    LocalMux I__2638 (
            .O(N__11252),
            .I(N__11238));
    Sp12to4 I__2637 (
            .O(N__11247),
            .I(N__11235));
    LocalMux I__2636 (
            .O(N__11244),
            .I(N__11232));
    Span12Mux_h I__2635 (
            .O(N__11241),
            .I(N__11229));
    Span12Mux_v I__2634 (
            .O(N__11238),
            .I(N__11226));
    Span12Mux_h I__2633 (
            .O(N__11235),
            .I(N__11223));
    Span12Mux_v I__2632 (
            .O(N__11232),
            .I(N__11220));
    Span12Mux_v I__2631 (
            .O(N__11229),
            .I(N__11217));
    Span12Mux_h I__2630 (
            .O(N__11226),
            .I(N__11214));
    Span12Mux_v I__2629 (
            .O(N__11223),
            .I(N__11209));
    Span12Mux_h I__2628 (
            .O(N__11220),
            .I(N__11209));
    Odrv12 I__2627 (
            .O(N__11217),
            .I(CASLn_c));
    Odrv12 I__2626 (
            .O(N__11214),
            .I(CASLn_c));
    Odrv12 I__2625 (
            .O(N__11209),
            .I(CASLn_c));
    IoInMux I__2624 (
            .O(N__11202),
            .I(N__11199));
    LocalMux I__2623 (
            .O(N__11199),
            .I(N__11195));
    CascadeMux I__2622 (
            .O(N__11198),
            .I(N__11191));
    IoSpan4Mux I__2621 (
            .O(N__11195),
            .I(N__11186));
    InMux I__2620 (
            .O(N__11194),
            .I(N__11183));
    InMux I__2619 (
            .O(N__11191),
            .I(N__11178));
    InMux I__2618 (
            .O(N__11190),
            .I(N__11178));
    InMux I__2617 (
            .O(N__11189),
            .I(N__11175));
    Span4Mux_s2_v I__2616 (
            .O(N__11186),
            .I(N__11172));
    LocalMux I__2615 (
            .O(N__11183),
            .I(N__11165));
    LocalMux I__2614 (
            .O(N__11178),
            .I(N__11165));
    LocalMux I__2613 (
            .O(N__11175),
            .I(N__11165));
    Sp12to4 I__2612 (
            .O(N__11172),
            .I(N__11162));
    Span4Mux_v I__2611 (
            .O(N__11165),
            .I(N__11159));
    Span12Mux_v I__2610 (
            .O(N__11162),
            .I(N__11155));
    Span4Mux_h I__2609 (
            .O(N__11159),
            .I(N__11152));
    InMux I__2608 (
            .O(N__11158),
            .I(N__11149));
    Odrv12 I__2607 (
            .O(N__11155),
            .I(DBENn_c));
    Odrv4 I__2606 (
            .O(N__11152),
            .I(DBENn_c));
    LocalMux I__2605 (
            .O(N__11149),
            .I(DBENn_c));
    CascadeMux I__2604 (
            .O(N__11142),
            .I(N__11136));
    InMux I__2603 (
            .O(N__11141),
            .I(N__11133));
    InMux I__2602 (
            .O(N__11140),
            .I(N__11130));
    InMux I__2601 (
            .O(N__11139),
            .I(N__11127));
    InMux I__2600 (
            .O(N__11136),
            .I(N__11123));
    LocalMux I__2599 (
            .O(N__11133),
            .I(N__11118));
    LocalMux I__2598 (
            .O(N__11130),
            .I(N__11118));
    LocalMux I__2597 (
            .O(N__11127),
            .I(N__11115));
    InMux I__2596 (
            .O(N__11126),
            .I(N__11112));
    LocalMux I__2595 (
            .O(N__11123),
            .I(N__11108));
    Span4Mux_h I__2594 (
            .O(N__11118),
            .I(N__11101));
    Span4Mux_v I__2593 (
            .O(N__11115),
            .I(N__11101));
    LocalMux I__2592 (
            .O(N__11112),
            .I(N__11101));
    InMux I__2591 (
            .O(N__11111),
            .I(N__11098));
    Span4Mux_v I__2590 (
            .O(N__11108),
            .I(N__11094));
    Span4Mux_h I__2589 (
            .O(N__11101),
            .I(N__11089));
    LocalMux I__2588 (
            .O(N__11098),
            .I(N__11089));
    InMux I__2587 (
            .O(N__11097),
            .I(N__11085));
    Span4Mux_h I__2586 (
            .O(N__11094),
            .I(N__11082));
    Span4Mux_h I__2585 (
            .O(N__11089),
            .I(N__11079));
    InMux I__2584 (
            .O(N__11088),
            .I(N__11076));
    LocalMux I__2583 (
            .O(N__11085),
            .I(N__11073));
    Odrv4 I__2582 (
            .O(N__11082),
            .I(DMA_CYCLEm));
    Odrv4 I__2581 (
            .O(N__11079),
            .I(DMA_CYCLEm));
    LocalMux I__2580 (
            .O(N__11076),
            .I(DMA_CYCLEm));
    Odrv4 I__2579 (
            .O(N__11073),
            .I(DMA_CYCLEm));
    InMux I__2578 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__2577 (
            .O(N__11061),
            .I(\U712_BYTE_ENABLE.N_456 ));
    IoInMux I__2576 (
            .O(N__11058),
            .I(N__11055));
    LocalMux I__2575 (
            .O(N__11055),
            .I(N__11052));
    Span4Mux_s0_v I__2574 (
            .O(N__11052),
            .I(N__11049));
    Span4Mux_v I__2573 (
            .O(N__11049),
            .I(N__11046));
    Odrv4 I__2572 (
            .O(N__11046),
            .I(N_412_i));
    CascadeMux I__2571 (
            .O(N__11043),
            .I(N__11039));
    InMux I__2570 (
            .O(N__11042),
            .I(N__11030));
    InMux I__2569 (
            .O(N__11039),
            .I(N__11027));
    InMux I__2568 (
            .O(N__11038),
            .I(N__11024));
    InMux I__2567 (
            .O(N__11037),
            .I(N__11021));
    InMux I__2566 (
            .O(N__11036),
            .I(N__11016));
    CascadeMux I__2565 (
            .O(N__11035),
            .I(N__11011));
    CascadeMux I__2564 (
            .O(N__11034),
            .I(N__11007));
    CascadeMux I__2563 (
            .O(N__11033),
            .I(N__11002));
    LocalMux I__2562 (
            .O(N__11030),
            .I(N__10998));
    LocalMux I__2561 (
            .O(N__11027),
            .I(N__10995));
    LocalMux I__2560 (
            .O(N__11024),
            .I(N__10989));
    LocalMux I__2559 (
            .O(N__11021),
            .I(N__10989));
    InMux I__2558 (
            .O(N__11020),
            .I(N__10986));
    InMux I__2557 (
            .O(N__11019),
            .I(N__10983));
    LocalMux I__2556 (
            .O(N__11016),
            .I(N__10977));
    InMux I__2555 (
            .O(N__11015),
            .I(N__10974));
    InMux I__2554 (
            .O(N__11014),
            .I(N__10963));
    InMux I__2553 (
            .O(N__11011),
            .I(N__10963));
    InMux I__2552 (
            .O(N__11010),
            .I(N__10963));
    InMux I__2551 (
            .O(N__11007),
            .I(N__10963));
    InMux I__2550 (
            .O(N__11006),
            .I(N__10963));
    InMux I__2549 (
            .O(N__11005),
            .I(N__10960));
    InMux I__2548 (
            .O(N__11002),
            .I(N__10955));
    InMux I__2547 (
            .O(N__11001),
            .I(N__10955));
    Span4Mux_v I__2546 (
            .O(N__10998),
            .I(N__10950));
    Span4Mux_v I__2545 (
            .O(N__10995),
            .I(N__10950));
    InMux I__2544 (
            .O(N__10994),
            .I(N__10947));
    Span4Mux_h I__2543 (
            .O(N__10989),
            .I(N__10940));
    LocalMux I__2542 (
            .O(N__10986),
            .I(N__10940));
    LocalMux I__2541 (
            .O(N__10983),
            .I(N__10940));
    InMux I__2540 (
            .O(N__10982),
            .I(N__10937));
    InMux I__2539 (
            .O(N__10981),
            .I(N__10934));
    InMux I__2538 (
            .O(N__10980),
            .I(N__10931));
    Span4Mux_v I__2537 (
            .O(N__10977),
            .I(N__10928));
    LocalMux I__2536 (
            .O(N__10974),
            .I(N__10919));
    LocalMux I__2535 (
            .O(N__10963),
            .I(N__10919));
    LocalMux I__2534 (
            .O(N__10960),
            .I(N__10919));
    LocalMux I__2533 (
            .O(N__10955),
            .I(N__10919));
    Sp12to4 I__2532 (
            .O(N__10950),
            .I(N__10915));
    LocalMux I__2531 (
            .O(N__10947),
            .I(N__10904));
    Span4Mux_h I__2530 (
            .O(N__10940),
            .I(N__10904));
    LocalMux I__2529 (
            .O(N__10937),
            .I(N__10904));
    LocalMux I__2528 (
            .O(N__10934),
            .I(N__10904));
    LocalMux I__2527 (
            .O(N__10931),
            .I(N__10904));
    Span4Mux_h I__2526 (
            .O(N__10928),
            .I(N__10899));
    Span4Mux_v I__2525 (
            .O(N__10919),
            .I(N__10899));
    InMux I__2524 (
            .O(N__10918),
            .I(N__10896));
    Span12Mux_h I__2523 (
            .O(N__10915),
            .I(N__10891));
    Sp12to4 I__2522 (
            .O(N__10904),
            .I(N__10891));
    Sp12to4 I__2521 (
            .O(N__10899),
            .I(N__10888));
    LocalMux I__2520 (
            .O(N__10896),
            .I(N__10885));
    Span12Mux_v I__2519 (
            .O(N__10891),
            .I(N__10882));
    Span12Mux_h I__2518 (
            .O(N__10888),
            .I(N__10879));
    Span12Mux_v I__2517 (
            .O(N__10885),
            .I(N__10876));
    Span12Mux_h I__2516 (
            .O(N__10882),
            .I(N__10873));
    Span12Mux_v I__2515 (
            .O(N__10879),
            .I(N__10868));
    Span12Mux_h I__2514 (
            .O(N__10876),
            .I(N__10868));
    Odrv12 I__2513 (
            .O(N__10873),
            .I(AGNUS_REV_c));
    Odrv12 I__2512 (
            .O(N__10868),
            .I(AGNUS_REV_c));
    InMux I__2511 (
            .O(N__10863),
            .I(N__10858));
    InMux I__2510 (
            .O(N__10862),
            .I(N__10855));
    InMux I__2509 (
            .O(N__10861),
            .I(N__10851));
    LocalMux I__2508 (
            .O(N__10858),
            .I(N__10848));
    LocalMux I__2507 (
            .O(N__10855),
            .I(N__10845));
    InMux I__2506 (
            .O(N__10854),
            .I(N__10842));
    LocalMux I__2505 (
            .O(N__10851),
            .I(N__10839));
    Span4Mux_v I__2504 (
            .O(N__10848),
            .I(N__10836));
    Span4Mux_h I__2503 (
            .O(N__10845),
            .I(N__10831));
    LocalMux I__2502 (
            .O(N__10842),
            .I(N__10831));
    Span4Mux_v I__2501 (
            .O(N__10839),
            .I(N__10828));
    Span4Mux_h I__2500 (
            .O(N__10836),
            .I(N__10823));
    Span4Mux_v I__2499 (
            .O(N__10831),
            .I(N__10823));
    Sp12to4 I__2498 (
            .O(N__10828),
            .I(N__10820));
    Sp12to4 I__2497 (
            .O(N__10823),
            .I(N__10817));
    Span12Mux_h I__2496 (
            .O(N__10820),
            .I(N__10814));
    Span12Mux_h I__2495 (
            .O(N__10817),
            .I(N__10811));
    Span12Mux_v I__2494 (
            .O(N__10814),
            .I(N__10808));
    Span12Mux_v I__2493 (
            .O(N__10811),
            .I(N__10805));
    Odrv12 I__2492 (
            .O(N__10808),
            .I(DRA_c_9));
    Odrv12 I__2491 (
            .O(N__10805),
            .I(DRA_c_9));
    InMux I__2490 (
            .O(N__10800),
            .I(N__10797));
    LocalMux I__2489 (
            .O(N__10797),
            .I(N__10794));
    Odrv12 I__2488 (
            .O(N__10794),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2487 (
            .O(N__10791),
            .I(N__10773));
    ClkMux I__2486 (
            .O(N__10790),
            .I(N__10773));
    ClkMux I__2485 (
            .O(N__10789),
            .I(N__10773));
    ClkMux I__2484 (
            .O(N__10788),
            .I(N__10773));
    ClkMux I__2483 (
            .O(N__10787),
            .I(N__10773));
    ClkMux I__2482 (
            .O(N__10786),
            .I(N__10773));
    GlobalMux I__2481 (
            .O(N__10773),
            .I(N__10770));
    gio2CtrlBuf I__2480 (
            .O(N__10770),
            .I(C3_c_g));
    CEMux I__2479 (
            .O(N__10767),
            .I(N__10731));
    CEMux I__2478 (
            .O(N__10766),
            .I(N__10731));
    CEMux I__2477 (
            .O(N__10765),
            .I(N__10731));
    CEMux I__2476 (
            .O(N__10764),
            .I(N__10731));
    CEMux I__2475 (
            .O(N__10763),
            .I(N__10731));
    CEMux I__2474 (
            .O(N__10762),
            .I(N__10731));
    CEMux I__2473 (
            .O(N__10761),
            .I(N__10731));
    CEMux I__2472 (
            .O(N__10760),
            .I(N__10731));
    CEMux I__2471 (
            .O(N__10759),
            .I(N__10731));
    CEMux I__2470 (
            .O(N__10758),
            .I(N__10731));
    CEMux I__2469 (
            .O(N__10757),
            .I(N__10731));
    CEMux I__2468 (
            .O(N__10756),
            .I(N__10731));
    GlobalMux I__2467 (
            .O(N__10731),
            .I(N__10728));
    gio2CtrlBuf I__2466 (
            .O(N__10728),
            .I(DBRn_c_i_0_g));
    InMux I__2465 (
            .O(N__10725),
            .I(N__10715));
    InMux I__2464 (
            .O(N__10724),
            .I(N__10712));
    InMux I__2463 (
            .O(N__10723),
            .I(N__10709));
    InMux I__2462 (
            .O(N__10722),
            .I(N__10704));
    InMux I__2461 (
            .O(N__10721),
            .I(N__10704));
    InMux I__2460 (
            .O(N__10720),
            .I(N__10699));
    InMux I__2459 (
            .O(N__10719),
            .I(N__10699));
    InMux I__2458 (
            .O(N__10718),
            .I(N__10696));
    LocalMux I__2457 (
            .O(N__10715),
            .I(N__10693));
    LocalMux I__2456 (
            .O(N__10712),
            .I(N__10678));
    LocalMux I__2455 (
            .O(N__10709),
            .I(N__10669));
    LocalMux I__2454 (
            .O(N__10704),
            .I(N__10661));
    LocalMux I__2453 (
            .O(N__10699),
            .I(N__10658));
    LocalMux I__2452 (
            .O(N__10696),
            .I(N__10643));
    Glb2LocalMux I__2451 (
            .O(N__10693),
            .I(N__10557));
    SRMux I__2450 (
            .O(N__10692),
            .I(N__10557));
    SRMux I__2449 (
            .O(N__10691),
            .I(N__10557));
    SRMux I__2448 (
            .O(N__10690),
            .I(N__10557));
    SRMux I__2447 (
            .O(N__10689),
            .I(N__10557));
    SRMux I__2446 (
            .O(N__10688),
            .I(N__10557));
    SRMux I__2445 (
            .O(N__10687),
            .I(N__10557));
    SRMux I__2444 (
            .O(N__10686),
            .I(N__10557));
    SRMux I__2443 (
            .O(N__10685),
            .I(N__10557));
    SRMux I__2442 (
            .O(N__10684),
            .I(N__10557));
    SRMux I__2441 (
            .O(N__10683),
            .I(N__10557));
    SRMux I__2440 (
            .O(N__10682),
            .I(N__10557));
    SRMux I__2439 (
            .O(N__10681),
            .I(N__10557));
    Glb2LocalMux I__2438 (
            .O(N__10678),
            .I(N__10557));
    SRMux I__2437 (
            .O(N__10677),
            .I(N__10557));
    SRMux I__2436 (
            .O(N__10676),
            .I(N__10557));
    SRMux I__2435 (
            .O(N__10675),
            .I(N__10557));
    SRMux I__2434 (
            .O(N__10674),
            .I(N__10557));
    SRMux I__2433 (
            .O(N__10673),
            .I(N__10557));
    SRMux I__2432 (
            .O(N__10672),
            .I(N__10557));
    Glb2LocalMux I__2431 (
            .O(N__10669),
            .I(N__10557));
    SRMux I__2430 (
            .O(N__10668),
            .I(N__10557));
    SRMux I__2429 (
            .O(N__10667),
            .I(N__10557));
    SRMux I__2428 (
            .O(N__10666),
            .I(N__10557));
    SRMux I__2427 (
            .O(N__10665),
            .I(N__10557));
    SRMux I__2426 (
            .O(N__10664),
            .I(N__10557));
    Glb2LocalMux I__2425 (
            .O(N__10661),
            .I(N__10557));
    Glb2LocalMux I__2424 (
            .O(N__10658),
            .I(N__10557));
    SRMux I__2423 (
            .O(N__10657),
            .I(N__10557));
    SRMux I__2422 (
            .O(N__10656),
            .I(N__10557));
    SRMux I__2421 (
            .O(N__10655),
            .I(N__10557));
    SRMux I__2420 (
            .O(N__10654),
            .I(N__10557));
    SRMux I__2419 (
            .O(N__10653),
            .I(N__10557));
    SRMux I__2418 (
            .O(N__10652),
            .I(N__10557));
    SRMux I__2417 (
            .O(N__10651),
            .I(N__10557));
    SRMux I__2416 (
            .O(N__10650),
            .I(N__10557));
    SRMux I__2415 (
            .O(N__10649),
            .I(N__10557));
    SRMux I__2414 (
            .O(N__10648),
            .I(N__10557));
    SRMux I__2413 (
            .O(N__10647),
            .I(N__10557));
    SRMux I__2412 (
            .O(N__10646),
            .I(N__10557));
    Glb2LocalMux I__2411 (
            .O(N__10643),
            .I(N__10557));
    SRMux I__2410 (
            .O(N__10642),
            .I(N__10557));
    GlobalMux I__2409 (
            .O(N__10557),
            .I(N__10554));
    gio2CtrlBuf I__2408 (
            .O(N__10554),
            .I(RESETn_c_i_g));
    InMux I__2407 (
            .O(N__10551),
            .I(N__10547));
    InMux I__2406 (
            .O(N__10550),
            .I(N__10544));
    LocalMux I__2405 (
            .O(N__10547),
            .I(N__10539));
    LocalMux I__2404 (
            .O(N__10544),
            .I(N__10539));
    Span4Mux_v I__2403 (
            .O(N__10539),
            .I(N__10536));
    Sp12to4 I__2402 (
            .O(N__10536),
            .I(N__10533));
    Span12Mux_h I__2401 (
            .O(N__10533),
            .I(N__10530));
    Odrv12 I__2400 (
            .O(N__10530),
            .I(RAS0n_c));
    InMux I__2399 (
            .O(N__10527),
            .I(N__10524));
    LocalMux I__2398 (
            .O(N__10524),
            .I(N__10521));
    Sp12to4 I__2397 (
            .O(N__10521),
            .I(N__10518));
    Span12Mux_v I__2396 (
            .O(N__10518),
            .I(N__10515));
    Span12Mux_h I__2395 (
            .O(N__10515),
            .I(N__10512));
    Odrv12 I__2394 (
            .O(N__10512),
            .I(RAS1n_c));
    InMux I__2393 (
            .O(N__10509),
            .I(N__10493));
    InMux I__2392 (
            .O(N__10508),
            .I(N__10488));
    InMux I__2391 (
            .O(N__10507),
            .I(N__10488));
    InMux I__2390 (
            .O(N__10506),
            .I(N__10485));
    InMux I__2389 (
            .O(N__10505),
            .I(N__10480));
    InMux I__2388 (
            .O(N__10504),
            .I(N__10480));
    InMux I__2387 (
            .O(N__10503),
            .I(N__10473));
    CascadeMux I__2386 (
            .O(N__10502),
            .I(N__10468));
    InMux I__2385 (
            .O(N__10501),
            .I(N__10461));
    InMux I__2384 (
            .O(N__10500),
            .I(N__10461));
    InMux I__2383 (
            .O(N__10499),
            .I(N__10461));
    InMux I__2382 (
            .O(N__10498),
            .I(N__10456));
    InMux I__2381 (
            .O(N__10497),
            .I(N__10456));
    InMux I__2380 (
            .O(N__10496),
            .I(N__10447));
    LocalMux I__2379 (
            .O(N__10493),
            .I(N__10436));
    LocalMux I__2378 (
            .O(N__10488),
            .I(N__10436));
    LocalMux I__2377 (
            .O(N__10485),
            .I(N__10436));
    LocalMux I__2376 (
            .O(N__10480),
            .I(N__10436));
    InMux I__2375 (
            .O(N__10479),
            .I(N__10431));
    InMux I__2374 (
            .O(N__10478),
            .I(N__10431));
    InMux I__2373 (
            .O(N__10477),
            .I(N__10426));
    InMux I__2372 (
            .O(N__10476),
            .I(N__10426));
    LocalMux I__2371 (
            .O(N__10473),
            .I(N__10422));
    InMux I__2370 (
            .O(N__10472),
            .I(N__10417));
    InMux I__2369 (
            .O(N__10471),
            .I(N__10417));
    InMux I__2368 (
            .O(N__10468),
            .I(N__10414));
    LocalMux I__2367 (
            .O(N__10461),
            .I(N__10409));
    LocalMux I__2366 (
            .O(N__10456),
            .I(N__10409));
    InMux I__2365 (
            .O(N__10455),
            .I(N__10398));
    InMux I__2364 (
            .O(N__10454),
            .I(N__10398));
    InMux I__2363 (
            .O(N__10453),
            .I(N__10398));
    InMux I__2362 (
            .O(N__10452),
            .I(N__10398));
    InMux I__2361 (
            .O(N__10451),
            .I(N__10398));
    CascadeMux I__2360 (
            .O(N__10450),
            .I(N__10395));
    LocalMux I__2359 (
            .O(N__10447),
            .I(N__10391));
    InMux I__2358 (
            .O(N__10446),
            .I(N__10386));
    InMux I__2357 (
            .O(N__10445),
            .I(N__10386));
    Span4Mux_v I__2356 (
            .O(N__10436),
            .I(N__10379));
    LocalMux I__2355 (
            .O(N__10431),
            .I(N__10379));
    LocalMux I__2354 (
            .O(N__10426),
            .I(N__10379));
    InMux I__2353 (
            .O(N__10425),
            .I(N__10376));
    Span4Mux_v I__2352 (
            .O(N__10422),
            .I(N__10366));
    LocalMux I__2351 (
            .O(N__10417),
            .I(N__10366));
    LocalMux I__2350 (
            .O(N__10414),
            .I(N__10366));
    Span4Mux_v I__2349 (
            .O(N__10409),
            .I(N__10360));
    LocalMux I__2348 (
            .O(N__10398),
            .I(N__10360));
    InMux I__2347 (
            .O(N__10395),
            .I(N__10357));
    InMux I__2346 (
            .O(N__10394),
            .I(N__10354));
    Span4Mux_v I__2345 (
            .O(N__10391),
            .I(N__10341));
    LocalMux I__2344 (
            .O(N__10386),
            .I(N__10341));
    Span4Mux_v I__2343 (
            .O(N__10379),
            .I(N__10336));
    LocalMux I__2342 (
            .O(N__10376),
            .I(N__10336));
    InMux I__2341 (
            .O(N__10375),
            .I(N__10331));
    InMux I__2340 (
            .O(N__10374),
            .I(N__10331));
    InMux I__2339 (
            .O(N__10373),
            .I(N__10328));
    Span4Mux_v I__2338 (
            .O(N__10366),
            .I(N__10325));
    InMux I__2337 (
            .O(N__10365),
            .I(N__10322));
    Span4Mux_h I__2336 (
            .O(N__10360),
            .I(N__10315));
    LocalMux I__2335 (
            .O(N__10357),
            .I(N__10315));
    LocalMux I__2334 (
            .O(N__10354),
            .I(N__10315));
    InMux I__2333 (
            .O(N__10353),
            .I(N__10310));
    InMux I__2332 (
            .O(N__10352),
            .I(N__10310));
    InMux I__2331 (
            .O(N__10351),
            .I(N__10297));
    InMux I__2330 (
            .O(N__10350),
            .I(N__10297));
    InMux I__2329 (
            .O(N__10349),
            .I(N__10297));
    InMux I__2328 (
            .O(N__10348),
            .I(N__10297));
    InMux I__2327 (
            .O(N__10347),
            .I(N__10297));
    InMux I__2326 (
            .O(N__10346),
            .I(N__10297));
    Span4Mux_h I__2325 (
            .O(N__10341),
            .I(N__10292));
    Span4Mux_v I__2324 (
            .O(N__10336),
            .I(N__10292));
    LocalMux I__2323 (
            .O(N__10331),
            .I(N__10289));
    LocalMux I__2322 (
            .O(N__10328),
            .I(N__10286));
    Span4Mux_h I__2321 (
            .O(N__10325),
            .I(N__10282));
    LocalMux I__2320 (
            .O(N__10322),
            .I(N__10273));
    Sp12to4 I__2319 (
            .O(N__10315),
            .I(N__10273));
    LocalMux I__2318 (
            .O(N__10310),
            .I(N__10273));
    LocalMux I__2317 (
            .O(N__10297),
            .I(N__10273));
    Span4Mux_h I__2316 (
            .O(N__10292),
            .I(N__10266));
    Span4Mux_v I__2315 (
            .O(N__10289),
            .I(N__10266));
    Span4Mux_v I__2314 (
            .O(N__10286),
            .I(N__10266));
    InMux I__2313 (
            .O(N__10285),
            .I(N__10263));
    Sp12to4 I__2312 (
            .O(N__10282),
            .I(N__10254));
    Span12Mux_v I__2311 (
            .O(N__10273),
            .I(N__10254));
    Sp12to4 I__2310 (
            .O(N__10266),
            .I(N__10254));
    LocalMux I__2309 (
            .O(N__10263),
            .I(N__10254));
    Span12Mux_h I__2308 (
            .O(N__10254),
            .I(N__10251));
    Odrv12 I__2307 (
            .O(N__10251),
            .I(RESETn_c));
    InMux I__2306 (
            .O(N__10248),
            .I(N__10245));
    LocalMux I__2305 (
            .O(N__10245),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2304 (
            .O(N__10242),
            .I(N__10239));
    LocalMux I__2303 (
            .O(N__10239),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2302 (
            .O(N__10236),
            .I(N__10233));
    LocalMux I__2301 (
            .O(N__10233),
            .I(N__10188));
    ClkMux I__2300 (
            .O(N__10232),
            .I(N__10095));
    ClkMux I__2299 (
            .O(N__10231),
            .I(N__10095));
    ClkMux I__2298 (
            .O(N__10230),
            .I(N__10095));
    ClkMux I__2297 (
            .O(N__10229),
            .I(N__10095));
    ClkMux I__2296 (
            .O(N__10228),
            .I(N__10095));
    ClkMux I__2295 (
            .O(N__10227),
            .I(N__10095));
    ClkMux I__2294 (
            .O(N__10226),
            .I(N__10095));
    ClkMux I__2293 (
            .O(N__10225),
            .I(N__10095));
    ClkMux I__2292 (
            .O(N__10224),
            .I(N__10095));
    ClkMux I__2291 (
            .O(N__10223),
            .I(N__10095));
    ClkMux I__2290 (
            .O(N__10222),
            .I(N__10095));
    ClkMux I__2289 (
            .O(N__10221),
            .I(N__10095));
    ClkMux I__2288 (
            .O(N__10220),
            .I(N__10095));
    ClkMux I__2287 (
            .O(N__10219),
            .I(N__10095));
    ClkMux I__2286 (
            .O(N__10218),
            .I(N__10095));
    ClkMux I__2285 (
            .O(N__10217),
            .I(N__10095));
    ClkMux I__2284 (
            .O(N__10216),
            .I(N__10095));
    ClkMux I__2283 (
            .O(N__10215),
            .I(N__10095));
    ClkMux I__2282 (
            .O(N__10214),
            .I(N__10095));
    ClkMux I__2281 (
            .O(N__10213),
            .I(N__10095));
    ClkMux I__2280 (
            .O(N__10212),
            .I(N__10095));
    ClkMux I__2279 (
            .O(N__10211),
            .I(N__10095));
    ClkMux I__2278 (
            .O(N__10210),
            .I(N__10095));
    ClkMux I__2277 (
            .O(N__10209),
            .I(N__10095));
    ClkMux I__2276 (
            .O(N__10208),
            .I(N__10095));
    ClkMux I__2275 (
            .O(N__10207),
            .I(N__10095));
    ClkMux I__2274 (
            .O(N__10206),
            .I(N__10095));
    ClkMux I__2273 (
            .O(N__10205),
            .I(N__10095));
    ClkMux I__2272 (
            .O(N__10204),
            .I(N__10095));
    ClkMux I__2271 (
            .O(N__10203),
            .I(N__10095));
    ClkMux I__2270 (
            .O(N__10202),
            .I(N__10095));
    ClkMux I__2269 (
            .O(N__10201),
            .I(N__10095));
    ClkMux I__2268 (
            .O(N__10200),
            .I(N__10095));
    ClkMux I__2267 (
            .O(N__10199),
            .I(N__10095));
    ClkMux I__2266 (
            .O(N__10198),
            .I(N__10095));
    ClkMux I__2265 (
            .O(N__10197),
            .I(N__10095));
    ClkMux I__2264 (
            .O(N__10196),
            .I(N__10095));
    ClkMux I__2263 (
            .O(N__10195),
            .I(N__10095));
    ClkMux I__2262 (
            .O(N__10194),
            .I(N__10095));
    ClkMux I__2261 (
            .O(N__10193),
            .I(N__10095));
    ClkMux I__2260 (
            .O(N__10192),
            .I(N__10095));
    ClkMux I__2259 (
            .O(N__10191),
            .I(N__10095));
    Glb2LocalMux I__2258 (
            .O(N__10188),
            .I(N__10095));
    ClkMux I__2257 (
            .O(N__10187),
            .I(N__10095));
    ClkMux I__2256 (
            .O(N__10186),
            .I(N__10095));
    GlobalMux I__2255 (
            .O(N__10095),
            .I(CLK80_PLL));
    InMux I__2254 (
            .O(N__10092),
            .I(N__10089));
    LocalMux I__2253 (
            .O(N__10089),
            .I(\U712_BYTE_ENABLE.N_467 ));
    CascadeMux I__2252 (
            .O(N__10086),
            .I(\U712_BYTE_ENABLE.N_455_cascade_ ));
    IoInMux I__2251 (
            .O(N__10083),
            .I(N__10080));
    LocalMux I__2250 (
            .O(N__10080),
            .I(N__10077));
    IoSpan4Mux I__2249 (
            .O(N__10077),
            .I(N__10074));
    IoSpan4Mux I__2248 (
            .O(N__10074),
            .I(N__10071));
    Span4Mux_s2_v I__2247 (
            .O(N__10071),
            .I(N__10068));
    Sp12to4 I__2246 (
            .O(N__10068),
            .I(N__10065));
    Span12Mux_v I__2245 (
            .O(N__10065),
            .I(N__10062));
    Odrv12 I__2244 (
            .O(N__10062),
            .I(N_38_i));
    InMux I__2243 (
            .O(N__10059),
            .I(N__10056));
    LocalMux I__2242 (
            .O(N__10056),
            .I(N__10053));
    Odrv4 I__2241 (
            .O(N__10053),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    InMux I__2240 (
            .O(N__10050),
            .I(N__10046));
    InMux I__2239 (
            .O(N__10049),
            .I(N__10043));
    LocalMux I__2238 (
            .O(N__10046),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__2237 (
            .O(N__10043),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__2236 (
            .O(N__10038),
            .I(N__10034));
    InMux I__2235 (
            .O(N__10037),
            .I(N__10031));
    LocalMux I__2234 (
            .O(N__10034),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__2233 (
            .O(N__10031),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__2232 (
            .O(N__10026),
            .I(N__10023));
    LocalMux I__2231 (
            .O(N__10023),
            .I(N__10020));
    Odrv4 I__2230 (
            .O(N__10020),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__2229 (
            .O(N__10017),
            .I(N__10014));
    LocalMux I__2228 (
            .O(N__10014),
            .I(N__10011));
    Span4Mux_v I__2227 (
            .O(N__10011),
            .I(N__10005));
    InMux I__2226 (
            .O(N__10010),
            .I(N__10000));
    InMux I__2225 (
            .O(N__10009),
            .I(N__10000));
    InMux I__2224 (
            .O(N__10008),
            .I(N__9997));
    Span4Mux_h I__2223 (
            .O(N__10005),
            .I(N__9989));
    LocalMux I__2222 (
            .O(N__10000),
            .I(N__9989));
    LocalMux I__2221 (
            .O(N__9997),
            .I(N__9989));
    InMux I__2220 (
            .O(N__9996),
            .I(N__9986));
    Span4Mux_h I__2219 (
            .O(N__9989),
            .I(N__9983));
    LocalMux I__2218 (
            .O(N__9986),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2217 (
            .O(N__9983),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2216 (
            .O(N__9978),
            .I(N__9975));
    LocalMux I__2215 (
            .O(N__9975),
            .I(N__9972));
    IoSpan4Mux I__2214 (
            .O(N__9972),
            .I(N__9969));
    Sp12to4 I__2213 (
            .O(N__9969),
            .I(N__9966));
    Span12Mux_s9_v I__2212 (
            .O(N__9966),
            .I(N__9963));
    Span12Mux_h I__2211 (
            .O(N__9963),
            .I(N__9960));
    Odrv12 I__2210 (
            .O(N__9960),
            .I(WEn_c));
    InMux I__2209 (
            .O(N__9957),
            .I(N__9952));
    InMux I__2208 (
            .O(N__9956),
            .I(N__9949));
    InMux I__2207 (
            .O(N__9955),
            .I(N__9945));
    LocalMux I__2206 (
            .O(N__9952),
            .I(N__9940));
    LocalMux I__2205 (
            .O(N__9949),
            .I(N__9940));
    InMux I__2204 (
            .O(N__9948),
            .I(N__9937));
    LocalMux I__2203 (
            .O(N__9945),
            .I(N__9934));
    Span4Mux_v I__2202 (
            .O(N__9940),
            .I(N__9931));
    LocalMux I__2201 (
            .O(N__9937),
            .I(N__9928));
    Span4Mux_v I__2200 (
            .O(N__9934),
            .I(N__9925));
    Span4Mux_h I__2199 (
            .O(N__9931),
            .I(N__9920));
    Span4Mux_h I__2198 (
            .O(N__9928),
            .I(N__9920));
    Span4Mux_v I__2197 (
            .O(N__9925),
            .I(N__9917));
    Span4Mux_v I__2196 (
            .O(N__9920),
            .I(N__9914));
    Sp12to4 I__2195 (
            .O(N__9917),
            .I(N__9909));
    Sp12to4 I__2194 (
            .O(N__9914),
            .I(N__9909));
    Span12Mux_h I__2193 (
            .O(N__9909),
            .I(N__9906));
    Odrv12 I__2192 (
            .O(N__9906),
            .I(DRA_c_4));
    CascadeMux I__2191 (
            .O(N__9903),
            .I(N__9900));
    InMux I__2190 (
            .O(N__9900),
            .I(N__9897));
    LocalMux I__2189 (
            .O(N__9897),
            .I(N__9894));
    Span4Mux_h I__2188 (
            .O(N__9894),
            .I(N__9891));
    Odrv4 I__2187 (
            .O(N__9891),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2186 (
            .O(N__9888),
            .I(N__9884));
    InMux I__2185 (
            .O(N__9887),
            .I(N__9881));
    LocalMux I__2184 (
            .O(N__9884),
            .I(N__9875));
    LocalMux I__2183 (
            .O(N__9881),
            .I(N__9875));
    InMux I__2182 (
            .O(N__9880),
            .I(N__9872));
    Span4Mux_h I__2181 (
            .O(N__9875),
            .I(N__9868));
    LocalMux I__2180 (
            .O(N__9872),
            .I(N__9865));
    InMux I__2179 (
            .O(N__9871),
            .I(N__9862));
    Span4Mux_v I__2178 (
            .O(N__9868),
            .I(N__9859));
    Sp12to4 I__2177 (
            .O(N__9865),
            .I(N__9854));
    LocalMux I__2176 (
            .O(N__9862),
            .I(N__9854));
    Sp12to4 I__2175 (
            .O(N__9859),
            .I(N__9849));
    Span12Mux_v I__2174 (
            .O(N__9854),
            .I(N__9849));
    Span12Mux_h I__2173 (
            .O(N__9849),
            .I(N__9846));
    Odrv12 I__2172 (
            .O(N__9846),
            .I(DRA_c_6));
    InMux I__2171 (
            .O(N__9843),
            .I(N__9840));
    LocalMux I__2170 (
            .O(N__9840),
            .I(N__9834));
    InMux I__2169 (
            .O(N__9839),
            .I(N__9831));
    InMux I__2168 (
            .O(N__9838),
            .I(N__9828));
    InMux I__2167 (
            .O(N__9837),
            .I(N__9825));
    Span4Mux_v I__2166 (
            .O(N__9834),
            .I(N__9820));
    LocalMux I__2165 (
            .O(N__9831),
            .I(N__9820));
    LocalMux I__2164 (
            .O(N__9828),
            .I(N__9815));
    LocalMux I__2163 (
            .O(N__9825),
            .I(N__9815));
    Span4Mux_v I__2162 (
            .O(N__9820),
            .I(N__9812));
    Span12Mux_v I__2161 (
            .O(N__9815),
            .I(N__9807));
    Sp12to4 I__2160 (
            .O(N__9812),
            .I(N__9807));
    Span12Mux_h I__2159 (
            .O(N__9807),
            .I(N__9804));
    Odrv12 I__2158 (
            .O(N__9804),
            .I(DRA_c_5));
    CascadeMux I__2157 (
            .O(N__9801),
            .I(N__9798));
    InMux I__2156 (
            .O(N__9798),
            .I(N__9795));
    LocalMux I__2155 (
            .O(N__9795),
            .I(N__9792));
    Odrv4 I__2154 (
            .O(N__9792),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2153 (
            .O(N__9789),
            .I(N__9784));
    InMux I__2152 (
            .O(N__9788),
            .I(N__9779));
    InMux I__2151 (
            .O(N__9787),
            .I(N__9779));
    LocalMux I__2150 (
            .O(N__9784),
            .I(N__9774));
    LocalMux I__2149 (
            .O(N__9779),
            .I(N__9774));
    Span4Mux_v I__2148 (
            .O(N__9774),
            .I(N__9770));
    InMux I__2147 (
            .O(N__9773),
            .I(N__9767));
    Span4Mux_v I__2146 (
            .O(N__9770),
            .I(N__9764));
    LocalMux I__2145 (
            .O(N__9767),
            .I(N__9761));
    Sp12to4 I__2144 (
            .O(N__9764),
            .I(N__9756));
    Span12Mux_v I__2143 (
            .O(N__9761),
            .I(N__9756));
    Span12Mux_h I__2142 (
            .O(N__9756),
            .I(N__9753));
    Odrv12 I__2141 (
            .O(N__9753),
            .I(DRA_c_3));
    InMux I__2140 (
            .O(N__9750),
            .I(N__9746));
    InMux I__2139 (
            .O(N__9749),
            .I(N__9743));
    LocalMux I__2138 (
            .O(N__9746),
            .I(N__9737));
    LocalMux I__2137 (
            .O(N__9743),
            .I(N__9737));
    InMux I__2136 (
            .O(N__9742),
            .I(N__9734));
    Span4Mux_v I__2135 (
            .O(N__9737),
            .I(N__9729));
    LocalMux I__2134 (
            .O(N__9734),
            .I(N__9729));
    Span4Mux_v I__2133 (
            .O(N__9729),
            .I(N__9725));
    InMux I__2132 (
            .O(N__9728),
            .I(N__9722));
    Span4Mux_v I__2131 (
            .O(N__9725),
            .I(N__9719));
    LocalMux I__2130 (
            .O(N__9722),
            .I(N__9716));
    Sp12to4 I__2129 (
            .O(N__9719),
            .I(N__9711));
    Span12Mux_v I__2128 (
            .O(N__9716),
            .I(N__9711));
    Span12Mux_h I__2127 (
            .O(N__9711),
            .I(N__9708));
    Odrv12 I__2126 (
            .O(N__9708),
            .I(DRA_c_2));
    InMux I__2125 (
            .O(N__9705),
            .I(N__9702));
    LocalMux I__2124 (
            .O(N__9702),
            .I(N__9699));
    Span12Mux_v I__2123 (
            .O(N__9699),
            .I(N__9696));
    Odrv12 I__2122 (
            .O(N__9696),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2121 (
            .O(N__9693),
            .I(N__9690));
    LocalMux I__2120 (
            .O(N__9690),
            .I(N__9687));
    Odrv4 I__2119 (
            .O(N__9687),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__2118 (
            .O(N__9684),
            .I(N__9681));
    LocalMux I__2117 (
            .O(N__9681),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2116 (
            .O(N__9678),
            .I(N__9675));
    LocalMux I__2115 (
            .O(N__9675),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__2114 (
            .O(N__9672),
            .I(bfn_13_12_0_));
    InMux I__2113 (
            .O(N__9669),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__2112 (
            .O(N__9666),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__2111 (
            .O(N__9663),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__2110 (
            .O(N__9660),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__2109 (
            .O(N__9657),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__2108 (
            .O(N__9654),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__2107 (
            .O(N__9651),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__2106 (
            .O(N__9648),
            .I(N__9645));
    LocalMux I__2105 (
            .O(N__9645),
            .I(N__9641));
    InMux I__2104 (
            .O(N__9644),
            .I(N__9638));
    Span4Mux_h I__2103 (
            .O(N__9641),
            .I(N__9635));
    LocalMux I__2102 (
            .O(N__9638),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__2101 (
            .O(N__9635),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__2100 (
            .O(N__9630),
            .I(N__9606));
    ClkMux I__2099 (
            .O(N__9629),
            .I(N__9606));
    ClkMux I__2098 (
            .O(N__9628),
            .I(N__9606));
    ClkMux I__2097 (
            .O(N__9627),
            .I(N__9606));
    ClkMux I__2096 (
            .O(N__9626),
            .I(N__9606));
    ClkMux I__2095 (
            .O(N__9625),
            .I(N__9606));
    ClkMux I__2094 (
            .O(N__9624),
            .I(N__9606));
    ClkMux I__2093 (
            .O(N__9623),
            .I(N__9606));
    GlobalMux I__2092 (
            .O(N__9606),
            .I(N__9603));
    gio2CtrlBuf I__2091 (
            .O(N__9603),
            .I(C1_c_g));
    SRMux I__2090 (
            .O(N__9600),
            .I(N__9597));
    LocalMux I__2089 (
            .O(N__9597),
            .I(N__9594));
    Span4Mux_h I__2088 (
            .O(N__9594),
            .I(N__9591));
    Odrv4 I__2087 (
            .O(N__9591),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__2086 (
            .O(N__9588),
            .I(N__9584));
    InMux I__2085 (
            .O(N__9587),
            .I(N__9581));
    LocalMux I__2084 (
            .O(N__9584),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__2083 (
            .O(N__9581),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__2082 (
            .O(N__9576),
            .I(N__9572));
    InMux I__2081 (
            .O(N__9575),
            .I(N__9569));
    LocalMux I__2080 (
            .O(N__9572),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__2079 (
            .O(N__9569),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__2078 (
            .O(N__9564),
            .I(N__9560));
    InMux I__2077 (
            .O(N__9563),
            .I(N__9557));
    InMux I__2076 (
            .O(N__9560),
            .I(N__9554));
    LocalMux I__2075 (
            .O(N__9557),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__2074 (
            .O(N__9554),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__2073 (
            .O(N__9549),
            .I(N__9545));
    InMux I__2072 (
            .O(N__9548),
            .I(N__9542));
    LocalMux I__2071 (
            .O(N__9545),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__2070 (
            .O(N__9542),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__2069 (
            .O(N__9537),
            .I(N__9534));
    LocalMux I__2068 (
            .O(N__9534),
            .I(\U712_REG_SM.N_351 ));
    CascadeMux I__2067 (
            .O(N__9531),
            .I(N__9528));
    InMux I__2066 (
            .O(N__9528),
            .I(N__9525));
    LocalMux I__2065 (
            .O(N__9525),
            .I(N__9522));
    Span4Mux_h I__2064 (
            .O(N__9522),
            .I(N__9518));
    InMux I__2063 (
            .O(N__9521),
            .I(N__9515));
    Odrv4 I__2062 (
            .O(N__9518),
            .I(\U712_REG_SM.N_435 ));
    LocalMux I__2061 (
            .O(N__9515),
            .I(\U712_REG_SM.N_435 ));
    InMux I__2060 (
            .O(N__9510),
            .I(N__9507));
    LocalMux I__2059 (
            .O(N__9507),
            .I(N__9503));
    InMux I__2058 (
            .O(N__9506),
            .I(N__9497));
    Span4Mux_h I__2057 (
            .O(N__9503),
            .I(N__9494));
    InMux I__2056 (
            .O(N__9502),
            .I(N__9491));
    InMux I__2055 (
            .O(N__9501),
            .I(N__9486));
    InMux I__2054 (
            .O(N__9500),
            .I(N__9486));
    LocalMux I__2053 (
            .O(N__9497),
            .I(\U712_REG_SM.N_345 ));
    Odrv4 I__2052 (
            .O(N__9494),
            .I(\U712_REG_SM.N_345 ));
    LocalMux I__2051 (
            .O(N__9491),
            .I(\U712_REG_SM.N_345 ));
    LocalMux I__2050 (
            .O(N__9486),
            .I(\U712_REG_SM.N_345 ));
    InMux I__2049 (
            .O(N__9477),
            .I(N__9474));
    LocalMux I__2048 (
            .O(N__9474),
            .I(N__9469));
    InMux I__2047 (
            .O(N__9473),
            .I(N__9465));
    InMux I__2046 (
            .O(N__9472),
            .I(N__9462));
    Span4Mux_h I__2045 (
            .O(N__9469),
            .I(N__9459));
    InMux I__2044 (
            .O(N__9468),
            .I(N__9456));
    LocalMux I__2043 (
            .O(N__9465),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__2042 (
            .O(N__9462),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    Odrv4 I__2041 (
            .O(N__9459),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__2040 (
            .O(N__9456),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__2039 (
            .O(N__9447),
            .I(N__9440));
    CascadeMux I__2038 (
            .O(N__9446),
            .I(N__9437));
    InMux I__2037 (
            .O(N__9445),
            .I(N__9433));
    InMux I__2036 (
            .O(N__9444),
            .I(N__9430));
    CascadeMux I__2035 (
            .O(N__9443),
            .I(N__9427));
    LocalMux I__2034 (
            .O(N__9440),
            .I(N__9424));
    InMux I__2033 (
            .O(N__9437),
            .I(N__9419));
    InMux I__2032 (
            .O(N__9436),
            .I(N__9419));
    LocalMux I__2031 (
            .O(N__9433),
            .I(N__9416));
    LocalMux I__2030 (
            .O(N__9430),
            .I(N__9413));
    InMux I__2029 (
            .O(N__9427),
            .I(N__9406));
    Span4Mux_v I__2028 (
            .O(N__9424),
            .I(N__9403));
    LocalMux I__2027 (
            .O(N__9419),
            .I(N__9396));
    Span4Mux_h I__2026 (
            .O(N__9416),
            .I(N__9396));
    Span4Mux_h I__2025 (
            .O(N__9413),
            .I(N__9396));
    InMux I__2024 (
            .O(N__9412),
            .I(N__9391));
    InMux I__2023 (
            .O(N__9411),
            .I(N__9391));
    InMux I__2022 (
            .O(N__9410),
            .I(N__9386));
    InMux I__2021 (
            .O(N__9409),
            .I(N__9386));
    LocalMux I__2020 (
            .O(N__9406),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2019 (
            .O(N__9403),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2018 (
            .O(N__9396),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2017 (
            .O(N__9391),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2016 (
            .O(N__9386),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__2015 (
            .O(N__9375),
            .I(N__9372));
    LocalMux I__2014 (
            .O(N__9372),
            .I(N__9369));
    Span4Mux_s1_v I__2013 (
            .O(N__9369),
            .I(N__9366));
    Sp12to4 I__2012 (
            .O(N__9366),
            .I(N__9363));
    Span12Mux_h I__2011 (
            .O(N__9363),
            .I(N__9360));
    Odrv12 I__2010 (
            .O(N__9360),
            .I(ASn_c));
    CEMux I__2009 (
            .O(N__9357),
            .I(N__9354));
    LocalMux I__2008 (
            .O(N__9354),
            .I(N__9351));
    Odrv4 I__2007 (
            .O(N__9351),
            .I(\U712_REG_SM.N_131_0 ));
    IoInMux I__2006 (
            .O(N__9348),
            .I(N__9345));
    LocalMux I__2005 (
            .O(N__9345),
            .I(N__9342));
    Odrv12 I__2004 (
            .O(N__9342),
            .I(RESETn_c_i));
    InMux I__2003 (
            .O(N__9339),
            .I(N__9333));
    InMux I__2002 (
            .O(N__9338),
            .I(N__9333));
    LocalMux I__2001 (
            .O(N__9333),
            .I(N__9330));
    Span4Mux_h I__2000 (
            .O(N__9330),
            .I(N__9327));
    Odrv4 I__1999 (
            .O(N__9327),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1998 (
            .O(N__9324),
            .I(N__9321));
    LocalMux I__1997 (
            .O(N__9321),
            .I(N__9318));
    Odrv4 I__1996 (
            .O(N__9318),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1995 (
            .O(N__9315),
            .I(N__9311));
    InMux I__1994 (
            .O(N__9314),
            .I(N__9308));
    LocalMux I__1993 (
            .O(N__9311),
            .I(N__9305));
    LocalMux I__1992 (
            .O(N__9308),
            .I(N__9302));
    Span4Mux_h I__1991 (
            .O(N__9305),
            .I(N__9295));
    Span4Mux_v I__1990 (
            .O(N__9302),
            .I(N__9295));
    InMux I__1989 (
            .O(N__9301),
            .I(N__9290));
    InMux I__1988 (
            .O(N__9300),
            .I(N__9290));
    Span4Mux_h I__1987 (
            .O(N__9295),
            .I(N__9287));
    LocalMux I__1986 (
            .O(N__9290),
            .I(N__9284));
    Sp12to4 I__1985 (
            .O(N__9287),
            .I(N__9281));
    Span12Mux_h I__1984 (
            .O(N__9284),
            .I(N__9278));
    Odrv12 I__1983 (
            .O(N__9281),
            .I(DRA_c_8));
    Odrv12 I__1982 (
            .O(N__9278),
            .I(DRA_c_8));
    InMux I__1981 (
            .O(N__9273),
            .I(N__9268));
    InMux I__1980 (
            .O(N__9272),
            .I(N__9265));
    InMux I__1979 (
            .O(N__9271),
            .I(N__9262));
    LocalMux I__1978 (
            .O(N__9268),
            .I(N__9259));
    LocalMux I__1977 (
            .O(N__9265),
            .I(N__9254));
    LocalMux I__1976 (
            .O(N__9262),
            .I(N__9254));
    Span4Mux_v I__1975 (
            .O(N__9259),
            .I(N__9250));
    Span4Mux_v I__1974 (
            .O(N__9254),
            .I(N__9247));
    InMux I__1973 (
            .O(N__9253),
            .I(N__9244));
    Sp12to4 I__1972 (
            .O(N__9250),
            .I(N__9237));
    Sp12to4 I__1971 (
            .O(N__9247),
            .I(N__9237));
    LocalMux I__1970 (
            .O(N__9244),
            .I(N__9237));
    Span12Mux_h I__1969 (
            .O(N__9237),
            .I(N__9234));
    Odrv12 I__1968 (
            .O(N__9234),
            .I(DRA_c_7));
    InMux I__1967 (
            .O(N__9231),
            .I(N__9228));
    LocalMux I__1966 (
            .O(N__9228),
            .I(N__9225));
    Odrv4 I__1965 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1964 (
            .O(N__9222),
            .I(N__9218));
    InMux I__1963 (
            .O(N__9221),
            .I(N__9215));
    LocalMux I__1962 (
            .O(N__9218),
            .I(N__9212));
    LocalMux I__1961 (
            .O(N__9215),
            .I(N__9209));
    Span4Mux_v I__1960 (
            .O(N__9212),
            .I(N__9204));
    Span4Mux_v I__1959 (
            .O(N__9209),
            .I(N__9204));
    Sp12to4 I__1958 (
            .O(N__9204),
            .I(N__9201));
    Span12Mux_h I__1957 (
            .O(N__9201),
            .I(N__9198));
    Span12Mux_v I__1956 (
            .O(N__9198),
            .I(N__9195));
    Odrv12 I__1955 (
            .O(N__9195),
            .I(DRA_c_0));
    InMux I__1954 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__1953 (
            .O(N__9189),
            .I(N__9184));
    InMux I__1952 (
            .O(N__9188),
            .I(N__9181));
    InMux I__1951 (
            .O(N__9187),
            .I(N__9178));
    Span4Mux_v I__1950 (
            .O(N__9184),
            .I(N__9175));
    LocalMux I__1949 (
            .O(N__9181),
            .I(N__9172));
    LocalMux I__1948 (
            .O(N__9178),
            .I(N__9169));
    Span4Mux_v I__1947 (
            .O(N__9175),
            .I(N__9165));
    Span4Mux_v I__1946 (
            .O(N__9172),
            .I(N__9160));
    Span4Mux_h I__1945 (
            .O(N__9169),
            .I(N__9160));
    InMux I__1944 (
            .O(N__9168),
            .I(N__9157));
    Span4Mux_v I__1943 (
            .O(N__9165),
            .I(N__9154));
    Span4Mux_h I__1942 (
            .O(N__9160),
            .I(N__9149));
    LocalMux I__1941 (
            .O(N__9157),
            .I(N__9149));
    Span4Mux_v I__1940 (
            .O(N__9154),
            .I(N__9146));
    Sp12to4 I__1939 (
            .O(N__9149),
            .I(N__9143));
    Sp12to4 I__1938 (
            .O(N__9146),
            .I(N__9138));
    Span12Mux_v I__1937 (
            .O(N__9143),
            .I(N__9138));
    Span12Mux_h I__1936 (
            .O(N__9138),
            .I(N__9135));
    Odrv12 I__1935 (
            .O(N__9135),
            .I(DRA_c_1));
    InMux I__1934 (
            .O(N__9132),
            .I(N__9129));
    LocalMux I__1933 (
            .O(N__9129),
            .I(N__9126));
    Odrv12 I__1932 (
            .O(N__9126),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1931 (
            .O(N__9123),
            .I(N__9120));
    LocalMux I__1930 (
            .O(N__9120),
            .I(N__9117));
    Span4Mux_h I__1929 (
            .O(N__9117),
            .I(N__9114));
    Odrv4 I__1928 (
            .O(N__9114),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1927 (
            .O(N__9111),
            .I(N__9105));
    InMux I__1926 (
            .O(N__9110),
            .I(N__9105));
    LocalMux I__1925 (
            .O(N__9105),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__1924 (
            .O(N__9102),
            .I(N__9098));
    InMux I__1923 (
            .O(N__9101),
            .I(N__9095));
    LocalMux I__1922 (
            .O(N__9098),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    LocalMux I__1921 (
            .O(N__9095),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    CascadeMux I__1920 (
            .O(N__9090),
            .I(N__9086));
    InMux I__1919 (
            .O(N__9089),
            .I(N__9083));
    InMux I__1918 (
            .O(N__9086),
            .I(N__9080));
    LocalMux I__1917 (
            .O(N__9083),
            .I(DBR_SYNC_i_1));
    LocalMux I__1916 (
            .O(N__9080),
            .I(DBR_SYNC_i_1));
    InMux I__1915 (
            .O(N__9075),
            .I(N__9072));
    LocalMux I__1914 (
            .O(N__9072),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    InMux I__1913 (
            .O(N__9069),
            .I(N__9065));
    InMux I__1912 (
            .O(N__9068),
            .I(N__9062));
    LocalMux I__1911 (
            .O(N__9065),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ));
    LocalMux I__1910 (
            .O(N__9062),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ));
    CascadeMux I__1909 (
            .O(N__9057),
            .I(N__9054));
    InMux I__1908 (
            .O(N__9054),
            .I(N__9051));
    LocalMux I__1907 (
            .O(N__9051),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    InMux I__1906 (
            .O(N__9048),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    InMux I__1905 (
            .O(N__9045),
            .I(N__9041));
    InMux I__1904 (
            .O(N__9044),
            .I(N__9038));
    LocalMux I__1903 (
            .O(N__9041),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    LocalMux I__1902 (
            .O(N__9038),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    CascadeMux I__1901 (
            .O(N__9033),
            .I(N__9030));
    InMux I__1900 (
            .O(N__9030),
            .I(N__9027));
    LocalMux I__1899 (
            .O(N__9027),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    InMux I__1898 (
            .O(N__9024),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__1897 (
            .O(N__9021),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    InMux I__1896 (
            .O(N__9018),
            .I(N__9015));
    LocalMux I__1895 (
            .O(N__9015),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__1894 (
            .O(N__9012),
            .I(N__9007));
    InMux I__1893 (
            .O(N__9011),
            .I(N__8997));
    InMux I__1892 (
            .O(N__9010),
            .I(N__8997));
    InMux I__1891 (
            .O(N__9007),
            .I(N__8997));
    InMux I__1890 (
            .O(N__9006),
            .I(N__8994));
    InMux I__1889 (
            .O(N__9005),
            .I(N__8991));
    InMux I__1888 (
            .O(N__9004),
            .I(N__8988));
    LocalMux I__1887 (
            .O(N__8997),
            .I(N__8985));
    LocalMux I__1886 (
            .O(N__8994),
            .I(N__8980));
    LocalMux I__1885 (
            .O(N__8991),
            .I(N__8975));
    LocalMux I__1884 (
            .O(N__8988),
            .I(N__8975));
    Span4Mux_h I__1883 (
            .O(N__8985),
            .I(N__8971));
    InMux I__1882 (
            .O(N__8984),
            .I(N__8968));
    InMux I__1881 (
            .O(N__8983),
            .I(N__8965));
    Span4Mux_h I__1880 (
            .O(N__8980),
            .I(N__8960));
    Span4Mux_v I__1879 (
            .O(N__8975),
            .I(N__8960));
    InMux I__1878 (
            .O(N__8974),
            .I(N__8957));
    Odrv4 I__1877 (
            .O(N__8971),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1876 (
            .O(N__8968),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1875 (
            .O(N__8965),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1874 (
            .O(N__8960),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1873 (
            .O(N__8957),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1872 (
            .O(N__8946),
            .I(N__8942));
    CascadeMux I__1871 (
            .O(N__8945),
            .I(N__8938));
    LocalMux I__1870 (
            .O(N__8942),
            .I(N__8935));
    CascadeMux I__1869 (
            .O(N__8941),
            .I(N__8928));
    InMux I__1868 (
            .O(N__8938),
            .I(N__8925));
    Span4Mux_h I__1867 (
            .O(N__8935),
            .I(N__8922));
    InMux I__1866 (
            .O(N__8934),
            .I(N__8913));
    InMux I__1865 (
            .O(N__8933),
            .I(N__8913));
    InMux I__1864 (
            .O(N__8932),
            .I(N__8913));
    InMux I__1863 (
            .O(N__8931),
            .I(N__8913));
    InMux I__1862 (
            .O(N__8928),
            .I(N__8910));
    LocalMux I__1861 (
            .O(N__8925),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__1860 (
            .O(N__8922),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1859 (
            .O(N__8913),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1858 (
            .O(N__8910),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1857 (
            .O(N__8901),
            .I(N__8898));
    LocalMux I__1856 (
            .O(N__8898),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ));
    InMux I__1855 (
            .O(N__8895),
            .I(N__8892));
    LocalMux I__1854 (
            .O(N__8892),
            .I(N__8889));
    Span4Mux_h I__1853 (
            .O(N__8889),
            .I(N__8885));
    InMux I__1852 (
            .O(N__8888),
            .I(N__8882));
    Odrv4 I__1851 (
            .O(N__8885),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    LocalMux I__1850 (
            .O(N__8882),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__1849 (
            .O(N__8877),
            .I(N__8874));
    LocalMux I__1848 (
            .O(N__8874),
            .I(N__8871));
    Odrv4 I__1847 (
            .O(N__8871),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1846 (
            .O(N__8868),
            .I(N__8865));
    LocalMux I__1845 (
            .O(N__8865),
            .I(N__8862));
    Odrv4 I__1844 (
            .O(N__8862),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1843 (
            .O(N__8859),
            .I(N__8856));
    LocalMux I__1842 (
            .O(N__8856),
            .I(N__8853));
    Odrv12 I__1841 (
            .O(N__8853),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1840 (
            .O(N__8850),
            .I(N__8847));
    LocalMux I__1839 (
            .O(N__8847),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ));
    InMux I__1838 (
            .O(N__8844),
            .I(N__8841));
    LocalMux I__1837 (
            .O(N__8841),
            .I(N__8837));
    CascadeMux I__1836 (
            .O(N__8840),
            .I(N__8834));
    Span4Mux_v I__1835 (
            .O(N__8837),
            .I(N__8831));
    InMux I__1834 (
            .O(N__8834),
            .I(N__8828));
    Span4Mux_h I__1833 (
            .O(N__8831),
            .I(N__8823));
    LocalMux I__1832 (
            .O(N__8828),
            .I(N__8823));
    Span4Mux_v I__1831 (
            .O(N__8823),
            .I(N__8818));
    InMux I__1830 (
            .O(N__8822),
            .I(N__8815));
    InMux I__1829 (
            .O(N__8821),
            .I(N__8812));
    Odrv4 I__1828 (
            .O(N__8818),
            .I(REG_CYCLEm));
    LocalMux I__1827 (
            .O(N__8815),
            .I(REG_CYCLEm));
    LocalMux I__1826 (
            .O(N__8812),
            .I(REG_CYCLEm));
    IoInMux I__1825 (
            .O(N__8805),
            .I(N__8802));
    LocalMux I__1824 (
            .O(N__8802),
            .I(N__8799));
    Span4Mux_s2_v I__1823 (
            .O(N__8799),
            .I(N__8796));
    Span4Mux_h I__1822 (
            .O(N__8796),
            .I(N__8793));
    Span4Mux_v I__1821 (
            .O(N__8793),
            .I(N__8790));
    Sp12to4 I__1820 (
            .O(N__8790),
            .I(N__8787));
    Span12Mux_h I__1819 (
            .O(N__8787),
            .I(N__8784));
    Odrv12 I__1818 (
            .O(N__8784),
            .I(N_196_i));
    InMux I__1817 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__1816 (
            .O(N__8778),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    InMux I__1815 (
            .O(N__8775),
            .I(N__8772));
    LocalMux I__1814 (
            .O(N__8772),
            .I(N__8769));
    Span4Mux_h I__1813 (
            .O(N__8769),
            .I(N__8766));
    Odrv4 I__1812 (
            .O(N__8766),
            .I(\U712_CHIP_RAM.N_492 ));
    InMux I__1811 (
            .O(N__8763),
            .I(N__8758));
    InMux I__1810 (
            .O(N__8762),
            .I(N__8755));
    InMux I__1809 (
            .O(N__8761),
            .I(N__8752));
    LocalMux I__1808 (
            .O(N__8758),
            .I(\U712_REG_SM.N_131 ));
    LocalMux I__1807 (
            .O(N__8755),
            .I(\U712_REG_SM.N_131 ));
    LocalMux I__1806 (
            .O(N__8752),
            .I(\U712_REG_SM.N_131 ));
    InMux I__1805 (
            .O(N__8745),
            .I(N__8742));
    LocalMux I__1804 (
            .O(N__8742),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_7 ));
    InMux I__1803 (
            .O(N__8739),
            .I(N__8736));
    LocalMux I__1802 (
            .O(N__8736),
            .I(N__8732));
    InMux I__1801 (
            .O(N__8735),
            .I(N__8729));
    Odrv4 I__1800 (
            .O(N__8732),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_5 ));
    LocalMux I__1799 (
            .O(N__8729),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_5 ));
    InMux I__1798 (
            .O(N__8724),
            .I(N__8721));
    LocalMux I__1797 (
            .O(N__8721),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_6 ));
    InMux I__1796 (
            .O(N__8718),
            .I(N__8715));
    LocalMux I__1795 (
            .O(N__8715),
            .I(N__8709));
    InMux I__1794 (
            .O(N__8714),
            .I(N__8706));
    InMux I__1793 (
            .O(N__8713),
            .I(N__8703));
    CascadeMux I__1792 (
            .O(N__8712),
            .I(N__8700));
    Span4Mux_v I__1791 (
            .O(N__8709),
            .I(N__8694));
    LocalMux I__1790 (
            .O(N__8706),
            .I(N__8694));
    LocalMux I__1789 (
            .O(N__8703),
            .I(N__8691));
    InMux I__1788 (
            .O(N__8700),
            .I(N__8688));
    InMux I__1787 (
            .O(N__8699),
            .I(N__8685));
    Span4Mux_h I__1786 (
            .O(N__8694),
            .I(N__8680));
    Span4Mux_h I__1785 (
            .O(N__8691),
            .I(N__8680));
    LocalMux I__1784 (
            .O(N__8688),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1783 (
            .O(N__8685),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1782 (
            .O(N__8680),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1781 (
            .O(N__8673),
            .I(N__8670));
    LocalMux I__1780 (
            .O(N__8670),
            .I(N__8667));
    Span4Mux_s3_v I__1779 (
            .O(N__8667),
            .I(N__8664));
    Span4Mux_v I__1778 (
            .O(N__8664),
            .I(N__8661));
    Sp12to4 I__1777 (
            .O(N__8661),
            .I(N__8658));
    Span12Mux_h I__1776 (
            .O(N__8658),
            .I(N__8655));
    Odrv12 I__1775 (
            .O(N__8655),
            .I(CRCSn_c));
    InMux I__1774 (
            .O(N__8652),
            .I(N__8649));
    LocalMux I__1773 (
            .O(N__8649),
            .I(N__8646));
    Span4Mux_h I__1772 (
            .O(N__8646),
            .I(N__8643));
    Odrv4 I__1771 (
            .O(N__8643),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1770 (
            .O(N__8640),
            .I(N__8637));
    LocalMux I__1769 (
            .O(N__8637),
            .I(N__8634));
    Span4Mux_v I__1768 (
            .O(N__8634),
            .I(N__8631));
    Odrv4 I__1767 (
            .O(N__8631),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1766 (
            .O(N__8628),
            .I(N__8625));
    LocalMux I__1765 (
            .O(N__8625),
            .I(N__8622));
    Odrv4 I__1764 (
            .O(N__8622),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1763 (
            .O(N__8619),
            .I(N__8616));
    LocalMux I__1762 (
            .O(N__8616),
            .I(N__8613));
    Span4Mux_h I__1761 (
            .O(N__8613),
            .I(N__8610));
    Odrv4 I__1760 (
            .O(N__8610),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1759 (
            .O(N__8607),
            .I(N__8604));
    LocalMux I__1758 (
            .O(N__8604),
            .I(N__8601));
    Span4Mux_h I__1757 (
            .O(N__8601),
            .I(N__8598));
    Odrv4 I__1756 (
            .O(N__8598),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1755 (
            .O(N__8595),
            .I(N__8592));
    LocalMux I__1754 (
            .O(N__8592),
            .I(N__8586));
    InMux I__1753 (
            .O(N__8591),
            .I(N__8583));
    InMux I__1752 (
            .O(N__8590),
            .I(N__8580));
    InMux I__1751 (
            .O(N__8589),
            .I(N__8577));
    Odrv4 I__1750 (
            .O(N__8586),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__1749 (
            .O(N__8583),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__1748 (
            .O(N__8580),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__1747 (
            .O(N__8577),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__1746 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1745 (
            .O(N__8565),
            .I(\U712_REG_SM.N_365 ));
    InMux I__1744 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__1743 (
            .O(N__8559),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_4 ));
    InMux I__1742 (
            .O(N__8556),
            .I(N__8553));
    LocalMux I__1741 (
            .O(N__8553),
            .I(\U712_REG_SM.N_588 ));
    InMux I__1740 (
            .O(N__8550),
            .I(N__8547));
    LocalMux I__1739 (
            .O(N__8547),
            .I(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ));
    InMux I__1738 (
            .O(N__8544),
            .I(N__8540));
    InMux I__1737 (
            .O(N__8543),
            .I(N__8537));
    LocalMux I__1736 (
            .O(N__8540),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1735 (
            .O(N__8537),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__1734 (
            .O(N__8532),
            .I(N__8529));
    InMux I__1733 (
            .O(N__8529),
            .I(N__8526));
    LocalMux I__1732 (
            .O(N__8526),
            .I(N__8521));
    InMux I__1731 (
            .O(N__8525),
            .I(N__8518));
    InMux I__1730 (
            .O(N__8524),
            .I(N__8510));
    Span4Mux_h I__1729 (
            .O(N__8521),
            .I(N__8505));
    LocalMux I__1728 (
            .O(N__8518),
            .I(N__8505));
    InMux I__1727 (
            .O(N__8517),
            .I(N__8498));
    InMux I__1726 (
            .O(N__8516),
            .I(N__8498));
    InMux I__1725 (
            .O(N__8515),
            .I(N__8498));
    InMux I__1724 (
            .O(N__8514),
            .I(N__8493));
    InMux I__1723 (
            .O(N__8513),
            .I(N__8493));
    LocalMux I__1722 (
            .O(N__8510),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1721 (
            .O(N__8505),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1720 (
            .O(N__8498),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1719 (
            .O(N__8493),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1718 (
            .O(N__8484),
            .I(N__8480));
    InMux I__1717 (
            .O(N__8483),
            .I(N__8476));
    InMux I__1716 (
            .O(N__8480),
            .I(N__8471));
    InMux I__1715 (
            .O(N__8479),
            .I(N__8468));
    LocalMux I__1714 (
            .O(N__8476),
            .I(N__8465));
    InMux I__1713 (
            .O(N__8475),
            .I(N__8460));
    InMux I__1712 (
            .O(N__8474),
            .I(N__8460));
    LocalMux I__1711 (
            .O(N__8471),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1710 (
            .O(N__8468),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    Odrv4 I__1709 (
            .O(N__8465),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1708 (
            .O(N__8460),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    CascadeMux I__1707 (
            .O(N__8451),
            .I(\U712_REG_SM.N_395_cascade_ ));
    CascadeMux I__1706 (
            .O(N__8448),
            .I(\U712_REG_SM.N_439_cascade_ ));
    InMux I__1705 (
            .O(N__8445),
            .I(N__8442));
    LocalMux I__1704 (
            .O(N__8442),
            .I(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ));
    InMux I__1703 (
            .O(N__8439),
            .I(N__8436));
    LocalMux I__1702 (
            .O(N__8436),
            .I(\U712_REG_SM.N_395 ));
    CascadeMux I__1701 (
            .O(N__8433),
            .I(N__8430));
    InMux I__1700 (
            .O(N__8430),
            .I(N__8424));
    InMux I__1699 (
            .O(N__8429),
            .I(N__8419));
    InMux I__1698 (
            .O(N__8428),
            .I(N__8419));
    InMux I__1697 (
            .O(N__8427),
            .I(N__8416));
    LocalMux I__1696 (
            .O(N__8424),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1695 (
            .O(N__8419),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1694 (
            .O(N__8416),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    IoInMux I__1693 (
            .O(N__8409),
            .I(N__8406));
    LocalMux I__1692 (
            .O(N__8406),
            .I(N__8403));
    Span4Mux_s2_v I__1691 (
            .O(N__8403),
            .I(N__8400));
    Span4Mux_v I__1690 (
            .O(N__8400),
            .I(N__8396));
    InMux I__1689 (
            .O(N__8399),
            .I(N__8393));
    Span4Mux_h I__1688 (
            .O(N__8396),
            .I(N__8390));
    LocalMux I__1687 (
            .O(N__8393),
            .I(N__8387));
    Odrv4 I__1686 (
            .O(N__8390),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1685 (
            .O(N__8387),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1684 (
            .O(N__8382),
            .I(N__8375));
    InMux I__1683 (
            .O(N__8381),
            .I(N__8370));
    InMux I__1682 (
            .O(N__8380),
            .I(N__8370));
    CascadeMux I__1681 (
            .O(N__8379),
            .I(N__8366));
    CascadeMux I__1680 (
            .O(N__8378),
            .I(N__8361));
    InMux I__1679 (
            .O(N__8375),
            .I(N__8354));
    LocalMux I__1678 (
            .O(N__8370),
            .I(N__8351));
    InMux I__1677 (
            .O(N__8369),
            .I(N__8346));
    InMux I__1676 (
            .O(N__8366),
            .I(N__8346));
    InMux I__1675 (
            .O(N__8365),
            .I(N__8343));
    InMux I__1674 (
            .O(N__8364),
            .I(N__8330));
    InMux I__1673 (
            .O(N__8361),
            .I(N__8325));
    InMux I__1672 (
            .O(N__8360),
            .I(N__8325));
    InMux I__1671 (
            .O(N__8359),
            .I(N__8318));
    InMux I__1670 (
            .O(N__8358),
            .I(N__8318));
    InMux I__1669 (
            .O(N__8357),
            .I(N__8318));
    LocalMux I__1668 (
            .O(N__8354),
            .I(N__8311));
    Span4Mux_h I__1667 (
            .O(N__8351),
            .I(N__8311));
    LocalMux I__1666 (
            .O(N__8346),
            .I(N__8311));
    LocalMux I__1665 (
            .O(N__8343),
            .I(N__8308));
    InMux I__1664 (
            .O(N__8342),
            .I(N__8301));
    InMux I__1663 (
            .O(N__8341),
            .I(N__8301));
    InMux I__1662 (
            .O(N__8340),
            .I(N__8301));
    InMux I__1661 (
            .O(N__8339),
            .I(N__8296));
    InMux I__1660 (
            .O(N__8338),
            .I(N__8296));
    InMux I__1659 (
            .O(N__8337),
            .I(N__8293));
    InMux I__1658 (
            .O(N__8336),
            .I(N__8290));
    InMux I__1657 (
            .O(N__8335),
            .I(N__8287));
    InMux I__1656 (
            .O(N__8334),
            .I(N__8282));
    InMux I__1655 (
            .O(N__8333),
            .I(N__8282));
    LocalMux I__1654 (
            .O(N__8330),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1653 (
            .O(N__8325),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1652 (
            .O(N__8318),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1651 (
            .O(N__8311),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1650 (
            .O(N__8308),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1649 (
            .O(N__8301),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1648 (
            .O(N__8296),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1647 (
            .O(N__8293),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1646 (
            .O(N__8290),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1645 (
            .O(N__8287),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1644 (
            .O(N__8282),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1643 (
            .O(N__8259),
            .I(N__8256));
    LocalMux I__1642 (
            .O(N__8256),
            .I(N__8253));
    Odrv12 I__1641 (
            .O(N__8253),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    IoInMux I__1640 (
            .O(N__8250),
            .I(N__8247));
    LocalMux I__1639 (
            .O(N__8247),
            .I(N__8244));
    Span4Mux_s2_v I__1638 (
            .O(N__8244),
            .I(N__8241));
    Sp12to4 I__1637 (
            .O(N__8241),
            .I(N__8238));
    Span12Mux_h I__1636 (
            .O(N__8238),
            .I(N__8235));
    Span12Mux_v I__1635 (
            .O(N__8235),
            .I(N__8231));
    InMux I__1634 (
            .O(N__8234),
            .I(N__8228));
    Odrv12 I__1633 (
            .O(N__8231),
            .I(PRnW_c));
    LocalMux I__1632 (
            .O(N__8228),
            .I(PRnW_c));
    InMux I__1631 (
            .O(N__8223),
            .I(N__8220));
    LocalMux I__1630 (
            .O(N__8220),
            .I(N__8215));
    InMux I__1629 (
            .O(N__8219),
            .I(N__8212));
    InMux I__1628 (
            .O(N__8218),
            .I(N__8209));
    Odrv4 I__1627 (
            .O(N__8215),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1626 (
            .O(N__8212),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1625 (
            .O(N__8209),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__1624 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1623 (
            .O(N__8199),
            .I(N__8194));
    InMux I__1622 (
            .O(N__8198),
            .I(N__8189));
    InMux I__1621 (
            .O(N__8197),
            .I(N__8186));
    Span4Mux_h I__1620 (
            .O(N__8194),
            .I(N__8183));
    InMux I__1619 (
            .O(N__8193),
            .I(N__8178));
    InMux I__1618 (
            .O(N__8192),
            .I(N__8178));
    LocalMux I__1617 (
            .O(N__8189),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1616 (
            .O(N__8186),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__1615 (
            .O(N__8183),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1614 (
            .O(N__8178),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__1613 (
            .O(N__8169),
            .I(\U712_REG_SM.N_351_cascade_ ));
    InMux I__1612 (
            .O(N__8166),
            .I(N__8162));
    InMux I__1611 (
            .O(N__8165),
            .I(N__8159));
    LocalMux I__1610 (
            .O(N__8162),
            .I(N__8156));
    LocalMux I__1609 (
            .O(N__8159),
            .I(\U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ));
    Odrv4 I__1608 (
            .O(N__8156),
            .I(\U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ));
    InMux I__1607 (
            .O(N__8151),
            .I(N__8142));
    InMux I__1606 (
            .O(N__8150),
            .I(N__8142));
    InMux I__1605 (
            .O(N__8149),
            .I(N__8142));
    LocalMux I__1604 (
            .O(N__8142),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1603 (
            .O(N__8139),
            .I(N__8135));
    InMux I__1602 (
            .O(N__8138),
            .I(N__8132));
    LocalMux I__1601 (
            .O(N__8135),
            .I(N__8127));
    LocalMux I__1600 (
            .O(N__8132),
            .I(N__8127));
    Span12Mux_h I__1599 (
            .O(N__8127),
            .I(N__8124));
    Span12Mux_v I__1598 (
            .O(N__8124),
            .I(N__8121));
    Odrv12 I__1597 (
            .O(N__8121),
            .I(TSn_c));
    InMux I__1596 (
            .O(N__8118),
            .I(N__8115));
    LocalMux I__1595 (
            .O(N__8115),
            .I(N__8111));
    IoInMux I__1594 (
            .O(N__8114),
            .I(N__8108));
    Span12Mux_h I__1593 (
            .O(N__8111),
            .I(N__8105));
    LocalMux I__1592 (
            .O(N__8108),
            .I(N__8102));
    Span12Mux_v I__1591 (
            .O(N__8105),
            .I(N__8099));
    IoSpan4Mux I__1590 (
            .O(N__8102),
            .I(N__8096));
    Odrv12 I__1589 (
            .O(N__8099),
            .I(RAMENn_c));
    Odrv4 I__1588 (
            .O(N__8096),
            .I(RAMENn_c));
    CascadeMux I__1587 (
            .O(N__8091),
            .I(\U712_CHIP_RAM.N_448_cascade_ ));
    InMux I__1586 (
            .O(N__8088),
            .I(N__8083));
    InMux I__1585 (
            .O(N__8087),
            .I(N__8078));
    InMux I__1584 (
            .O(N__8086),
            .I(N__8078));
    LocalMux I__1583 (
            .O(N__8083),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1582 (
            .O(N__8078),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__1581 (
            .O(N__8073),
            .I(N__8070));
    LocalMux I__1580 (
            .O(N__8070),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    CascadeMux I__1579 (
            .O(N__8067),
            .I(N__8064));
    InMux I__1578 (
            .O(N__8064),
            .I(N__8061));
    LocalMux I__1577 (
            .O(N__8061),
            .I(\U712_CHIP_RAM.N_450 ));
    InMux I__1576 (
            .O(N__8058),
            .I(N__8055));
    LocalMux I__1575 (
            .O(N__8055),
            .I(N__8052));
    Sp12to4 I__1574 (
            .O(N__8052),
            .I(N__8049));
    Span12Mux_v I__1573 (
            .O(N__8049),
            .I(N__8046));
    Span12Mux_h I__1572 (
            .O(N__8046),
            .I(N__8043));
    Odrv12 I__1571 (
            .O(N__8043),
            .I(A_c_15));
    InMux I__1570 (
            .O(N__8040),
            .I(N__8037));
    LocalMux I__1569 (
            .O(N__8037),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    CascadeMux I__1568 (
            .O(N__8034),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1567 (
            .O(N__8031),
            .I(N__8028));
    LocalMux I__1566 (
            .O(N__8028),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    InMux I__1565 (
            .O(N__8025),
            .I(N__8022));
    LocalMux I__1564 (
            .O(N__8022),
            .I(N__8019));
    Sp12to4 I__1563 (
            .O(N__8019),
            .I(N__8016));
    Span12Mux_v I__1562 (
            .O(N__8016),
            .I(N__8013));
    Span12Mux_h I__1561 (
            .O(N__8013),
            .I(N__8010));
    Odrv12 I__1560 (
            .O(N__8010),
            .I(A_c_13));
    CascadeMux I__1559 (
            .O(N__8007),
            .I(N__8004));
    InMux I__1558 (
            .O(N__8004),
            .I(N__7995));
    InMux I__1557 (
            .O(N__8003),
            .I(N__7990));
    InMux I__1556 (
            .O(N__8002),
            .I(N__7990));
    InMux I__1555 (
            .O(N__8001),
            .I(N__7986));
    InMux I__1554 (
            .O(N__8000),
            .I(N__7974));
    InMux I__1553 (
            .O(N__7999),
            .I(N__7974));
    InMux I__1552 (
            .O(N__7998),
            .I(N__7974));
    LocalMux I__1551 (
            .O(N__7995),
            .I(N__7969));
    LocalMux I__1550 (
            .O(N__7990),
            .I(N__7969));
    CascadeMux I__1549 (
            .O(N__7989),
            .I(N__7960));
    LocalMux I__1548 (
            .O(N__7986),
            .I(N__7950));
    InMux I__1547 (
            .O(N__7985),
            .I(N__7947));
    InMux I__1546 (
            .O(N__7984),
            .I(N__7942));
    InMux I__1545 (
            .O(N__7983),
            .I(N__7942));
    InMux I__1544 (
            .O(N__7982),
            .I(N__7939));
    InMux I__1543 (
            .O(N__7981),
            .I(N__7936));
    LocalMux I__1542 (
            .O(N__7974),
            .I(N__7931));
    Span4Mux_v I__1541 (
            .O(N__7969),
            .I(N__7931));
    InMux I__1540 (
            .O(N__7968),
            .I(N__7926));
    InMux I__1539 (
            .O(N__7967),
            .I(N__7926));
    InMux I__1538 (
            .O(N__7966),
            .I(N__7921));
    InMux I__1537 (
            .O(N__7965),
            .I(N__7921));
    InMux I__1536 (
            .O(N__7964),
            .I(N__7910));
    InMux I__1535 (
            .O(N__7963),
            .I(N__7910));
    InMux I__1534 (
            .O(N__7960),
            .I(N__7910));
    InMux I__1533 (
            .O(N__7959),
            .I(N__7910));
    InMux I__1532 (
            .O(N__7958),
            .I(N__7910));
    InMux I__1531 (
            .O(N__7957),
            .I(N__7899));
    InMux I__1530 (
            .O(N__7956),
            .I(N__7899));
    InMux I__1529 (
            .O(N__7955),
            .I(N__7899));
    InMux I__1528 (
            .O(N__7954),
            .I(N__7899));
    InMux I__1527 (
            .O(N__7953),
            .I(N__7899));
    Span4Mux_v I__1526 (
            .O(N__7950),
            .I(N__7892));
    LocalMux I__1525 (
            .O(N__7947),
            .I(N__7892));
    LocalMux I__1524 (
            .O(N__7942),
            .I(N__7892));
    LocalMux I__1523 (
            .O(N__7939),
            .I(N__7889));
    LocalMux I__1522 (
            .O(N__7936),
            .I(N__7884));
    Span4Mux_v I__1521 (
            .O(N__7931),
            .I(N__7884));
    LocalMux I__1520 (
            .O(N__7926),
            .I(N__7879));
    LocalMux I__1519 (
            .O(N__7921),
            .I(N__7879));
    LocalMux I__1518 (
            .O(N__7910),
            .I(N__7874));
    LocalMux I__1517 (
            .O(N__7899),
            .I(N__7874));
    Odrv4 I__1516 (
            .O(N__7892),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1515 (
            .O(N__7889),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1514 (
            .O(N__7884),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1513 (
            .O(N__7879),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1512 (
            .O(N__7874),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1511 (
            .O(N__7863),
            .I(N__7860));
    LocalMux I__1510 (
            .O(N__7860),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1509 (
            .O(N__7857),
            .I(N__7854));
    LocalMux I__1508 (
            .O(N__7854),
            .I(N__7851));
    Span4Mux_v I__1507 (
            .O(N__7851),
            .I(N__7848));
    Sp12to4 I__1506 (
            .O(N__7848),
            .I(N__7845));
    Span12Mux_h I__1505 (
            .O(N__7845),
            .I(N__7842));
    Odrv12 I__1504 (
            .O(N__7842),
            .I(A_c_6));
    InMux I__1503 (
            .O(N__7839),
            .I(N__7836));
    LocalMux I__1502 (
            .O(N__7836),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CEMux I__1501 (
            .O(N__7833),
            .I(N__7830));
    LocalMux I__1500 (
            .O(N__7830),
            .I(N__7826));
    CEMux I__1499 (
            .O(N__7829),
            .I(N__7823));
    Span4Mux_v I__1498 (
            .O(N__7826),
            .I(N__7820));
    LocalMux I__1497 (
            .O(N__7823),
            .I(N__7817));
    Odrv4 I__1496 (
            .O(N__7820),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv12 I__1495 (
            .O(N__7817),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    InMux I__1494 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__1493 (
            .O(N__7809),
            .I(N__7806));
    Span4Mux_h I__1492 (
            .O(N__7806),
            .I(N__7803));
    Span4Mux_v I__1491 (
            .O(N__7803),
            .I(N__7800));
    Sp12to4 I__1490 (
            .O(N__7800),
            .I(N__7797));
    Span12Mux_h I__1489 (
            .O(N__7797),
            .I(N__7794));
    Odrv12 I__1488 (
            .O(N__7794),
            .I(A_c_20));
    InMux I__1487 (
            .O(N__7791),
            .I(N__7786));
    InMux I__1486 (
            .O(N__7790),
            .I(N__7781));
    InMux I__1485 (
            .O(N__7789),
            .I(N__7781));
    LocalMux I__1484 (
            .O(N__7786),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1483 (
            .O(N__7781),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    InMux I__1482 (
            .O(N__7776),
            .I(N__7773));
    LocalMux I__1481 (
            .O(N__7773),
            .I(N__7769));
    InMux I__1480 (
            .O(N__7772),
            .I(N__7766));
    Span4Mux_h I__1479 (
            .O(N__7769),
            .I(N__7763));
    LocalMux I__1478 (
            .O(N__7766),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__1477 (
            .O(N__7763),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__1476 (
            .O(N__7758),
            .I(N__7754));
    InMux I__1475 (
            .O(N__7757),
            .I(N__7751));
    LocalMux I__1474 (
            .O(N__7754),
            .I(N__7748));
    LocalMux I__1473 (
            .O(N__7751),
            .I(N__7745));
    Span4Mux_h I__1472 (
            .O(N__7748),
            .I(N__7742));
    Odrv12 I__1471 (
            .O(N__7745),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ));
    Odrv4 I__1470 (
            .O(N__7742),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ));
    InMux I__1469 (
            .O(N__7737),
            .I(N__7733));
    InMux I__1468 (
            .O(N__7736),
            .I(N__7730));
    LocalMux I__1467 (
            .O(N__7733),
            .I(N__7724));
    LocalMux I__1466 (
            .O(N__7730),
            .I(N__7724));
    InMux I__1465 (
            .O(N__7729),
            .I(N__7719));
    Span4Mux_h I__1464 (
            .O(N__7724),
            .I(N__7716));
    InMux I__1463 (
            .O(N__7723),
            .I(N__7713));
    InMux I__1462 (
            .O(N__7722),
            .I(N__7710));
    LocalMux I__1461 (
            .O(N__7719),
            .I(\U712_CHIP_RAM.N_510 ));
    Odrv4 I__1460 (
            .O(N__7716),
            .I(\U712_CHIP_RAM.N_510 ));
    LocalMux I__1459 (
            .O(N__7713),
            .I(\U712_CHIP_RAM.N_510 ));
    LocalMux I__1458 (
            .O(N__7710),
            .I(\U712_CHIP_RAM.N_510 ));
    InMux I__1457 (
            .O(N__7701),
            .I(N__7698));
    LocalMux I__1456 (
            .O(N__7698),
            .I(N__7695));
    Span4Mux_h I__1455 (
            .O(N__7695),
            .I(N__7691));
    InMux I__1454 (
            .O(N__7694),
            .I(N__7688));
    Odrv4 I__1453 (
            .O(N__7691),
            .I(\U712_CHIP_RAM.N_461 ));
    LocalMux I__1452 (
            .O(N__7688),
            .I(\U712_CHIP_RAM.N_461 ));
    CascadeMux I__1451 (
            .O(N__7683),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ));
    IoInMux I__1450 (
            .O(N__7680),
            .I(N__7677));
    LocalMux I__1449 (
            .O(N__7677),
            .I(N__7674));
    Span4Mux_s3_v I__1448 (
            .O(N__7674),
            .I(N__7671));
    Sp12to4 I__1447 (
            .O(N__7671),
            .I(N__7668));
    Span12Mux_h I__1446 (
            .O(N__7668),
            .I(N__7664));
    InMux I__1445 (
            .O(N__7667),
            .I(N__7661));
    Odrv12 I__1444 (
            .O(N__7664),
            .I(LATCH_CLK_c));
    LocalMux I__1443 (
            .O(N__7661),
            .I(LATCH_CLK_c));
    InMux I__1442 (
            .O(N__7656),
            .I(N__7653));
    LocalMux I__1441 (
            .O(N__7653),
            .I(\U712_REG_SM.N_357 ));
    CascadeMux I__1440 (
            .O(N__7650),
            .I(N__7646));
    InMux I__1439 (
            .O(N__7649),
            .I(N__7643));
    InMux I__1438 (
            .O(N__7646),
            .I(N__7640));
    LocalMux I__1437 (
            .O(N__7643),
            .I(\U712_REG_SM.N_353 ));
    LocalMux I__1436 (
            .O(N__7640),
            .I(\U712_REG_SM.N_353 ));
    IoInMux I__1435 (
            .O(N__7635),
            .I(N__7632));
    LocalMux I__1434 (
            .O(N__7632),
            .I(N__7629));
    Span4Mux_s1_v I__1433 (
            .O(N__7629),
            .I(N__7626));
    Sp12to4 I__1432 (
            .O(N__7626),
            .I(N__7623));
    Span12Mux_h I__1431 (
            .O(N__7623),
            .I(N__7620));
    Odrv12 I__1430 (
            .O(N__7620),
            .I(CASn_c));
    InMux I__1429 (
            .O(N__7617),
            .I(N__7613));
    CascadeMux I__1428 (
            .O(N__7616),
            .I(N__7607));
    LocalMux I__1427 (
            .O(N__7613),
            .I(N__7604));
    InMux I__1426 (
            .O(N__7612),
            .I(N__7601));
    InMux I__1425 (
            .O(N__7611),
            .I(N__7598));
    InMux I__1424 (
            .O(N__7610),
            .I(N__7593));
    InMux I__1423 (
            .O(N__7607),
            .I(N__7593));
    Span4Mux_v I__1422 (
            .O(N__7604),
            .I(N__7583));
    LocalMux I__1421 (
            .O(N__7601),
            .I(N__7583));
    LocalMux I__1420 (
            .O(N__7598),
            .I(N__7583));
    LocalMux I__1419 (
            .O(N__7593),
            .I(N__7583));
    InMux I__1418 (
            .O(N__7592),
            .I(N__7580));
    Span4Mux_h I__1417 (
            .O(N__7583),
            .I(N__7577));
    LocalMux I__1416 (
            .O(N__7580),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1415 (
            .O(N__7577),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1414 (
            .O(N__7572),
            .I(N__7569));
    LocalMux I__1413 (
            .O(N__7569),
            .I(N__7566));
    Span4Mux_s2_v I__1412 (
            .O(N__7566),
            .I(N__7563));
    Span4Mux_h I__1411 (
            .O(N__7563),
            .I(N__7560));
    Sp12to4 I__1410 (
            .O(N__7560),
            .I(N__7557));
    Span12Mux_v I__1409 (
            .O(N__7557),
            .I(N__7554));
    Odrv12 I__1408 (
            .O(N__7554),
            .I(RASn_c));
    CascadeMux I__1407 (
            .O(N__7551),
            .I(N__7548));
    InMux I__1406 (
            .O(N__7548),
            .I(N__7545));
    LocalMux I__1405 (
            .O(N__7545),
            .I(N__7541));
    InMux I__1404 (
            .O(N__7544),
            .I(N__7538));
    Span4Mux_h I__1403 (
            .O(N__7541),
            .I(N__7535));
    LocalMux I__1402 (
            .O(N__7538),
            .I(N__7532));
    Span4Mux_v I__1401 (
            .O(N__7535),
            .I(N__7527));
    Span4Mux_v I__1400 (
            .O(N__7532),
            .I(N__7527));
    Odrv4 I__1399 (
            .O(N__7527),
            .I(DBRn_c_i));
    InMux I__1398 (
            .O(N__7524),
            .I(N__7520));
    InMux I__1397 (
            .O(N__7523),
            .I(N__7517));
    LocalMux I__1396 (
            .O(N__7520),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    LocalMux I__1395 (
            .O(N__7517),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1394 (
            .O(N__7512),
            .I(N__7509));
    LocalMux I__1393 (
            .O(N__7509),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1392 (
            .O(N__7506),
            .I(N__7503));
    LocalMux I__1391 (
            .O(N__7503),
            .I(N__7500));
    Span4Mux_h I__1390 (
            .O(N__7500),
            .I(N__7497));
    Odrv4 I__1389 (
            .O(N__7497),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    IoInMux I__1388 (
            .O(N__7494),
            .I(N__7491));
    LocalMux I__1387 (
            .O(N__7491),
            .I(N__7488));
    IoSpan4Mux I__1386 (
            .O(N__7488),
            .I(N__7485));
    IoSpan4Mux I__1385 (
            .O(N__7485),
            .I(N__7482));
    Span4Mux_s3_h I__1384 (
            .O(N__7482),
            .I(N__7479));
    Span4Mux_h I__1383 (
            .O(N__7479),
            .I(N__7476));
    Sp12to4 I__1382 (
            .O(N__7476),
            .I(N__7472));
    InMux I__1381 (
            .O(N__7475),
            .I(N__7469));
    Span12Mux_h I__1380 (
            .O(N__7472),
            .I(N__7464));
    LocalMux I__1379 (
            .O(N__7469),
            .I(N__7464));
    Span12Mux_h I__1378 (
            .O(N__7464),
            .I(N__7461));
    Odrv12 I__1377 (
            .O(N__7461),
            .I(C3_c));
    IoInMux I__1376 (
            .O(N__7458),
            .I(N__7455));
    LocalMux I__1375 (
            .O(N__7455),
            .I(N__7451));
    IoInMux I__1374 (
            .O(N__7454),
            .I(N__7448));
    IoSpan4Mux I__1373 (
            .O(N__7451),
            .I(N__7445));
    LocalMux I__1372 (
            .O(N__7448),
            .I(N__7442));
    Span4Mux_s1_v I__1371 (
            .O(N__7445),
            .I(N__7439));
    Span4Mux_s1_v I__1370 (
            .O(N__7442),
            .I(N__7436));
    Span4Mux_v I__1369 (
            .O(N__7439),
            .I(N__7433));
    Span4Mux_v I__1368 (
            .O(N__7436),
            .I(N__7430));
    Sp12to4 I__1367 (
            .O(N__7433),
            .I(N__7427));
    Sp12to4 I__1366 (
            .O(N__7430),
            .I(N__7424));
    Span12Mux_h I__1365 (
            .O(N__7427),
            .I(N__7418));
    Span12Mux_h I__1364 (
            .O(N__7424),
            .I(N__7418));
    InMux I__1363 (
            .O(N__7423),
            .I(N__7415));
    Odrv12 I__1362 (
            .O(N__7418),
            .I(BLSn_c));
    LocalMux I__1361 (
            .O(N__7415),
            .I(BLSn_c));
    InMux I__1360 (
            .O(N__7410),
            .I(N__7407));
    LocalMux I__1359 (
            .O(N__7407),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__1358 (
            .O(N__7404),
            .I(\U712_REG_SM.N_345_cascade_ ));
    InMux I__1357 (
            .O(N__7401),
            .I(N__7396));
    InMux I__1356 (
            .O(N__7400),
            .I(N__7391));
    InMux I__1355 (
            .O(N__7399),
            .I(N__7391));
    LocalMux I__1354 (
            .O(N__7396),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1353 (
            .O(N__7391),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    InMux I__1352 (
            .O(N__7386),
            .I(N__7383));
    LocalMux I__1351 (
            .O(N__7383),
            .I(\U712_REG_SM.N_396 ));
    CascadeMux I__1350 (
            .O(N__7380),
            .I(\U712_REG_SM.N_435_cascade_ ));
    InMux I__1349 (
            .O(N__7377),
            .I(N__7371));
    InMux I__1348 (
            .O(N__7376),
            .I(N__7371));
    LocalMux I__1347 (
            .O(N__7371),
            .I(\U712_REG_SM.N_352 ));
    InMux I__1346 (
            .O(N__7368),
            .I(N__7362));
    InMux I__1345 (
            .O(N__7367),
            .I(N__7362));
    LocalMux I__1344 (
            .O(N__7362),
            .I(\U712_CHIP_RAM.N_500 ));
    CascadeMux I__1343 (
            .O(N__7359),
            .I(N__7350));
    InMux I__1342 (
            .O(N__7358),
            .I(N__7346));
    InMux I__1341 (
            .O(N__7357),
            .I(N__7343));
    InMux I__1340 (
            .O(N__7356),
            .I(N__7340));
    InMux I__1339 (
            .O(N__7355),
            .I(N__7337));
    InMux I__1338 (
            .O(N__7354),
            .I(N__7334));
    InMux I__1337 (
            .O(N__7353),
            .I(N__7331));
    InMux I__1336 (
            .O(N__7350),
            .I(N__7326));
    InMux I__1335 (
            .O(N__7349),
            .I(N__7326));
    LocalMux I__1334 (
            .O(N__7346),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1333 (
            .O(N__7343),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1332 (
            .O(N__7340),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1331 (
            .O(N__7337),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1330 (
            .O(N__7334),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1329 (
            .O(N__7331),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1328 (
            .O(N__7326),
            .I(\U712_CHIP_RAM.N_503 ));
    CascadeMux I__1327 (
            .O(N__7311),
            .I(\U712_CHIP_RAM.N_500_cascade_ ));
    InMux I__1326 (
            .O(N__7308),
            .I(N__7305));
    LocalMux I__1325 (
            .O(N__7305),
            .I(N__7300));
    InMux I__1324 (
            .O(N__7304),
            .I(N__7293));
    InMux I__1323 (
            .O(N__7303),
            .I(N__7293));
    Span4Mux_h I__1322 (
            .O(N__7300),
            .I(N__7290));
    InMux I__1321 (
            .O(N__7299),
            .I(N__7287));
    InMux I__1320 (
            .O(N__7298),
            .I(N__7284));
    LocalMux I__1319 (
            .O(N__7293),
            .I(\U712_CHIP_RAM.N_514 ));
    Odrv4 I__1318 (
            .O(N__7290),
            .I(\U712_CHIP_RAM.N_514 ));
    LocalMux I__1317 (
            .O(N__7287),
            .I(\U712_CHIP_RAM.N_514 ));
    LocalMux I__1316 (
            .O(N__7284),
            .I(\U712_CHIP_RAM.N_514 ));
    InMux I__1315 (
            .O(N__7275),
            .I(N__7270));
    InMux I__1314 (
            .O(N__7274),
            .I(N__7267));
    InMux I__1313 (
            .O(N__7273),
            .I(N__7264));
    LocalMux I__1312 (
            .O(N__7270),
            .I(N__7261));
    LocalMux I__1311 (
            .O(N__7267),
            .I(N__7256));
    LocalMux I__1310 (
            .O(N__7264),
            .I(N__7246));
    Span4Mux_h I__1309 (
            .O(N__7261),
            .I(N__7246));
    InMux I__1308 (
            .O(N__7260),
            .I(N__7241));
    InMux I__1307 (
            .O(N__7259),
            .I(N__7241));
    Span4Mux_h I__1306 (
            .O(N__7256),
            .I(N__7238));
    InMux I__1305 (
            .O(N__7255),
            .I(N__7233));
    InMux I__1304 (
            .O(N__7254),
            .I(N__7233));
    InMux I__1303 (
            .O(N__7253),
            .I(N__7226));
    InMux I__1302 (
            .O(N__7252),
            .I(N__7226));
    InMux I__1301 (
            .O(N__7251),
            .I(N__7226));
    Odrv4 I__1300 (
            .O(N__7246),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1299 (
            .O(N__7241),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1298 (
            .O(N__7238),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1297 (
            .O(N__7233),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1296 (
            .O(N__7226),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1295 (
            .O(N__7215),
            .I(N__7211));
    InMux I__1294 (
            .O(N__7214),
            .I(N__7208));
    LocalMux I__1293 (
            .O(N__7211),
            .I(N__7203));
    LocalMux I__1292 (
            .O(N__7208),
            .I(N__7203));
    Odrv4 I__1291 (
            .O(N__7203),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    InMux I__1290 (
            .O(N__7200),
            .I(N__7197));
    LocalMux I__1289 (
            .O(N__7197),
            .I(N__7194));
    Span4Mux_h I__1288 (
            .O(N__7194),
            .I(N__7190));
    InMux I__1287 (
            .O(N__7193),
            .I(N__7187));
    Odrv4 I__1286 (
            .O(N__7190),
            .I(\U712_CHIP_RAM.N_337 ));
    LocalMux I__1285 (
            .O(N__7187),
            .I(\U712_CHIP_RAM.N_337 ));
    InMux I__1284 (
            .O(N__7182),
            .I(N__7179));
    LocalMux I__1283 (
            .O(N__7179),
            .I(N__7176));
    Odrv4 I__1282 (
            .O(N__7176),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1 ));
    InMux I__1281 (
            .O(N__7173),
            .I(N__7168));
    CascadeMux I__1280 (
            .O(N__7172),
            .I(N__7165));
    InMux I__1279 (
            .O(N__7171),
            .I(N__7160));
    LocalMux I__1278 (
            .O(N__7168),
            .I(N__7154));
    InMux I__1277 (
            .O(N__7165),
            .I(N__7151));
    InMux I__1276 (
            .O(N__7164),
            .I(N__7148));
    CascadeMux I__1275 (
            .O(N__7163),
            .I(N__7145));
    LocalMux I__1274 (
            .O(N__7160),
            .I(N__7142));
    InMux I__1273 (
            .O(N__7159),
            .I(N__7139));
    CascadeMux I__1272 (
            .O(N__7158),
            .I(N__7135));
    CascadeMux I__1271 (
            .O(N__7157),
            .I(N__7131));
    Span4Mux_h I__1270 (
            .O(N__7154),
            .I(N__7125));
    LocalMux I__1269 (
            .O(N__7151),
            .I(N__7125));
    LocalMux I__1268 (
            .O(N__7148),
            .I(N__7120));
    InMux I__1267 (
            .O(N__7145),
            .I(N__7117));
    Span4Mux_h I__1266 (
            .O(N__7142),
            .I(N__7112));
    LocalMux I__1265 (
            .O(N__7139),
            .I(N__7112));
    InMux I__1264 (
            .O(N__7138),
            .I(N__7109));
    InMux I__1263 (
            .O(N__7135),
            .I(N__7106));
    InMux I__1262 (
            .O(N__7134),
            .I(N__7101));
    InMux I__1261 (
            .O(N__7131),
            .I(N__7101));
    InMux I__1260 (
            .O(N__7130),
            .I(N__7098));
    Span4Mux_h I__1259 (
            .O(N__7125),
            .I(N__7095));
    InMux I__1258 (
            .O(N__7124),
            .I(N__7090));
    InMux I__1257 (
            .O(N__7123),
            .I(N__7090));
    Span4Mux_h I__1256 (
            .O(N__7120),
            .I(N__7087));
    LocalMux I__1255 (
            .O(N__7117),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1254 (
            .O(N__7112),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1253 (
            .O(N__7109),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1252 (
            .O(N__7106),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1251 (
            .O(N__7101),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1250 (
            .O(N__7098),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1249 (
            .O(N__7095),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1248 (
            .O(N__7090),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1247 (
            .O(N__7087),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1246 (
            .O(N__7068),
            .I(N__7062));
    InMux I__1245 (
            .O(N__7067),
            .I(N__7059));
    CascadeMux I__1244 (
            .O(N__7066),
            .I(N__7055));
    InMux I__1243 (
            .O(N__7065),
            .I(N__7050));
    InMux I__1242 (
            .O(N__7062),
            .I(N__7050));
    LocalMux I__1241 (
            .O(N__7059),
            .I(N__7046));
    CascadeMux I__1240 (
            .O(N__7058),
            .I(N__7043));
    InMux I__1239 (
            .O(N__7055),
            .I(N__7039));
    LocalMux I__1238 (
            .O(N__7050),
            .I(N__7036));
    CascadeMux I__1237 (
            .O(N__7049),
            .I(N__7031));
    Span4Mux_v I__1236 (
            .O(N__7046),
            .I(N__7026));
    InMux I__1235 (
            .O(N__7043),
            .I(N__7023));
    InMux I__1234 (
            .O(N__7042),
            .I(N__7020));
    LocalMux I__1233 (
            .O(N__7039),
            .I(N__7015));
    Span4Mux_h I__1232 (
            .O(N__7036),
            .I(N__7015));
    InMux I__1231 (
            .O(N__7035),
            .I(N__7012));
    InMux I__1230 (
            .O(N__7034),
            .I(N__7009));
    InMux I__1229 (
            .O(N__7031),
            .I(N__7004));
    InMux I__1228 (
            .O(N__7030),
            .I(N__7004));
    InMux I__1227 (
            .O(N__7029),
            .I(N__7001));
    Odrv4 I__1226 (
            .O(N__7026),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1225 (
            .O(N__7023),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1224 (
            .O(N__7020),
            .I(\U712_CHIP_RAM.N_332 ));
    Odrv4 I__1223 (
            .O(N__7015),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1222 (
            .O(N__7012),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1221 (
            .O(N__7009),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1220 (
            .O(N__7004),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__1219 (
            .O(N__7001),
            .I(\U712_CHIP_RAM.N_332 ));
    InMux I__1218 (
            .O(N__6984),
            .I(N__6978));
    InMux I__1217 (
            .O(N__6983),
            .I(N__6978));
    LocalMux I__1216 (
            .O(N__6978),
            .I(CPU_TACKm));
    CEMux I__1215 (
            .O(N__6975),
            .I(N__6972));
    LocalMux I__1214 (
            .O(N__6972),
            .I(N__6969));
    Odrv4 I__1213 (
            .O(N__6969),
            .I(\U712_CHIP_RAM.N_248_0 ));
    InMux I__1212 (
            .O(N__6966),
            .I(N__6962));
    InMux I__1211 (
            .O(N__6965),
            .I(N__6959));
    LocalMux I__1210 (
            .O(N__6962),
            .I(N__6953));
    LocalMux I__1209 (
            .O(N__6959),
            .I(N__6953));
    InMux I__1208 (
            .O(N__6958),
            .I(N__6949));
    Span4Mux_v I__1207 (
            .O(N__6953),
            .I(N__6946));
    InMux I__1206 (
            .O(N__6952),
            .I(N__6943));
    LocalMux I__1205 (
            .O(N__6949),
            .I(N__6939));
    Span4Mux_v I__1204 (
            .O(N__6946),
            .I(N__6934));
    LocalMux I__1203 (
            .O(N__6943),
            .I(N__6934));
    CascadeMux I__1202 (
            .O(N__6942),
            .I(N__6931));
    Span4Mux_v I__1201 (
            .O(N__6939),
            .I(N__6926));
    Span4Mux_v I__1200 (
            .O(N__6934),
            .I(N__6926));
    InMux I__1199 (
            .O(N__6931),
            .I(N__6923));
    Sp12to4 I__1198 (
            .O(N__6926),
            .I(N__6918));
    LocalMux I__1197 (
            .O(N__6923),
            .I(N__6918));
    Span12Mux_h I__1196 (
            .O(N__6918),
            .I(N__6915));
    Odrv12 I__1195 (
            .O(N__6915),
            .I(RnW_c));
    InMux I__1194 (
            .O(N__6912),
            .I(N__6909));
    LocalMux I__1193 (
            .O(N__6909),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__1192 (
            .O(N__6906),
            .I(N__6903));
    InMux I__1191 (
            .O(N__6903),
            .I(N__6898));
    InMux I__1190 (
            .O(N__6902),
            .I(N__6893));
    InMux I__1189 (
            .O(N__6901),
            .I(N__6893));
    LocalMux I__1188 (
            .O(N__6898),
            .I(REG_TACK));
    LocalMux I__1187 (
            .O(N__6893),
            .I(REG_TACK));
    InMux I__1186 (
            .O(N__6888),
            .I(N__6884));
    InMux I__1185 (
            .O(N__6887),
            .I(N__6881));
    LocalMux I__1184 (
            .O(N__6884),
            .I(N__6878));
    LocalMux I__1183 (
            .O(N__6881),
            .I(\U712_REG_SM.START_RSTZ0 ));
    Odrv4 I__1182 (
            .O(N__6878),
            .I(\U712_REG_SM.START_RSTZ0 ));
    CascadeMux I__1181 (
            .O(N__6873),
            .I(\U712_CHIP_RAM.N_514_cascade_ ));
    InMux I__1180 (
            .O(N__6870),
            .I(N__6866));
    InMux I__1179 (
            .O(N__6869),
            .I(N__6863));
    LocalMux I__1178 (
            .O(N__6866),
            .I(N__6860));
    LocalMux I__1177 (
            .O(N__6863),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ));
    Odrv4 I__1176 (
            .O(N__6860),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ));
    InMux I__1175 (
            .O(N__6855),
            .I(N__6851));
    InMux I__1174 (
            .O(N__6854),
            .I(N__6848));
    LocalMux I__1173 (
            .O(N__6851),
            .I(\U712_CHIP_RAM.N_350 ));
    LocalMux I__1172 (
            .O(N__6848),
            .I(\U712_CHIP_RAM.N_350 ));
    CascadeMux I__1171 (
            .O(N__6843),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ));
    CEMux I__1170 (
            .O(N__6840),
            .I(N__6837));
    LocalMux I__1169 (
            .O(N__6837),
            .I(N__6834));
    Span4Mux_v I__1168 (
            .O(N__6834),
            .I(N__6831));
    Odrv4 I__1167 (
            .O(N__6831),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ));
    InMux I__1166 (
            .O(N__6828),
            .I(N__6825));
    LocalMux I__1165 (
            .O(N__6825),
            .I(N__6820));
    InMux I__1164 (
            .O(N__6824),
            .I(N__6817));
    InMux I__1163 (
            .O(N__6823),
            .I(N__6813));
    Span4Mux_h I__1162 (
            .O(N__6820),
            .I(N__6808));
    LocalMux I__1161 (
            .O(N__6817),
            .I(N__6805));
    InMux I__1160 (
            .O(N__6816),
            .I(N__6802));
    LocalMux I__1159 (
            .O(N__6813),
            .I(N__6799));
    InMux I__1158 (
            .O(N__6812),
            .I(N__6794));
    InMux I__1157 (
            .O(N__6811),
            .I(N__6794));
    Odrv4 I__1156 (
            .O(N__6808),
            .I(\U712_CHIP_RAM.N_501 ));
    Odrv12 I__1155 (
            .O(N__6805),
            .I(\U712_CHIP_RAM.N_501 ));
    LocalMux I__1154 (
            .O(N__6802),
            .I(\U712_CHIP_RAM.N_501 ));
    Odrv4 I__1153 (
            .O(N__6799),
            .I(\U712_CHIP_RAM.N_501 ));
    LocalMux I__1152 (
            .O(N__6794),
            .I(\U712_CHIP_RAM.N_501 ));
    InMux I__1151 (
            .O(N__6783),
            .I(N__6780));
    LocalMux I__1150 (
            .O(N__6780),
            .I(N__6777));
    Odrv4 I__1149 (
            .O(N__6777),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ));
    InMux I__1148 (
            .O(N__6774),
            .I(N__6767));
    InMux I__1147 (
            .O(N__6773),
            .I(N__6767));
    InMux I__1146 (
            .O(N__6772),
            .I(N__6763));
    LocalMux I__1145 (
            .O(N__6767),
            .I(N__6760));
    InMux I__1144 (
            .O(N__6766),
            .I(N__6757));
    LocalMux I__1143 (
            .O(N__6763),
            .I(N__6754));
    Odrv4 I__1142 (
            .O(N__6760),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1141 (
            .O(N__6757),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    Odrv4 I__1140 (
            .O(N__6754),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__1139 (
            .O(N__6747),
            .I(\U712_CHIP_RAM.N_481_cascade_ ));
    CascadeMux I__1138 (
            .O(N__6744),
            .I(\U712_REG_SM.N_428_cascade_ ));
    InMux I__1137 (
            .O(N__6741),
            .I(N__6738));
    LocalMux I__1136 (
            .O(N__6738),
            .I(N__6735));
    Span4Mux_h I__1135 (
            .O(N__6735),
            .I(N__6732));
    Span4Mux_h I__1134 (
            .O(N__6732),
            .I(N__6729));
    Sp12to4 I__1133 (
            .O(N__6729),
            .I(N__6726));
    Span12Mux_v I__1132 (
            .O(N__6726),
            .I(N__6723));
    Odrv12 I__1131 (
            .O(N__6723),
            .I(REGSPACEn_c));
    InMux I__1130 (
            .O(N__6720),
            .I(N__6717));
    LocalMux I__1129 (
            .O(N__6717),
            .I(N__6714));
    Span12Mux_v I__1128 (
            .O(N__6714),
            .I(N__6711));
    Span12Mux_h I__1127 (
            .O(N__6711),
            .I(N__6708));
    Odrv12 I__1126 (
            .O(N__6708),
            .I(A_c_3));
    InMux I__1125 (
            .O(N__6705),
            .I(N__6702));
    LocalMux I__1124 (
            .O(N__6702),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1123 (
            .O(N__6699),
            .I(N__6696));
    LocalMux I__1122 (
            .O(N__6696),
            .I(N__6693));
    Span4Mux_v I__1121 (
            .O(N__6693),
            .I(N__6690));
    Sp12to4 I__1120 (
            .O(N__6690),
            .I(N__6687));
    Span12Mux_h I__1119 (
            .O(N__6687),
            .I(N__6684));
    Odrv12 I__1118 (
            .O(N__6684),
            .I(A_c_4));
    InMux I__1117 (
            .O(N__6681),
            .I(N__6678));
    LocalMux I__1116 (
            .O(N__6678),
            .I(N__6675));
    Span4Mux_h I__1115 (
            .O(N__6675),
            .I(N__6672));
    Odrv4 I__1114 (
            .O(N__6672),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__1113 (
            .O(N__6669),
            .I(N__6666));
    LocalMux I__1112 (
            .O(N__6666),
            .I(N__6663));
    Span4Mux_v I__1111 (
            .O(N__6663),
            .I(N__6660));
    Span4Mux_h I__1110 (
            .O(N__6660),
            .I(N__6657));
    Sp12to4 I__1109 (
            .O(N__6657),
            .I(N__6654));
    Odrv12 I__1108 (
            .O(N__6654),
            .I(A_c_7));
    InMux I__1107 (
            .O(N__6651),
            .I(N__6648));
    LocalMux I__1106 (
            .O(N__6648),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1105 (
            .O(N__6645),
            .I(N__6642));
    LocalMux I__1104 (
            .O(N__6642),
            .I(N__6639));
    Span12Mux_h I__1103 (
            .O(N__6639),
            .I(N__6636));
    Odrv12 I__1102 (
            .O(N__6636),
            .I(A_c_8));
    InMux I__1101 (
            .O(N__6633),
            .I(N__6630));
    LocalMux I__1100 (
            .O(N__6630),
            .I(N__6627));
    Span4Mux_v I__1099 (
            .O(N__6627),
            .I(N__6624));
    Sp12to4 I__1098 (
            .O(N__6624),
            .I(N__6621));
    Span12Mux_h I__1097 (
            .O(N__6621),
            .I(N__6618));
    Odrv12 I__1096 (
            .O(N__6618),
            .I(A_c_5));
    InMux I__1095 (
            .O(N__6615),
            .I(N__6612));
    LocalMux I__1094 (
            .O(N__6612),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__1093 (
            .O(N__6609),
            .I(N__6606));
    LocalMux I__1092 (
            .O(N__6606),
            .I(N__6603));
    Span12Mux_v I__1091 (
            .O(N__6603),
            .I(N__6600));
    Span12Mux_v I__1090 (
            .O(N__6600),
            .I(N__6597));
    Span12Mux_h I__1089 (
            .O(N__6597),
            .I(N__6594));
    Odrv12 I__1088 (
            .O(N__6594),
            .I(A_c_18));
    InMux I__1087 (
            .O(N__6591),
            .I(N__6588));
    LocalMux I__1086 (
            .O(N__6588),
            .I(N__6585));
    Span4Mux_h I__1085 (
            .O(N__6585),
            .I(N__6582));
    Odrv4 I__1084 (
            .O(N__6582),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    CascadeMux I__1083 (
            .O(N__6579),
            .I(N__6576));
    InMux I__1082 (
            .O(N__6576),
            .I(N__6568));
    InMux I__1081 (
            .O(N__6575),
            .I(N__6568));
    InMux I__1080 (
            .O(N__6574),
            .I(N__6565));
    InMux I__1079 (
            .O(N__6573),
            .I(N__6562));
    LocalMux I__1078 (
            .O(N__6568),
            .I(N__6544));
    LocalMux I__1077 (
            .O(N__6565),
            .I(N__6539));
    LocalMux I__1076 (
            .O(N__6562),
            .I(N__6539));
    InMux I__1075 (
            .O(N__6561),
            .I(N__6532));
    InMux I__1074 (
            .O(N__6560),
            .I(N__6532));
    InMux I__1073 (
            .O(N__6559),
            .I(N__6532));
    InMux I__1072 (
            .O(N__6558),
            .I(N__6527));
    InMux I__1071 (
            .O(N__6557),
            .I(N__6527));
    InMux I__1070 (
            .O(N__6556),
            .I(N__6520));
    InMux I__1069 (
            .O(N__6555),
            .I(N__6520));
    InMux I__1068 (
            .O(N__6554),
            .I(N__6520));
    InMux I__1067 (
            .O(N__6553),
            .I(N__6513));
    InMux I__1066 (
            .O(N__6552),
            .I(N__6513));
    InMux I__1065 (
            .O(N__6551),
            .I(N__6513));
    InMux I__1064 (
            .O(N__6550),
            .I(N__6510));
    InMux I__1063 (
            .O(N__6549),
            .I(N__6505));
    InMux I__1062 (
            .O(N__6548),
            .I(N__6505));
    InMux I__1061 (
            .O(N__6547),
            .I(N__6502));
    Span4Mux_h I__1060 (
            .O(N__6544),
            .I(N__6499));
    Odrv4 I__1059 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1058 (
            .O(N__6532),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1057 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1056 (
            .O(N__6520),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1055 (
            .O(N__6513),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1054 (
            .O(N__6510),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1053 (
            .O(N__6505),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1052 (
            .O(N__6502),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1051 (
            .O(N__6499),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1050 (
            .O(N__6480),
            .I(N__6477));
    LocalMux I__1049 (
            .O(N__6477),
            .I(N__6468));
    InMux I__1048 (
            .O(N__6476),
            .I(N__6461));
    InMux I__1047 (
            .O(N__6475),
            .I(N__6456));
    InMux I__1046 (
            .O(N__6474),
            .I(N__6456));
    InMux I__1045 (
            .O(N__6473),
            .I(N__6451));
    InMux I__1044 (
            .O(N__6472),
            .I(N__6448));
    InMux I__1043 (
            .O(N__6471),
            .I(N__6445));
    Span4Mux_h I__1042 (
            .O(N__6468),
            .I(N__6442));
    InMux I__1041 (
            .O(N__6467),
            .I(N__6435));
    InMux I__1040 (
            .O(N__6466),
            .I(N__6435));
    InMux I__1039 (
            .O(N__6465),
            .I(N__6435));
    InMux I__1038 (
            .O(N__6464),
            .I(N__6432));
    LocalMux I__1037 (
            .O(N__6461),
            .I(N__6427));
    LocalMux I__1036 (
            .O(N__6456),
            .I(N__6427));
    InMux I__1035 (
            .O(N__6455),
            .I(N__6422));
    InMux I__1034 (
            .O(N__6454),
            .I(N__6422));
    LocalMux I__1033 (
            .O(N__6451),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1032 (
            .O(N__6448),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1031 (
            .O(N__6445),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1030 (
            .O(N__6442),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1029 (
            .O(N__6435),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1028 (
            .O(N__6432),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1027 (
            .O(N__6427),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1026 (
            .O(N__6422),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1025 (
            .O(N__6405),
            .I(N__6402));
    LocalMux I__1024 (
            .O(N__6402),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__1023 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1022 (
            .O(N__6396),
            .I(N__6393));
    Span4Mux_v I__1021 (
            .O(N__6393),
            .I(N__6390));
    Sp12to4 I__1020 (
            .O(N__6390),
            .I(N__6387));
    Span12Mux_h I__1019 (
            .O(N__6387),
            .I(N__6384));
    Span12Mux_v I__1018 (
            .O(N__6384),
            .I(N__6381));
    Odrv12 I__1017 (
            .O(N__6381),
            .I(A_c_19));
    IoInMux I__1016 (
            .O(N__6378),
            .I(N__6375));
    LocalMux I__1015 (
            .O(N__6375),
            .I(N__6372));
    Span4Mux_s3_h I__1014 (
            .O(N__6372),
            .I(N__6369));
    Sp12to4 I__1013 (
            .O(N__6369),
            .I(N__6366));
    Span12Mux_v I__1012 (
            .O(N__6366),
            .I(N__6363));
    Span12Mux_h I__1011 (
            .O(N__6363),
            .I(N__6360));
    Odrv12 I__1010 (
            .O(N__6360),
            .I(CMA_c_9));
    InMux I__1009 (
            .O(N__6357),
            .I(N__6353));
    InMux I__1008 (
            .O(N__6356),
            .I(N__6350));
    LocalMux I__1007 (
            .O(N__6353),
            .I(N__6342));
    LocalMux I__1006 (
            .O(N__6350),
            .I(N__6339));
    InMux I__1005 (
            .O(N__6349),
            .I(N__6328));
    InMux I__1004 (
            .O(N__6348),
            .I(N__6328));
    InMux I__1003 (
            .O(N__6347),
            .I(N__6328));
    InMux I__1002 (
            .O(N__6346),
            .I(N__6328));
    InMux I__1001 (
            .O(N__6345),
            .I(N__6328));
    Odrv4 I__1000 (
            .O(N__6342),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__999 (
            .O(N__6339),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__998 (
            .O(N__6328),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    CascadeMux I__997 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    CascadeMux I__996 (
            .O(N__6318),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ));
    CEMux I__995 (
            .O(N__6315),
            .I(N__6311));
    CEMux I__994 (
            .O(N__6314),
            .I(N__6308));
    LocalMux I__993 (
            .O(N__6311),
            .I(N__6303));
    LocalMux I__992 (
            .O(N__6308),
            .I(N__6300));
    CEMux I__991 (
            .O(N__6307),
            .I(N__6297));
    CEMux I__990 (
            .O(N__6306),
            .I(N__6294));
    Span4Mux_h I__989 (
            .O(N__6303),
            .I(N__6289));
    Span4Mux_v I__988 (
            .O(N__6300),
            .I(N__6289));
    LocalMux I__987 (
            .O(N__6297),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    LocalMux I__986 (
            .O(N__6294),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__985 (
            .O(N__6289),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    InMux I__984 (
            .O(N__6282),
            .I(N__6279));
    LocalMux I__983 (
            .O(N__6279),
            .I(N__6276));
    Span12Mux_v I__982 (
            .O(N__6276),
            .I(N__6273));
    Span12Mux_h I__981 (
            .O(N__6273),
            .I(N__6270));
    Odrv12 I__980 (
            .O(N__6270),
            .I(A_c_12));
    CascadeMux I__979 (
            .O(N__6267),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__978 (
            .O(N__6264),
            .I(N__6261));
    LocalMux I__977 (
            .O(N__6261),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__976 (
            .O(N__6258),
            .I(N__6255));
    LocalMux I__975 (
            .O(N__6255),
            .I(N__6252));
    Span4Mux_h I__974 (
            .O(N__6252),
            .I(N__6249));
    Sp12to4 I__973 (
            .O(N__6249),
            .I(N__6246));
    Span12Mux_v I__972 (
            .O(N__6246),
            .I(N__6243));
    Odrv12 I__971 (
            .O(N__6243),
            .I(A_c_2));
    InMux I__970 (
            .O(N__6240),
            .I(N__6237));
    LocalMux I__969 (
            .O(N__6237),
            .I(N__6234));
    Span4Mux_h I__968 (
            .O(N__6234),
            .I(N__6231));
    Odrv4 I__967 (
            .O(N__6231),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    InMux I__966 (
            .O(N__6228),
            .I(N__6225));
    LocalMux I__965 (
            .O(N__6225),
            .I(N__6222));
    Span12Mux_v I__964 (
            .O(N__6222),
            .I(N__6219));
    Span12Mux_h I__963 (
            .O(N__6219),
            .I(N__6216));
    Odrv12 I__962 (
            .O(N__6216),
            .I(A_c_16));
    CascadeMux I__961 (
            .O(N__6213),
            .I(N__6210));
    InMux I__960 (
            .O(N__6210),
            .I(N__6207));
    LocalMux I__959 (
            .O(N__6207),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__958 (
            .O(N__6204),
            .I(N__6201));
    LocalMux I__957 (
            .O(N__6201),
            .I(N__6198));
    Span4Mux_v I__956 (
            .O(N__6198),
            .I(N__6195));
    Span4Mux_h I__955 (
            .O(N__6195),
            .I(N__6192));
    Span4Mux_v I__954 (
            .O(N__6192),
            .I(N__6189));
    Span4Mux_v I__953 (
            .O(N__6189),
            .I(N__6186));
    Sp12to4 I__952 (
            .O(N__6186),
            .I(N__6183));
    Odrv12 I__951 (
            .O(N__6183),
            .I(A_c_17));
    CascadeMux I__950 (
            .O(N__6180),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__949 (
            .O(N__6177),
            .I(N__6174));
    LocalMux I__948 (
            .O(N__6174),
            .I(N__6171));
    Span12Mux_v I__947 (
            .O(N__6171),
            .I(N__6168));
    Span12Mux_h I__946 (
            .O(N__6168),
            .I(N__6165));
    Odrv12 I__945 (
            .O(N__6165),
            .I(A_c_14));
    InMux I__944 (
            .O(N__6162),
            .I(N__6159));
    LocalMux I__943 (
            .O(N__6159),
            .I(\U712_CHIP_RAM.N_383 ));
    IoInMux I__942 (
            .O(N__6156),
            .I(N__6153));
    LocalMux I__941 (
            .O(N__6153),
            .I(N__6150));
    IoSpan4Mux I__940 (
            .O(N__6150),
            .I(N__6147));
    Span4Mux_s2_v I__939 (
            .O(N__6147),
            .I(N__6144));
    Sp12to4 I__938 (
            .O(N__6144),
            .I(N__6141));
    Span12Mux_s10_h I__937 (
            .O(N__6141),
            .I(N__6138));
    Span12Mux_v I__936 (
            .O(N__6138),
            .I(N__6135));
    Odrv12 I__935 (
            .O(N__6135),
            .I(CMA_c_3));
    IoInMux I__934 (
            .O(N__6132),
            .I(N__6129));
    LocalMux I__933 (
            .O(N__6129),
            .I(N__6126));
    Span12Mux_s11_h I__932 (
            .O(N__6126),
            .I(N__6123));
    Span12Mux_v I__931 (
            .O(N__6123),
            .I(N__6120));
    Odrv12 I__930 (
            .O(N__6120),
            .I(CMA_c_4));
    IoInMux I__929 (
            .O(N__6117),
            .I(N__6114));
    LocalMux I__928 (
            .O(N__6114),
            .I(N__6111));
    IoSpan4Mux I__927 (
            .O(N__6111),
            .I(N__6108));
    Span4Mux_s2_v I__926 (
            .O(N__6108),
            .I(N__6105));
    Sp12to4 I__925 (
            .O(N__6105),
            .I(N__6102));
    Span12Mux_h I__924 (
            .O(N__6102),
            .I(N__6099));
    Span12Mux_v I__923 (
            .O(N__6099),
            .I(N__6096));
    Odrv12 I__922 (
            .O(N__6096),
            .I(CMA_c_6));
    CascadeMux I__921 (
            .O(N__6093),
            .I(N__6090));
    InMux I__920 (
            .O(N__6090),
            .I(N__6087));
    LocalMux I__919 (
            .O(N__6087),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__918 (
            .O(N__6084),
            .I(N__6081));
    LocalMux I__917 (
            .O(N__6081),
            .I(N__6078));
    Span4Mux_s2_h I__916 (
            .O(N__6078),
            .I(N__6075));
    Span4Mux_h I__915 (
            .O(N__6075),
            .I(N__6072));
    Sp12to4 I__914 (
            .O(N__6072),
            .I(N__6069));
    Span12Mux_v I__913 (
            .O(N__6069),
            .I(N__6066));
    Span12Mux_h I__912 (
            .O(N__6066),
            .I(N__6063));
    Odrv12 I__911 (
            .O(N__6063),
            .I(CMA_c_7));
    CascadeMux I__910 (
            .O(N__6060),
            .I(N__6054));
    CascadeMux I__909 (
            .O(N__6059),
            .I(N__6046));
    CascadeMux I__908 (
            .O(N__6058),
            .I(N__6043));
    CascadeMux I__907 (
            .O(N__6057),
            .I(N__6040));
    InMux I__906 (
            .O(N__6054),
            .I(N__6037));
    InMux I__905 (
            .O(N__6053),
            .I(N__6033));
    InMux I__904 (
            .O(N__6052),
            .I(N__6028));
    InMux I__903 (
            .O(N__6051),
            .I(N__6028));
    InMux I__902 (
            .O(N__6050),
            .I(N__6023));
    InMux I__901 (
            .O(N__6049),
            .I(N__6023));
    InMux I__900 (
            .O(N__6046),
            .I(N__6016));
    InMux I__899 (
            .O(N__6043),
            .I(N__6016));
    InMux I__898 (
            .O(N__6040),
            .I(N__6016));
    LocalMux I__897 (
            .O(N__6037),
            .I(N__6013));
    InMux I__896 (
            .O(N__6036),
            .I(N__6010));
    LocalMux I__895 (
            .O(N__6033),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__894 (
            .O(N__6028),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__893 (
            .O(N__6023),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__892 (
            .O(N__6016),
            .I(\U712_CHIP_RAM.N_343 ));
    Odrv4 I__891 (
            .O(N__6013),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__890 (
            .O(N__6010),
            .I(\U712_CHIP_RAM.N_343 ));
    InMux I__889 (
            .O(N__5997),
            .I(N__5994));
    LocalMux I__888 (
            .O(N__5994),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    IoInMux I__887 (
            .O(N__5991),
            .I(N__5988));
    LocalMux I__886 (
            .O(N__5988),
            .I(N__5985));
    Span4Mux_s2_h I__885 (
            .O(N__5985),
            .I(N__5982));
    Sp12to4 I__884 (
            .O(N__5982),
            .I(N__5979));
    Span12Mux_v I__883 (
            .O(N__5979),
            .I(N__5976));
    Span12Mux_h I__882 (
            .O(N__5976),
            .I(N__5973));
    Odrv12 I__881 (
            .O(N__5973),
            .I(CMA_c_8));
    CascadeMux I__880 (
            .O(N__5970),
            .I(\U712_REG_SM.N_352_cascade_ ));
    IoInMux I__879 (
            .O(N__5967),
            .I(N__5964));
    LocalMux I__878 (
            .O(N__5964),
            .I(N__5960));
    InMux I__877 (
            .O(N__5963),
            .I(N__5957));
    IoSpan4Mux I__876 (
            .O(N__5960),
            .I(N__5954));
    LocalMux I__875 (
            .O(N__5957),
            .I(N__5951));
    IoSpan4Mux I__874 (
            .O(N__5954),
            .I(N__5948));
    Span12Mux_h I__873 (
            .O(N__5951),
            .I(N__5945));
    IoSpan4Mux I__872 (
            .O(N__5948),
            .I(N__5942));
    Odrv12 I__871 (
            .O(N__5945),
            .I(C1_c));
    Odrv4 I__870 (
            .O(N__5942),
            .I(C1_c));
    InMux I__869 (
            .O(N__5937),
            .I(N__5934));
    LocalMux I__868 (
            .O(N__5934),
            .I(N__5931));
    Odrv4 I__867 (
            .O(N__5931),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    IoInMux I__866 (
            .O(N__5928),
            .I(N__5925));
    LocalMux I__865 (
            .O(N__5925),
            .I(N__5922));
    Span4Mux_s2_v I__864 (
            .O(N__5922),
            .I(N__5919));
    Span4Mux_v I__863 (
            .O(N__5919),
            .I(N__5916));
    Sp12to4 I__862 (
            .O(N__5916),
            .I(N__5913));
    Span12Mux_h I__861 (
            .O(N__5913),
            .I(N__5909));
    InMux I__860 (
            .O(N__5912),
            .I(N__5906));
    Odrv12 I__859 (
            .O(N__5909),
            .I(UDSn_c));
    LocalMux I__858 (
            .O(N__5906),
            .I(UDSn_c));
    InMux I__857 (
            .O(N__5901),
            .I(N__5898));
    LocalMux I__856 (
            .O(N__5898),
            .I(\U712_REG_SM.N_429 ));
    IoInMux I__855 (
            .O(N__5895),
            .I(N__5892));
    LocalMux I__854 (
            .O(N__5892),
            .I(N__5889));
    Span4Mux_s3_v I__853 (
            .O(N__5889),
            .I(N__5886));
    Span4Mux_h I__852 (
            .O(N__5886),
            .I(N__5883));
    Sp12to4 I__851 (
            .O(N__5883),
            .I(N__5879));
    CascadeMux I__850 (
            .O(N__5882),
            .I(N__5876));
    Span12Mux_h I__849 (
            .O(N__5879),
            .I(N__5873));
    InMux I__848 (
            .O(N__5876),
            .I(N__5870));
    Odrv12 I__847 (
            .O(N__5873),
            .I(LDSn_c));
    LocalMux I__846 (
            .O(N__5870),
            .I(LDSn_c));
    InMux I__845 (
            .O(N__5865),
            .I(N__5862));
    LocalMux I__844 (
            .O(N__5862),
            .I(\U712_REG_SM.N_493 ));
    InMux I__843 (
            .O(N__5859),
            .I(N__5852));
    InMux I__842 (
            .O(N__5858),
            .I(N__5852));
    InMux I__841 (
            .O(N__5857),
            .I(N__5849));
    LocalMux I__840 (
            .O(N__5852),
            .I(N__5846));
    LocalMux I__839 (
            .O(N__5849),
            .I(N__5843));
    Odrv4 I__838 (
            .O(N__5846),
            .I(\U712_CHIP_RAM.N_590 ));
    Odrv4 I__837 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.N_590 ));
    InMux I__836 (
            .O(N__5838),
            .I(N__5834));
    InMux I__835 (
            .O(N__5837),
            .I(N__5831));
    LocalMux I__834 (
            .O(N__5834),
            .I(\U712_CHIP_RAM.N_476 ));
    LocalMux I__833 (
            .O(N__5831),
            .I(\U712_CHIP_RAM.N_476 ));
    CascadeMux I__832 (
            .O(N__5826),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_ ));
    CascadeMux I__831 (
            .O(N__5823),
            .I(\U712_CHIP_RAM.N_248_cascade_ ));
    InMux I__830 (
            .O(N__5820),
            .I(N__5817));
    LocalMux I__829 (
            .O(N__5817),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__828 (
            .O(N__5814),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__827 (
            .O(N__5811),
            .I(N__5808));
    LocalMux I__826 (
            .O(N__5808),
            .I(N__5805));
    Odrv12 I__825 (
            .O(N__5805),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__824 (
            .O(N__5802),
            .I(N__5799));
    InMux I__823 (
            .O(N__5799),
            .I(N__5793));
    InMux I__822 (
            .O(N__5798),
            .I(N__5793));
    LocalMux I__821 (
            .O(N__5793),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__820 (
            .O(N__5790),
            .I(N__5784));
    InMux I__819 (
            .O(N__5789),
            .I(N__5784));
    LocalMux I__818 (
            .O(N__5784),
            .I(N__5781));
    Odrv12 I__817 (
            .O(N__5781),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__816 (
            .O(N__5778),
            .I(\U712_CYCLE_TERM.N_358_i_cascade_ ));
    IoInMux I__815 (
            .O(N__5775),
            .I(N__5771));
    IoInMux I__814 (
            .O(N__5774),
            .I(N__5767));
    LocalMux I__813 (
            .O(N__5771),
            .I(N__5764));
    IoInMux I__812 (
            .O(N__5770),
            .I(N__5761));
    LocalMux I__811 (
            .O(N__5767),
            .I(N__5758));
    IoSpan4Mux I__810 (
            .O(N__5764),
            .I(N__5755));
    LocalMux I__809 (
            .O(N__5761),
            .I(N__5752));
    Span12Mux_s7_v I__808 (
            .O(N__5758),
            .I(N__5749));
    Sp12to4 I__807 (
            .O(N__5755),
            .I(N__5746));
    IoSpan4Mux I__806 (
            .O(N__5752),
            .I(N__5743));
    Span12Mux_h I__805 (
            .O(N__5749),
            .I(N__5740));
    Span12Mux_s7_v I__804 (
            .O(N__5746),
            .I(N__5737));
    Sp12to4 I__803 (
            .O(N__5743),
            .I(N__5734));
    Span12Mux_v I__802 (
            .O(N__5740),
            .I(N__5728));
    Span12Mux_v I__801 (
            .O(N__5737),
            .I(N__5728));
    Span12Mux_h I__800 (
            .O(N__5734),
            .I(N__5725));
    InMux I__799 (
            .O(N__5733),
            .I(N__5722));
    Odrv12 I__798 (
            .O(N__5728),
            .I(TACK_EN));
    Odrv12 I__797 (
            .O(N__5725),
            .I(TACK_EN));
    LocalMux I__796 (
            .O(N__5722),
            .I(TACK_EN));
    InMux I__795 (
            .O(N__5715),
            .I(N__5707));
    InMux I__794 (
            .O(N__5714),
            .I(N__5707));
    InMux I__793 (
            .O(N__5713),
            .I(N__5704));
    InMux I__792 (
            .O(N__5712),
            .I(N__5701));
    LocalMux I__791 (
            .O(N__5707),
            .I(N__5698));
    LocalMux I__790 (
            .O(N__5704),
            .I(N__5695));
    LocalMux I__789 (
            .O(N__5701),
            .I(N__5692));
    Span4Mux_v I__788 (
            .O(N__5698),
            .I(N__5689));
    Span4Mux_v I__787 (
            .O(N__5695),
            .I(N__5684));
    Span4Mux_v I__786 (
            .O(N__5692),
            .I(N__5684));
    Span4Mux_h I__785 (
            .O(N__5689),
            .I(N__5681));
    Sp12to4 I__784 (
            .O(N__5684),
            .I(N__5678));
    Sp12to4 I__783 (
            .O(N__5681),
            .I(N__5673));
    Span12Mux_h I__782 (
            .O(N__5678),
            .I(N__5673));
    Span12Mux_v I__781 (
            .O(N__5673),
            .I(N__5670));
    Odrv12 I__780 (
            .O(N__5670),
            .I(CLK40_PLL_i));
    InMux I__779 (
            .O(N__5667),
            .I(N__5661));
    InMux I__778 (
            .O(N__5666),
            .I(N__5654));
    InMux I__777 (
            .O(N__5665),
            .I(N__5654));
    InMux I__776 (
            .O(N__5664),
            .I(N__5654));
    LocalMux I__775 (
            .O(N__5661),
            .I(N__5651));
    LocalMux I__774 (
            .O(N__5654),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__773 (
            .O(N__5651),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__772 (
            .O(N__5646),
            .I(N__5642));
    InMux I__771 (
            .O(N__5645),
            .I(N__5639));
    LocalMux I__770 (
            .O(N__5642),
            .I(N__5636));
    LocalMux I__769 (
            .O(N__5639),
            .I(N__5633));
    Odrv4 I__768 (
            .O(N__5636),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    Odrv4 I__767 (
            .O(N__5633),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__766 (
            .O(N__5628),
            .I(N__5624));
    InMux I__765 (
            .O(N__5627),
            .I(N__5621));
    LocalMux I__764 (
            .O(N__5624),
            .I(N__5618));
    LocalMux I__763 (
            .O(N__5621),
            .I(N__5615));
    Span4Mux_v I__762 (
            .O(N__5618),
            .I(N__5612));
    Span4Mux_v I__761 (
            .O(N__5615),
            .I(N__5609));
    Span4Mux_h I__760 (
            .O(N__5612),
            .I(N__5606));
    Sp12to4 I__759 (
            .O(N__5609),
            .I(N__5603));
    Sp12to4 I__758 (
            .O(N__5606),
            .I(N__5598));
    Span12Mux_h I__757 (
            .O(N__5603),
            .I(N__5598));
    Odrv12 I__756 (
            .O(N__5598),
            .I(DBRn_c));
    InMux I__755 (
            .O(N__5595),
            .I(N__5586));
    InMux I__754 (
            .O(N__5594),
            .I(N__5586));
    InMux I__753 (
            .O(N__5593),
            .I(N__5586));
    LocalMux I__752 (
            .O(N__5586),
            .I(DMA_WRITE_CYCLE));
    IoInMux I__751 (
            .O(N__5583),
            .I(N__5580));
    LocalMux I__750 (
            .O(N__5580),
            .I(N__5577));
    IoSpan4Mux I__749 (
            .O(N__5577),
            .I(N__5574));
    IoSpan4Mux I__748 (
            .O(N__5574),
            .I(N__5571));
    Sp12to4 I__747 (
            .O(N__5571),
            .I(N__5568));
    Span12Mux_s7_h I__746 (
            .O(N__5568),
            .I(N__5565));
    Span12Mux_h I__745 (
            .O(N__5565),
            .I(N__5562));
    Odrv12 I__744 (
            .O(N__5562),
            .I(DRDDIR_c));
    CascadeMux I__743 (
            .O(N__5559),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ));
    CEMux I__742 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__741 (
            .O(N__5553),
            .I(N__5550));
    Odrv4 I__740 (
            .O(N__5550),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ));
    CascadeMux I__739 (
            .O(N__5547),
            .I(N__5543));
    InMux I__738 (
            .O(N__5546),
            .I(N__5537));
    InMux I__737 (
            .O(N__5543),
            .I(N__5534));
    CascadeMux I__736 (
            .O(N__5542),
            .I(N__5528));
    CascadeMux I__735 (
            .O(N__5541),
            .I(N__5522));
    CascadeMux I__734 (
            .O(N__5540),
            .I(N__5519));
    LocalMux I__733 (
            .O(N__5537),
            .I(N__5515));
    LocalMux I__732 (
            .O(N__5534),
            .I(N__5512));
    InMux I__731 (
            .O(N__5533),
            .I(N__5507));
    InMux I__730 (
            .O(N__5532),
            .I(N__5507));
    InMux I__729 (
            .O(N__5531),
            .I(N__5503));
    InMux I__728 (
            .O(N__5528),
            .I(N__5500));
    InMux I__727 (
            .O(N__5527),
            .I(N__5497));
    InMux I__726 (
            .O(N__5526),
            .I(N__5494));
    InMux I__725 (
            .O(N__5525),
            .I(N__5485));
    InMux I__724 (
            .O(N__5522),
            .I(N__5485));
    InMux I__723 (
            .O(N__5519),
            .I(N__5485));
    InMux I__722 (
            .O(N__5518),
            .I(N__5485));
    Span4Mux_v I__721 (
            .O(N__5515),
            .I(N__5478));
    Span4Mux_h I__720 (
            .O(N__5512),
            .I(N__5478));
    LocalMux I__719 (
            .O(N__5507),
            .I(N__5478));
    InMux I__718 (
            .O(N__5506),
            .I(N__5475));
    LocalMux I__717 (
            .O(N__5503),
            .I(N__5470));
    LocalMux I__716 (
            .O(N__5500),
            .I(N__5470));
    LocalMux I__715 (
            .O(N__5497),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__714 (
            .O(N__5494),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__713 (
            .O(N__5485),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__712 (
            .O(N__5478),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__711 (
            .O(N__5475),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__710 (
            .O(N__5470),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__709 (
            .O(N__5457),
            .I(\U712_CHIP_RAM.N_503_cascade_ ));
    InMux I__708 (
            .O(N__5454),
            .I(N__5451));
    LocalMux I__707 (
            .O(N__5451),
            .I(\U712_CHIP_RAM.N_420 ));
    CEMux I__706 (
            .O(N__5448),
            .I(N__5445));
    LocalMux I__705 (
            .O(N__5445),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ));
    InMux I__704 (
            .O(N__5442),
            .I(N__5438));
    InMux I__703 (
            .O(N__5441),
            .I(N__5435));
    LocalMux I__702 (
            .O(N__5438),
            .I(N__5432));
    LocalMux I__701 (
            .O(N__5435),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    Odrv4 I__700 (
            .O(N__5432),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__699 (
            .O(N__5427),
            .I(N__5424));
    LocalMux I__698 (
            .O(N__5424),
            .I(N__5421));
    Odrv4 I__697 (
            .O(N__5421),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1 ));
    CascadeMux I__696 (
            .O(N__5418),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    InMux I__695 (
            .O(N__5415),
            .I(N__5412));
    LocalMux I__694 (
            .O(N__5412),
            .I(N__5408));
    InMux I__693 (
            .O(N__5411),
            .I(N__5405));
    Odrv4 I__692 (
            .O(N__5408),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ));
    LocalMux I__691 (
            .O(N__5405),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ));
    CascadeMux I__690 (
            .O(N__5400),
            .I(N__5397));
    InMux I__689 (
            .O(N__5397),
            .I(N__5390));
    InMux I__688 (
            .O(N__5396),
            .I(N__5385));
    InMux I__687 (
            .O(N__5395),
            .I(N__5382));
    InMux I__686 (
            .O(N__5394),
            .I(N__5379));
    InMux I__685 (
            .O(N__5393),
            .I(N__5376));
    LocalMux I__684 (
            .O(N__5390),
            .I(N__5373));
    InMux I__683 (
            .O(N__5389),
            .I(N__5370));
    InMux I__682 (
            .O(N__5388),
            .I(N__5367));
    LocalMux I__681 (
            .O(N__5385),
            .I(N__5360));
    LocalMux I__680 (
            .O(N__5382),
            .I(N__5360));
    LocalMux I__679 (
            .O(N__5379),
            .I(N__5360));
    LocalMux I__678 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__677 (
            .O(N__5373),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__676 (
            .O(N__5370),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__675 (
            .O(N__5367),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__674 (
            .O(N__5360),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__673 (
            .O(N__5349),
            .I(\U712_CHIP_RAM.N_366_cascade_ ));
    InMux I__672 (
            .O(N__5346),
            .I(N__5343));
    LocalMux I__671 (
            .O(N__5343),
            .I(N__5340));
    Span4Mux_v I__670 (
            .O(N__5340),
            .I(N__5336));
    InMux I__669 (
            .O(N__5339),
            .I(N__5333));
    Odrv4 I__668 (
            .O(N__5336),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__667 (
            .O(N__5333),
            .I(\U712_CHIP_RAM.N_335 ));
    CascadeMux I__666 (
            .O(N__5328),
            .I(\U712_CHIP_RAM.DBENn_8_1_cascade_ ));
    IoInMux I__665 (
            .O(N__5325),
            .I(N__5322));
    LocalMux I__664 (
            .O(N__5322),
            .I(N__5319));
    IoSpan4Mux I__663 (
            .O(N__5319),
            .I(N__5316));
    Span4Mux_s2_v I__662 (
            .O(N__5316),
            .I(N__5313));
    Sp12to4 I__661 (
            .O(N__5313),
            .I(N__5310));
    Span12Mux_s11_v I__660 (
            .O(N__5310),
            .I(N__5306));
    InMux I__659 (
            .O(N__5309),
            .I(N__5303));
    Odrv12 I__658 (
            .O(N__5306),
            .I(DBDIR_c));
    LocalMux I__657 (
            .O(N__5303),
            .I(DBDIR_c));
    CascadeMux I__656 (
            .O(N__5298),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_ ));
    InMux I__655 (
            .O(N__5295),
            .I(N__5289));
    InMux I__654 (
            .O(N__5294),
            .I(N__5289));
    LocalMux I__653 (
            .O(N__5289),
            .I(N__5285));
    InMux I__652 (
            .O(N__5288),
            .I(N__5282));
    Span4Mux_h I__651 (
            .O(N__5285),
            .I(N__5277));
    LocalMux I__650 (
            .O(N__5282),
            .I(N__5277));
    Span4Mux_v I__649 (
            .O(N__5277),
            .I(N__5274));
    Sp12to4 I__648 (
            .O(N__5274),
            .I(N__5271));
    Span12Mux_h I__647 (
            .O(N__5271),
            .I(N__5268));
    Odrv12 I__646 (
            .O(N__5268),
            .I(AWEn_c));
    IoInMux I__645 (
            .O(N__5265),
            .I(N__5262));
    LocalMux I__644 (
            .O(N__5262),
            .I(N__5259));
    Span4Mux_s2_v I__643 (
            .O(N__5259),
            .I(N__5256));
    Sp12to4 I__642 (
            .O(N__5256),
            .I(N__5253));
    Span12Mux_h I__641 (
            .O(N__5253),
            .I(N__5250));
    Span12Mux_v I__640 (
            .O(N__5250),
            .I(N__5247));
    Odrv12 I__639 (
            .O(N__5247),
            .I(DMA_LATCH_EN_c));
    CascadeMux I__638 (
            .O(N__5244),
            .I(\U712_CHIP_RAM.N_343_cascade_ ));
    InMux I__637 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__636 (
            .O(N__5238),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    IoInMux I__635 (
            .O(N__5235),
            .I(N__5232));
    LocalMux I__634 (
            .O(N__5232),
            .I(N__5229));
    IoSpan4Mux I__633 (
            .O(N__5229),
            .I(N__5226));
    Span4Mux_s2_v I__632 (
            .O(N__5226),
            .I(N__5222));
    InMux I__631 (
            .O(N__5225),
            .I(N__5219));
    Sp12to4 I__630 (
            .O(N__5222),
            .I(N__5216));
    LocalMux I__629 (
            .O(N__5219),
            .I(N__5213));
    Span12Mux_s8_v I__628 (
            .O(N__5216),
            .I(N__5210));
    Span4Mux_v I__627 (
            .O(N__5213),
            .I(N__5207));
    Span12Mux_v I__626 (
            .O(N__5210),
            .I(N__5202));
    Sp12to4 I__625 (
            .O(N__5207),
            .I(N__5202));
    Span12Mux_h I__624 (
            .O(N__5202),
            .I(N__5199));
    Odrv12 I__623 (
            .O(N__5199),
            .I(A_c_10));
    CascadeMux I__622 (
            .O(N__5196),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__621 (
            .O(N__5193),
            .I(N__5190));
    LocalMux I__620 (
            .O(N__5190),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__619 (
            .O(N__5187),
            .I(N__5184));
    LocalMux I__618 (
            .O(N__5184),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__617 (
            .O(N__5181),
            .I(N__5177));
    InMux I__616 (
            .O(N__5180),
            .I(N__5174));
    LocalMux I__615 (
            .O(N__5177),
            .I(N__5171));
    LocalMux I__614 (
            .O(N__5174),
            .I(N__5168));
    Odrv4 I__613 (
            .O(N__5171),
            .I(\U712_CHIP_RAM.N_334 ));
    Odrv12 I__612 (
            .O(N__5168),
            .I(\U712_CHIP_RAM.N_334 ));
    InMux I__611 (
            .O(N__5163),
            .I(N__5159));
    InMux I__610 (
            .O(N__5162),
            .I(N__5156));
    LocalMux I__609 (
            .O(N__5159),
            .I(N__5153));
    LocalMux I__608 (
            .O(N__5156),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0 ));
    Odrv4 I__607 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0 ));
    InMux I__606 (
            .O(N__5148),
            .I(N__5145));
    LocalMux I__605 (
            .O(N__5145),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1 ));
    InMux I__604 (
            .O(N__5142),
            .I(N__5138));
    InMux I__603 (
            .O(N__5141),
            .I(N__5135));
    LocalMux I__602 (
            .O(N__5138),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__601 (
            .O(N__5135),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__600 (
            .O(N__5130),
            .I(N__5126));
    InMux I__599 (
            .O(N__5129),
            .I(N__5123));
    LocalMux I__598 (
            .O(N__5126),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__597 (
            .O(N__5123),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__596 (
            .O(N__5118),
            .I(N__5114));
    InMux I__595 (
            .O(N__5117),
            .I(N__5111));
    InMux I__594 (
            .O(N__5114),
            .I(N__5108));
    LocalMux I__593 (
            .O(N__5111),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__592 (
            .O(N__5108),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__591 (
            .O(N__5103),
            .I(N__5099));
    InMux I__590 (
            .O(N__5102),
            .I(N__5096));
    LocalMux I__589 (
            .O(N__5099),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__588 (
            .O(N__5096),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__587 (
            .O(N__5091),
            .I(\U712_CHIP_RAM.N_332_cascade_ ));
    CascadeMux I__586 (
            .O(N__5088),
            .I(\U712_CHIP_RAM.N_510_cascade_ ));
    InMux I__585 (
            .O(N__5085),
            .I(N__5082));
    LocalMux I__584 (
            .O(N__5082),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__583 (
            .O(N__5079),
            .I(N__5076));
    LocalMux I__582 (
            .O(N__5076),
            .I(N__5073));
    Span4Mux_s1_v I__581 (
            .O(N__5073),
            .I(N__5070));
    Sp12to4 I__580 (
            .O(N__5070),
            .I(N__5067));
    Span12Mux_h I__579 (
            .O(N__5067),
            .I(N__5064));
    Span12Mux_v I__578 (
            .O(N__5064),
            .I(N__5061));
    Odrv12 I__577 (
            .O(N__5061),
            .I(CMA_c_0));
    IoInMux I__576 (
            .O(N__5058),
            .I(N__5055));
    LocalMux I__575 (
            .O(N__5055),
            .I(N__5052));
    IoSpan4Mux I__574 (
            .O(N__5052),
            .I(N__5049));
    Span4Mux_s2_v I__573 (
            .O(N__5049),
            .I(N__5046));
    Sp12to4 I__572 (
            .O(N__5046),
            .I(N__5043));
    Odrv12 I__571 (
            .O(N__5043),
            .I(CMA_c_1));
    IoInMux I__570 (
            .O(N__5040),
            .I(N__5037));
    LocalMux I__569 (
            .O(N__5037),
            .I(N__5034));
    IoSpan4Mux I__568 (
            .O(N__5034),
            .I(N__5031));
    IoSpan4Mux I__567 (
            .O(N__5031),
            .I(N__5028));
    Sp12to4 I__566 (
            .O(N__5028),
            .I(N__5025));
    Span12Mux_s7_h I__565 (
            .O(N__5025),
            .I(N__5022));
    Span12Mux_h I__564 (
            .O(N__5022),
            .I(N__5019));
    Odrv12 I__563 (
            .O(N__5019),
            .I(CMA_c_5));
    InMux I__562 (
            .O(N__5016),
            .I(N__5013));
    LocalMux I__561 (
            .O(N__5013),
            .I(\U712_CHIP_RAM.N_389 ));
    InMux I__560 (
            .O(N__5010),
            .I(N__5007));
    LocalMux I__559 (
            .O(N__5007),
            .I(\U712_CHIP_RAM.N_504 ));
    CascadeMux I__558 (
            .O(N__5004),
            .I(\U712_CHIP_RAM.N_583_cascade_ ));
    InMux I__557 (
            .O(N__5001),
            .I(N__4998));
    LocalMux I__556 (
            .O(N__4998),
            .I(\U712_CHIP_RAM.N_591 ));
    CascadeMux I__555 (
            .O(N__4995),
            .I(\U712_CHIP_RAM.N_402_cascade_ ));
    InMux I__554 (
            .O(N__4992),
            .I(N__4983));
    InMux I__553 (
            .O(N__4991),
            .I(N__4976));
    InMux I__552 (
            .O(N__4990),
            .I(N__4976));
    InMux I__551 (
            .O(N__4989),
            .I(N__4976));
    InMux I__550 (
            .O(N__4988),
            .I(N__4969));
    InMux I__549 (
            .O(N__4987),
            .I(N__4969));
    InMux I__548 (
            .O(N__4986),
            .I(N__4969));
    LocalMux I__547 (
            .O(N__4983),
            .I(\U712_CHIP_RAM.N_375_0_i ));
    LocalMux I__546 (
            .O(N__4976),
            .I(\U712_CHIP_RAM.N_375_0_i ));
    LocalMux I__545 (
            .O(N__4969),
            .I(\U712_CHIP_RAM.N_375_0_i ));
    InMux I__544 (
            .O(N__4962),
            .I(N__4959));
    LocalMux I__543 (
            .O(N__4959),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0 ));
    CascadeMux I__542 (
            .O(N__4956),
            .I(\U712_CHIP_RAM.N_375_0_i_cascade_ ));
    InMux I__541 (
            .O(N__4953),
            .I(N__4950));
    LocalMux I__540 (
            .O(N__4950),
            .I(\U712_CHIP_RAM.N_402 ));
    CEMux I__539 (
            .O(N__4947),
            .I(N__4943));
    CEMux I__538 (
            .O(N__4946),
            .I(N__4940));
    LocalMux I__537 (
            .O(N__4943),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    LocalMux I__536 (
            .O(N__4940),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__535 (
            .O(N__4935),
            .I(N__4932));
    LocalMux I__534 (
            .O(N__4932),
            .I(\U712_CHIP_RAM.N_426 ));
    IoInMux I__533 (
            .O(N__4929),
            .I(N__4926));
    LocalMux I__532 (
            .O(N__4926),
            .I(N__4923));
    IoSpan4Mux I__531 (
            .O(N__4923),
            .I(N__4920));
    Span4Mux_s1_h I__530 (
            .O(N__4920),
            .I(N__4917));
    Sp12to4 I__529 (
            .O(N__4917),
            .I(N__4914));
    Span12Mux_h I__528 (
            .O(N__4914),
            .I(N__4911));
    Span12Mux_v I__527 (
            .O(N__4911),
            .I(N__4908));
    Odrv12 I__526 (
            .O(N__4908),
            .I(CLK_EN_c));
    InMux I__525 (
            .O(N__4905),
            .I(N__4901));
    InMux I__524 (
            .O(N__4904),
            .I(N__4898));
    LocalMux I__523 (
            .O(N__4901),
            .I(N__4893));
    LocalMux I__522 (
            .O(N__4898),
            .I(N__4893));
    Odrv4 I__521 (
            .O(N__4893),
            .I(\U712_CHIP_RAM.N_586 ));
    InMux I__520 (
            .O(N__4890),
            .I(N__4887));
    LocalMux I__519 (
            .O(N__4887),
            .I(N__4884));
    Odrv4 I__518 (
            .O(N__4884),
            .I(\U712_CHIP_RAM.N_359 ));
    CascadeMux I__517 (
            .O(N__4881),
            .I(\U712_CHIP_RAM.N_586_cascade_ ));
    CascadeMux I__516 (
            .O(N__4878),
            .I(\U712_CHIP_RAM.N_419_cascade_ ));
    CascadeMux I__515 (
            .O(N__4875),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ));
    CascadeMux I__514 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.N_349_cascade_ ));
    InMux I__513 (
            .O(N__4869),
            .I(N__4866));
    LocalMux I__512 (
            .O(N__4866),
            .I(\U712_CHIP_RAM.N_349 ));
    InMux I__511 (
            .O(N__4863),
            .I(N__4860));
    LocalMux I__510 (
            .O(N__4860),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__509 (
            .O(N__4857),
            .I(N__4854));
    InMux I__508 (
            .O(N__4854),
            .I(N__4849));
    InMux I__507 (
            .O(N__4853),
            .I(N__4846));
    InMux I__506 (
            .O(N__4852),
            .I(N__4843));
    LocalMux I__505 (
            .O(N__4849),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__504 (
            .O(N__4846),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__503 (
            .O(N__4843),
            .I(\U712_CHIP_RAM.N_509 ));
    CascadeMux I__502 (
            .O(N__4836),
            .I(\U712_CHIP_RAM.N_509_cascade_ ));
    IoInMux I__501 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__500 (
            .O(N__4830),
            .I(N__4826));
    InMux I__499 (
            .O(N__4829),
            .I(N__4823));
    Span12Mux_s4_v I__498 (
            .O(N__4826),
            .I(N__4820));
    LocalMux I__497 (
            .O(N__4823),
            .I(N__4817));
    Span12Mux_h I__496 (
            .O(N__4820),
            .I(N__4814));
    Span4Mux_v I__495 (
            .O(N__4817),
            .I(N__4811));
    Span12Mux_v I__494 (
            .O(N__4814),
            .I(N__4808));
    Sp12to4 I__493 (
            .O(N__4811),
            .I(N__4805));
    Odrv12 I__492 (
            .O(N__4808),
            .I(A_c_9));
    Odrv12 I__491 (
            .O(N__4805),
            .I(A_c_9));
    CascadeMux I__490 (
            .O(N__4800),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    IoInMux I__489 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__488 (
            .O(N__4794),
            .I(N__4791));
    Span12Mux_s8_v I__487 (
            .O(N__4791),
            .I(N__4788));
    Odrv12 I__486 (
            .O(N__4788),
            .I(VBENn_c));
    IoInMux I__485 (
            .O(N__4785),
            .I(N__4782));
    LocalMux I__484 (
            .O(N__4782),
            .I(N__4779));
    Span12Mux_s6_v I__483 (
            .O(N__4779),
            .I(N__4776));
    Span12Mux_h I__482 (
            .O(N__4776),
            .I(N__4773));
    Odrv12 I__481 (
            .O(N__4773),
            .I(CMA_c_10));
    IoInMux I__480 (
            .O(N__4770),
            .I(N__4767));
    LocalMux I__479 (
            .O(N__4767),
            .I(N__4764));
    IoSpan4Mux I__478 (
            .O(N__4764),
            .I(N__4761));
    Span4Mux_s2_v I__477 (
            .O(N__4761),
            .I(N__4758));
    Sp12to4 I__476 (
            .O(N__4758),
            .I(N__4755));
    Span12Mux_s8_v I__475 (
            .O(N__4755),
            .I(N__4751));
    InMux I__474 (
            .O(N__4754),
            .I(N__4748));
    Span12Mux_v I__473 (
            .O(N__4751),
            .I(N__4745));
    LocalMux I__472 (
            .O(N__4748),
            .I(N__4742));
    Span12Mux_h I__471 (
            .O(N__4745),
            .I(N__4737));
    Span12Mux_v I__470 (
            .O(N__4742),
            .I(N__4737));
    Odrv12 I__469 (
            .O(N__4737),
            .I(A_c_11));
    CascadeMux I__468 (
            .O(N__4734),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    CascadeMux I__467 (
            .O(N__4731),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ));
    IoInMux I__466 (
            .O(N__4728),
            .I(N__4725));
    LocalMux I__465 (
            .O(N__4725),
            .I(N__4722));
    Span4Mux_s3_v I__464 (
            .O(N__4722),
            .I(N__4719));
    Sp12to4 I__463 (
            .O(N__4719),
            .I(N__4716));
    Span12Mux_h I__462 (
            .O(N__4716),
            .I(N__4713));
    Span12Mux_v I__461 (
            .O(N__4713),
            .I(N__4710));
    Odrv12 I__460 (
            .O(N__4710),
            .I(CMA_c_2));
    CascadeMux I__459 (
            .O(N__4707),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER19_cascade_ ));
    CascadeMux I__458 (
            .O(N__4704),
            .I(\U712_CHIP_RAM.N_335_cascade_ ));
    CascadeMux I__457 (
            .O(N__4701),
            .I(\U712_CHIP_RAM.N_507_cascade_ ));
    InMux I__456 (
            .O(N__4698),
            .I(N__4695));
    LocalMux I__455 (
            .O(N__4695),
            .I(N__4692));
    Odrv4 I__454 (
            .O(N__4692),
            .I(\U712_CHIP_RAM.N_477 ));
    CascadeMux I__453 (
            .O(N__4689),
            .I(\U712_CHIP_RAM.N_477_cascade_ ));
    InMux I__452 (
            .O(N__4686),
            .I(N__4679));
    InMux I__451 (
            .O(N__4685),
            .I(N__4679));
    InMux I__450 (
            .O(N__4684),
            .I(N__4676));
    LocalMux I__449 (
            .O(N__4679),
            .I(N__4673));
    LocalMux I__448 (
            .O(N__4676),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__447 (
            .O(N__4673),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__446 (
            .O(N__4668),
            .I(\U712_CYCLE_TERM.N_406_cascade_ ));
    IoInMux I__445 (
            .O(N__4665),
            .I(N__4662));
    LocalMux I__444 (
            .O(N__4662),
            .I(N__4659));
    Span4Mux_s3_h I__443 (
            .O(N__4659),
            .I(N__4656));
    Sp12to4 I__442 (
            .O(N__4656),
            .I(N__4653));
    Span12Mux_v I__441 (
            .O(N__4653),
            .I(N__4649));
    InMux I__440 (
            .O(N__4652),
            .I(N__4646));
    Odrv12 I__439 (
            .O(N__4649),
            .I(TACK_OUT));
    LocalMux I__438 (
            .O(N__4646),
            .I(TACK_OUT));
    InMux I__437 (
            .O(N__4641),
            .I(N__4638));
    LocalMux I__436 (
            .O(N__4638),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0 ));
    InMux I__435 (
            .O(N__4635),
            .I(N__4632));
    LocalMux I__434 (
            .O(N__4632),
            .I(\U712_CHIP_RAM.N_478 ));
    InMux I__433 (
            .O(N__4629),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__432 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__431 (
            .O(N__4623),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__430 (
            .O(N__4620),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__429 (
            .O(N__4617),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__428 (
            .O(N__4614),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__427 (
            .O(N__4611),
            .I(N__4608));
    LocalMux I__426 (
            .O(N__4608),
            .I(N__4605));
    Odrv4 I__425 (
            .O(N__4605),
            .I(\U712_CHIP_RAM.N_483 ));
    IoInMux I__424 (
            .O(N__4602),
            .I(N__4598));
    IoInMux I__423 (
            .O(N__4601),
            .I(N__4595));
    LocalMux I__422 (
            .O(N__4598),
            .I(N__4592));
    LocalMux I__421 (
            .O(N__4595),
            .I(N__4589));
    IoSpan4Mux I__420 (
            .O(N__4592),
            .I(N__4584));
    IoSpan4Mux I__419 (
            .O(N__4589),
            .I(N__4584));
    Span4Mux_s3_v I__418 (
            .O(N__4584),
            .I(N__4581));
    Sp12to4 I__417 (
            .O(N__4581),
            .I(N__4577));
    IoInMux I__416 (
            .O(N__4580),
            .I(N__4574));
    Span12Mux_v I__415 (
            .O(N__4577),
            .I(N__4571));
    LocalMux I__414 (
            .O(N__4574),
            .I(N__4568));
    Span12Mux_h I__413 (
            .O(N__4571),
            .I(N__4563));
    Span12Mux_s5_h I__412 (
            .O(N__4568),
            .I(N__4563));
    Odrv12 I__411 (
            .O(N__4563),
            .I(CLK40_PLL_i_i));
    CascadeMux I__410 (
            .O(N__4560),
            .I(\U712_CHIP_RAM.N_592_cascade_ ));
    CascadeMux I__409 (
            .O(N__4557),
            .I(\U712_CHIP_RAM.N_482_cascade_ ));
    InMux I__408 (
            .O(N__4554),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    IoInMux I__407 (
            .O(N__4551),
            .I(N__4548));
    LocalMux I__406 (
            .O(N__4548),
            .I(N__4545));
    Span4Mux_s3_h I__405 (
            .O(N__4545),
            .I(N__4542));
    Odrv4 I__404 (
            .O(N__4542),
            .I(DBRn_c_i_0));
    IoInMux I__403 (
            .O(N__4539),
            .I(N__4536));
    LocalMux I__402 (
            .O(N__4536),
            .I(N__4533));
    IoSpan4Mux I__401 (
            .O(N__4533),
            .I(N__4530));
    Span4Mux_s2_v I__400 (
            .O(N__4530),
            .I(N__4527));
    Span4Mux_v I__399 (
            .O(N__4527),
            .I(N__4524));
    Odrv4 I__398 (
            .O(N__4524),
            .I(CLK80_PLL_iso_i));
    IoInMux I__397 (
            .O(N__4521),
            .I(N__4518));
    LocalMux I__396 (
            .O(N__4518),
            .I(N__4515));
    Span4Mux_s0_v I__395 (
            .O(N__4515),
            .I(N__4512));
    Span4Mux_v I__394 (
            .O(N__4512),
            .I(N__4509));
    Sp12to4 I__393 (
            .O(N__4509),
            .I(N__4506));
    Span12Mux_h I__392 (
            .O(N__4506),
            .I(N__4503));
    Span12Mux_v I__391 (
            .O(N__4503),
            .I(N__4500));
    Odrv12 I__390 (
            .O(N__4500),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__9627));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__9624));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__9625));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__9626));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__9629));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__9628));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__9630));
    INV \INVU712_CYCLE_TERM.TACK_STATE_1C  (
            .O(\INVU712_CYCLE_TERM.TACK_STATE_1C_net ),
            .I(N__10220));
    INV \INVU712_CYCLE_TERM.TACK_OUTC  (
            .O(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .I(N__10228));
    INV \INVU712_CYCLE_TERM.TACK_STATE_3C  (
            .O(\INVU712_CYCLE_TERM.TACK_STATE_3C_net ),
            .I(N__10231));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5967),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9348),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4551),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__7494),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__7544),
            .in2(_gnd_net_),
            .in3(N__10725),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_5.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_5.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10236),
            .lcout(CLK80_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_6_12_4.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5628),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_6_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5646),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_3C_net ),
            .ce(),
            .sr(N__10673));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4684),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_3C_net ),
            .ce(),
            .sr(N__10673));
    defparam pll_RNI8MQ3_LC_7_10_1.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_7_10_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_7_10_1 (
            .in0(N__5713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_7_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_7_11_0  (
            .in0(N__5506),
            .in1(N__7130),
            .in2(_gnd_net_),
            .in3(N__6548),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_11_1  (
            .in0(N__10446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5858),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_11_2 .LUT_INIT=16'b1010101100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_11_2  (
            .in0(N__6774),
            .in1(N__4698),
            .in2(N__4560),
            .in3(N__8699),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10213),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_11_4 .LUT_INIT=16'b0000010000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_11_4  (
            .in0(N__6472),
            .in1(N__6549),
            .in2(N__7158),
            .in3(N__8338),
            .lcout(\U712_CHIP_RAM.N_334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_11_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_11_6  (
            .in0(N__5859),
            .in1(N__10445),
            .in2(N__5400),
            .in3(N__8339),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_7_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_7_11_7 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_7_11_7  (
            .in0(N__4611),
            .in1(N__6773),
            .in2(N__4557),
            .in3(N__9996),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10213),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_7_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_7_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__8335),
            .in2(_gnd_net_),
            .in3(N__11097),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_12_1  (
            .in0(N__4989),
            .in1(N__7138),
            .in2(_gnd_net_),
            .in3(N__4554),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__6574),
            .in2(_gnd_net_),
            .in3(N__4629),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_12_3  (
            .in0(N__4990),
            .in1(N__6473),
            .in2(_gnd_net_),
            .in3(N__4626),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_12_4  (
            .in0(N__4986),
            .in1(N__5117),
            .in2(_gnd_net_),
            .in3(N__4623),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_12_5  (
            .in0(N__4991),
            .in1(N__5130),
            .in2(_gnd_net_),
            .in3(N__4620),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_12_6  (
            .in0(N__4987),
            .in1(N__5142),
            .in2(_gnd_net_),
            .in3(N__4617),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_12_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_12_7  (
            .in0(N__5103),
            .in1(N__4988),
            .in2(_gnd_net_),
            .in3(N__4614),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10218),
            .ce(N__4947),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_7_13_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_7_13_0  (
            .in0(N__10500),
            .in1(N__8364),
            .in2(_gnd_net_),
            .in3(N__6552),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_13_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_13_1  (
            .in0(N__4852),
            .in1(N__8359),
            .in2(N__7049),
            .in3(N__5533),
            .lcout(\U712_CHIP_RAM.N_483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2EV43_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2EV43_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2EV43_LC_7_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2EV43_LC_7_13_2  (
            .in0(N__5532),
            .in1(N__6551),
            .in2(N__7157),
            .in3(N__7030),
            .lcout(\U712_CHIP_RAM.N_590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_7_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_7_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__8357),
            .in2(_gnd_net_),
            .in3(N__7134),
            .lcout(\U712_CHIP_RAM.N_335 ),
            .ltout(\U712_CHIP_RAM.N_335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_3_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_3_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_3_LC_7_13_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_3_LC_7_13_4  (
            .in0(N__10501),
            .in1(N__6471),
            .in2(N__4704),
            .in3(N__6553),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5EAU6_3_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5EAU6_3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5EAU6_3_LC_7_13_5 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5EAU6_3_LC_7_13_5  (
            .in0(N__5163),
            .in1(N__7042),
            .in2(N__4701),
            .in3(N__5181),
            .lcout(\U712_CHIP_RAM.N_477 ),
            .ltout(\U712_CHIP_RAM.N_477_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_7_13_6 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_7_13_6  (
            .in0(N__4635),
            .in1(N__6766),
            .in2(N__4689),
            .in3(N__7592),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10223),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIN90C1_LC_7_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIN90C1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIN90C1_LC_7_13_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIN90C1_LC_7_13_7  (
            .in0(N__11088),
            .in1(N__10499),
            .in2(N__5547),
            .in3(N__8358),
            .lcout(\U712_CHIP_RAM.N_504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_14_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__4685),
            .in2(_gnd_net_),
            .in3(N__5645),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_7_14_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_7_14_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__5712),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_7_14_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_7_14_3 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_LC_7_14_3  (
            .in0(N__10496),
            .in1(N__4686),
            .in2(N__4668),
            .in3(N__4652),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_14_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_14_5  (
            .in0(N__7159),
            .in1(N__4641),
            .in2(N__7058),
            .in3(N__5546),
            .lcout(\U712_CHIP_RAM.N_478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5  (
            .in0(N__4829),
            .in1(N__6240),
            .in2(_gnd_net_),
            .in3(N__8002),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_8_8_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_8_8_6  (
            .in0(N__8003),
            .in1(N__11893),
            .in2(N__4800),
            .in3(N__8652),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_9_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_9_6  (
            .in0(N__8844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11902),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_8_10_3 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_8_10_3  (
            .in0(N__8000),
            .in1(N__6051),
            .in2(N__8712),
            .in3(_gnd_net_),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10204),
            .ce(N__6315),
            .sr(N__10686));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_10_5  (
            .in0(N__7998),
            .in1(N__4754),
            .in2(_gnd_net_),
            .in3(N__6681),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_8_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_8_10_6  (
            .in0(N__11901),
            .in1(N__7999),
            .in2(N__4734),
            .in3(N__8859),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_8_10_7 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_8_10_7  (
            .in0(N__6356),
            .in1(N__6052),
            .in2(N__4731),
            .in3(N__9705),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10204),
            .ce(N__6315),
            .sr(N__10686));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_11_0  (
            .in0(N__8342),
            .in1(N__4904),
            .in2(N__7163),
            .in3(N__6561),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_11_1 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__10451),
            .in2(N__4707),
            .in3(N__5525),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10210),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIGDNC1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIGDNC1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIGDNC1_LC_8_11_2 .LUT_INIT=16'b0000011100010111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIGDNC1_LC_8_11_2  (
            .in0(N__8340),
            .in1(N__6559),
            .in2(N__5540),
            .in3(N__5389),
            .lcout(\U712_CHIP_RAM.N_349 ),
            .ltout(\U712_CHIP_RAM.N_349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI6NJS1_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI6NJS1_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI6NJS1_LC_8_11_3 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI6NJS1_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__10455),
            .in2(N__4872),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_11_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_11_4  (
            .in0(N__8341),
            .in1(N__6560),
            .in2(N__5541),
            .in3(N__6816),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__10452),
            .in2(_gnd_net_),
            .in3(N__5518),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_11_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_11_6  (
            .in0(N__10454),
            .in1(N__4853),
            .in2(_gnd_net_),
            .in3(N__4869),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_11_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__10453),
            .in2(_gnd_net_),
            .in3(N__6464),
            .lcout(\U712_CHIP_RAM.N_501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0  (
            .in0(N__4863),
            .in1(N__6870),
            .in2(N__4857),
            .in3(N__4992),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10214),
            .ce(N__4946),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILQND1_3_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILQND1_3_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILQND1_3_LC_8_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILQND1_3_LC_8_12_1  (
            .in0(N__6466),
            .in1(N__10497),
            .in2(_gnd_net_),
            .in3(N__6557),
            .lcout(\U712_CHIP_RAM.N_509 ),
            .ltout(\U712_CHIP_RAM.N_509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_2 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_2  (
            .in0(N__7274),
            .in1(N__7200),
            .in2(N__4836),
            .in3(N__7356),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7F93_1_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7F93_1_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7F93_1_LC_8_12_3 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7F93_1_LC_8_12_3  (
            .in0(N__6465),
            .in1(N__10498),
            .in2(N__7066),
            .in3(N__7173),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_583_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI615I6_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI615I6_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI615I6_LC_8_12_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI615I6_LC_8_12_4  (
            .in0(N__5010),
            .in1(N__6812),
            .in2(N__5004),
            .in3(N__5339),
            .lcout(\U712_CHIP_RAM.N_402 ),
            .ltout(\U712_CHIP_RAM.N_402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSQMA_3_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSQMA_3_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISSQMA_3_LC_8_12_5 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISSQMA_3_LC_8_12_5  (
            .in0(N__6467),
            .in1(N__5001),
            .in2(N__4995),
            .in3(N__4935),
            .lcout(\U712_CHIP_RAM.N_375_0_i ),
            .ltout(\U712_CHIP_RAM.N_375_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_12_6 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_12_6  (
            .in0(N__4962),
            .in1(N__8259),
            .in2(N__4956),
            .in3(N__4953),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10214),
            .ce(N__4946),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_8_12_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_8_12_7  (
            .in0(N__6811),
            .in1(N__6558),
            .in2(_gnd_net_),
            .in3(N__5527),
            .lcout(\U712_CHIP_RAM.N_426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_8_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_8_13_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_8_13_0  (
            .in0(N__6556),
            .in1(N__7124),
            .in2(N__8378),
            .in3(N__4905),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10219),
            .ce(N__5556),
            .sr(N__10665));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_8_13_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__6454),
            .in2(_gnd_net_),
            .in3(N__7035),
            .lcout(\U712_CHIP_RAM.N_586 ),
            .ltout(\U712_CHIP_RAM.N_586_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_13_2  (
            .in0(N__8360),
            .in1(N__4890),
            .in2(N__4881),
            .in3(N__10471),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_419_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIADE59_2_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIADE59_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIADE59_2_LC_8_13_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIADE59_2_LC_8_13_3  (
            .in0(N__6824),
            .in1(N__6555),
            .in2(N__4878),
            .in3(N__7354),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOV5BI_2_LC_8_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOV5BI_2_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOV5BI_2_LC_8_13_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOV5BI_2_LC_8_13_4  (
            .in0(N__5454),
            .in1(N__7729),
            .in2(N__4875),
            .in3(N__10472),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_13_5  (
            .in0(N__5141),
            .in1(N__5129),
            .in2(N__5118),
            .in3(N__5102),
            .lcout(\U712_CHIP_RAM.N_332 ),
            .ltout(\U712_CHIP_RAM.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_8_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_8_13_6  (
            .in0(N__6455),
            .in1(N__7123),
            .in2(N__5091),
            .in3(N__5531),
            .lcout(\U712_CHIP_RAM.N_510 ),
            .ltout(\U712_CHIP_RAM.N_510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_13_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_13_7  (
            .in0(N__8365),
            .in1(N__6554),
            .in2(N__5088),
            .in3(N__5395),
            .lcout(\U712_CHIP_RAM.N_461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_14_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_14_0  (
            .in0(N__7275),
            .in1(N__7308),
            .in2(_gnd_net_),
            .in3(N__7358),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10224),
            .ce(N__5448),
            .sr(N__10654));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_17_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_17_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_8_17_0  (
            .in0(N__11621),
            .in1(N__11558),
            .in2(N__6942),
            .in3(N__11430),
            .lcout(\U712_REG_SM.N_429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_9_8_5 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_9_8_5  (
            .in0(N__6357),
            .in1(N__8640),
            .in2(N__6060),
            .in3(N__5085),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10193),
            .ce(N__6314),
            .sr(N__10691));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_9_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_9_9_2  (
            .in0(N__5241),
            .in1(N__5187),
            .in2(_gnd_net_),
            .in3(N__5193),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10196),
            .ce(N__6307),
            .sr(N__10687));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_9_6 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_9_9_6  (
            .in0(N__6162),
            .in1(N__6053),
            .in2(N__8007),
            .in3(N__5016),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10196),
            .ce(N__6307),
            .sr(N__10687));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_10_0  (
            .in0(N__11869),
            .in1(N__6651),
            .in2(_gnd_net_),
            .in3(N__7506),
            .lcout(\U712_CHIP_RAM.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__7611),
            .in2(_gnd_net_),
            .in3(N__10009),
            .lcout(\U712_CHIP_RAM.N_343 ),
            .ltout(\U712_CHIP_RAM.N_343_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_10_2 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_10_2  (
            .in0(N__9339),
            .in1(N__11868),
            .in2(N__5244),
            .in3(N__7963),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_10_4  (
            .in0(N__5225),
            .in1(N__6705),
            .in2(_gnd_net_),
            .in3(N__7958),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_10_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_10_5  (
            .in0(N__7964),
            .in1(N__11871),
            .in2(N__5196),
            .in3(N__8868),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_10_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_10_6  (
            .in0(N__10010),
            .in1(N__7612),
            .in2(_gnd_net_),
            .in3(N__7959),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_10_7 .LUT_INIT=16'b0000010110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_10_7  (
            .in0(N__6036),
            .in1(N__9338),
            .in2(N__7989),
            .in3(N__11870),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_11_0 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_11_0  (
            .in0(N__5180),
            .in1(N__5162),
            .in2(N__7068),
            .in3(N__5148),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_11_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_11_1  (
            .in0(N__8336),
            .in1(N__5388),
            .in2(_gnd_net_),
            .in3(N__6550),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_2  (
            .in0(N__7273),
            .in1(N__6966),
            .in2(_gnd_net_),
            .in3(N__5295),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3  (
            .in0(N__5393),
            .in1(N__6869),
            .in2(N__5349),
            .in3(N__7304),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10205),
            .ce(),
            .sr(N__10674));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_11_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_9_11_5  (
            .in0(N__5346),
            .in1(N__7303),
            .in2(_gnd_net_),
            .in3(N__7065),
            .lcout(),
            .ltout(\U712_CHIP_RAM.DBENn_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_9_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_9_11_6 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_9_11_6  (
            .in0(N__11158),
            .in1(N__5415),
            .in2(N__5328),
            .in3(N__9132),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10205),
            .ce(),
            .sr(N__10674));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_11_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_11_7  (
            .in0(N__5294),
            .in1(N__5309),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10205),
            .ce(),
            .sr(N__10674));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__5394),
            .in2(_gnd_net_),
            .in3(N__6547),
            .lcout(\U712_CHIP_RAM.N_350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQS0H1_1_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQS0H1_1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQS0H1_1_LC_9_12_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQS0H1_1_LC_9_12_1  (
            .in0(N__8337),
            .in1(N__6476),
            .in2(N__7172),
            .in3(N__11813),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN2IA4_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN2IA4_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN2IA4_LC_9_12_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN2IA4_LC_9_12_2  (
            .in0(N__6854),
            .in1(N__5526),
            .in2(N__5298),
            .in3(N__7034),
            .lcout(\U712_CHIP_RAM.N_476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_12_3 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_12_3  (
            .in0(N__5288),
            .in1(N__5593),
            .in2(N__10502),
            .in3(N__5441),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10211),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_9_12_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_9_12_4  (
            .in0(N__5594),
            .in1(N__11357),
            .in2(_gnd_net_),
            .in3(N__11268),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_9_12_5 .LUT_INIT=16'b0010000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_9_12_5  (
            .in0(N__11358),
            .in1(N__6965),
            .in2(N__11276),
            .in3(N__5595),
            .lcout(DRDDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_9_12_6 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_9_12_6  (
            .in0(N__6573),
            .in1(N__5837),
            .in2(N__8382),
            .in3(N__7723),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_12_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5559),
            .in3(N__10723),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_9_13_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_9_13_0  (
            .in0(N__7164),
            .in1(N__8333),
            .in2(N__5542),
            .in3(N__7029),
            .lcout(\U712_CHIP_RAM.N_503 ),
            .ltout(\U712_CHIP_RAM.N_503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNILPRG5_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNILPRG5_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNILPRG5_LC_9_13_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNILPRG5_LC_9_13_1  (
            .in0(N__7193),
            .in1(N__7254),
            .in2(N__5457),
            .in3(N__6823),
            .lcout(\U712_CHIP_RAM.N_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_2  (
            .in0(N__10722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5411),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_13_3  (
            .in0(N__7299),
            .in1(N__7255),
            .in2(_gnd_net_),
            .in3(N__7353),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIAGI99_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIAGI99_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIAGI99_LC_9_13_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIAGI99_LC_9_13_4  (
            .in0(N__5427),
            .in1(N__7758),
            .in2(N__5418),
            .in3(N__7722),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_13_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_13_5  (
            .in0(N__8334),
            .in1(N__5396),
            .in2(_gnd_net_),
            .in3(N__6480),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_13_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_13_6  (
            .in0(N__5857),
            .in1(N__5838),
            .in2(N__5826),
            .in3(N__7694),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_13_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5823),
            .in3(N__10721),
            .lcout(\U712_CHIP_RAM.N_248_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_14_0 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_14_0  (
            .in0(N__5666),
            .in1(N__5714),
            .in2(N__5802),
            .in3(N__5820),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_1C_net ),
            .ce(),
            .sr(N__10651));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_14_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_14_1  (
            .in0(N__6901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6983),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_2 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_2  (
            .in0(N__5665),
            .in1(N__5790),
            .in2(N__5814),
            .in3(N__5811),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_1C_net ),
            .ce(),
            .sr(N__10651));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_14_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_14_3  (
            .in0(N__6902),
            .in1(N__5798),
            .in2(_gnd_net_),
            .in3(N__6984),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_358_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_14_4 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__5789),
            .in2(N__5778),
            .in3(N__5733),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_1C_net ),
            .ce(),
            .sr(N__10651));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_14_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_14_5  (
            .in0(N__5715),
            .in1(N__5664),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_1C_net ),
            .ce(),
            .sr(N__10651));
    defparam DBR_SYNC_0_LC_9_15_3.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_9_15_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_9_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_9_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5627),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10225),
            .ce(),
            .sr(N__10649));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5937),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10225),
            .ce(),
            .sr(N__10649));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_16_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__8513),
            .in2(_gnd_net_),
            .in3(N__9409),
            .lcout(\U712_REG_SM.N_352 ),
            .ltout(\U712_REG_SM.N_352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_16_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_16_2  (
            .in0(N__10503),
            .in1(N__8198),
            .in2(N__5970),
            .in3(N__7401),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10229),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_9_16_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_9_16_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__8514),
            .in2(_gnd_net_),
            .in3(N__9410),
            .lcout(\U712_REG_SM.N_353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_17_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_17_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_17_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_17_0  (
            .in0(N__5963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(),
            .sr(N__10647));
    defparam \U712_REG_SM.UDSn_LC_9_17_3 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_9_17_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_9_17_3 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_REG_SM.UDSn_LC_9_17_3  (
            .in0(N__5912),
            .in1(N__8762),
            .in2(N__9446),
            .in3(N__5865),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(),
            .sr(N__10647));
    defparam \U712_REG_SM.LDSn_LC_9_17_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_9_17_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_9_17_6 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U712_REG_SM.LDSn_LC_9_17_6  (
            .in0(N__5901),
            .in1(N__9436),
            .in2(N__5882),
            .in3(N__8763),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(),
            .sr(N__10647));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_18_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_18_7 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_9_18_7  (
            .in0(N__6952),
            .in1(N__11638),
            .in2(N__11575),
            .in3(N__11453),
            .lcout(\U712_REG_SM.N_493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_8_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_8_0  (
            .in0(N__7967),
            .in1(N__11873),
            .in2(N__6213),
            .in3(N__7512),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_8_1  (
            .in0(N__7965),
            .in1(N__6591),
            .in2(_gnd_net_),
            .in3(N__6228),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_2  (
            .in0(N__6204),
            .in1(N__7966),
            .in2(_gnd_net_),
            .in3(N__7776),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_3  (
            .in0(N__11874),
            .in1(N__7968),
            .in2(N__6180),
            .in3(N__7523),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_6  (
            .in0(N__6177),
            .in1(N__11872),
            .in2(_gnd_net_),
            .in3(N__8607),
            .lcout(\U712_CHIP_RAM.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_9_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_10_9_0  (
            .in0(N__6345),
            .in1(N__8619),
            .in2(N__6057),
            .in3(N__6264),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_10_9_1 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_10_9_1  (
            .in0(N__6049),
            .in1(N__6346),
            .in2(N__9903),
            .in3(N__8073),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_10_9_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_10_9_2  (
            .in0(N__6347),
            .in1(N__9324),
            .in2(N__6058),
            .in3(N__8031),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_10_9_3 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_10_9_3  (
            .in0(N__6050),
            .in1(N__6348),
            .in2(N__6093),
            .in3(N__8877),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_10_9_4 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_10_9_4  (
            .in0(N__6349),
            .in1(N__8628),
            .in2(N__6059),
            .in3(N__5997),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_10_9_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_10_9_5  (
            .in0(N__6405),
            .in1(N__6399),
            .in2(N__11903),
            .in3(N__10800),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10194),
            .ce(N__6306),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_10_10_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_10_10_0  (
            .in0(N__7955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11863),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_1  (
            .in0(N__10008),
            .in1(N__7953),
            .in2(N__7616),
            .in3(N__8713),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_10_2 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_10_2  (
            .in0(N__7954),
            .in1(N__7610),
            .in2(N__6321),
            .in3(N__8714),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_10_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6318),
            .in3(N__10724),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_10_4 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_10_4  (
            .in0(N__10425),
            .in1(N__8946),
            .in2(N__8067),
            .in3(N__9005),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10197),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_5  (
            .in0(N__6282),
            .in1(N__6615),
            .in2(_gnd_net_),
            .in3(N__7956),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_10_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_10_6  (
            .in0(N__7957),
            .in1(N__11864),
            .in2(N__6267),
            .in3(N__9123),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_10_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6258),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_11_1  (
            .in0(N__6720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_10_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_10_11_2  (
            .in0(N__6699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_10_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_10_11_3  (
            .in0(N__6669),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6645),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_11_5  (
            .in0(N__6633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6609),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10200),
            .ce(N__7829),
            .sr(N__10666));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_12_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_12_0  (
            .in0(N__6475),
            .in1(N__8369),
            .in2(N__6579),
            .in3(N__11839),
            .lcout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__6575),
            .in2(_gnd_net_),
            .in3(N__6474),
            .lcout(\U712_CHIP_RAM.N_514 ),
            .ltout(\U712_CHIP_RAM.N_514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_12_2  (
            .in0(N__7260),
            .in1(N__7357),
            .in2(N__6873),
            .in3(N__7368),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10206),
            .ce(N__6840),
            .sr(N__10655));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIVM1I4_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIVM1I4_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIVM1I4_LC_10_12_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIVM1I4_LC_10_12_3  (
            .in0(N__7367),
            .in1(N__7259),
            .in2(_gnd_net_),
            .in3(N__7355),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_0_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_0_LC_10_12_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_0_LC_10_12_4  (
            .in0(N__7790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10720),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_5 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_5  (
            .in0(N__6855),
            .in1(N__7736),
            .in2(N__8379),
            .in3(N__7789),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6843),
            .in3(N__10719),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_13_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_13_0  (
            .in0(N__8151),
            .in1(N__7252),
            .in2(N__7359),
            .in3(N__6828),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_481_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_13_1 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_13_1  (
            .in0(N__6783),
            .in1(N__6772),
            .in2(N__6747),
            .in3(N__7981),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10212),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_10_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__6888),
            .in2(_gnd_net_),
            .in3(N__8219),
            .lcout(),
            .ltout(\U712_REG_SM.N_428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_3 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_10_13_3  (
            .in0(N__10477),
            .in1(N__8138),
            .in2(N__6744),
            .in3(N__6741),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10212),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_0_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_0_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_0_LC_10_13_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_0_LC_10_13_4  (
            .in0(N__8149),
            .in1(N__7214),
            .in2(_gnd_net_),
            .in3(N__8086),
            .lcout(\U712_CHIP_RAM.N_500 ),
            .ltout(\U712_CHIP_RAM.N_500_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_13_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_13_5  (
            .in0(N__7251),
            .in1(N__7349),
            .in2(N__7311),
            .in3(N__7298),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_13_6 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_13_6  (
            .in0(N__8775),
            .in1(N__10476),
            .in2(N__11142),
            .in3(N__7253),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10212),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_13_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_13_7  (
            .in0(N__8087),
            .in1(N__8150),
            .in2(_gnd_net_),
            .in3(N__7215),
            .lcout(\U712_CHIP_RAM.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_10_14_2 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_LC_10_14_2  (
            .in0(N__7182),
            .in1(N__7171),
            .in2(_gnd_net_),
            .in3(N__7067),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10215),
            .ce(N__6975),
            .sr(N__10650));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_15_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_10_15_0  (
            .in0(N__8591),
            .in1(N__7399),
            .in2(_gnd_net_),
            .in3(N__6958),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam DBR_SYNC_1_LC_10_15_1.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_10_15_1.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_10_15_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_1_LC_10_15_1 (
            .in0(N__6912),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.REG_TACK_LC_10_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_15_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_15_2  (
            .in0(N__8550),
            .in1(N__8556),
            .in2(N__6906),
            .in3(N__8568),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.START_RST_LC_10_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_10_15_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_10_15_3  (
            .in0(N__7400),
            .in1(N__6887),
            .in2(_gnd_net_),
            .in3(N__8197),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7475),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.REGENn_LC_10_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_10_15_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_10_15_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \U712_REG_SM.REGENn_LC_10_15_6  (
            .in0(N__8166),
            .in1(N__7423),
            .in2(_gnd_net_),
            .in3(N__9506),
            .lcout(BLSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7410),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10221),
            .ce(),
            .sr(N__10648));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_10_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_10_16_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__8516),
            .in2(_gnd_net_),
            .in3(N__9412),
            .lcout(\U712_REG_SM.N_345 ),
            .ltout(\U712_REG_SM.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_10_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_10_16_1 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__9477),
            .in2(N__7404),
            .in3(N__8223),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_16_2 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_10_16_2  (
            .in0(N__7656),
            .in1(N__7386),
            .in2(N__9443),
            .in3(N__10506),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10226),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_16_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_16_3  (
            .in0(N__8193),
            .in1(N__8544),
            .in2(_gnd_net_),
            .in3(N__7377),
            .lcout(\U712_REG_SM.N_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_10_16_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_10_16_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_10_16_4  (
            .in0(N__8474),
            .in1(N__8515),
            .in2(_gnd_net_),
            .in3(N__9411),
            .lcout(\U712_REG_SM.N_435 ),
            .ltout(\U712_REG_SM.N_435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_10_16_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_10_16_5 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_10_16_5  (
            .in0(N__8192),
            .in1(_gnd_net_),
            .in2(N__7380),
            .in3(N__7376),
            .lcout(\U712_REG_SM.N_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_16_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__8983),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(\U712_REG_SM.N_357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_16_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_16_7  (
            .in0(N__8590),
            .in1(N__8475),
            .in2(N__7650),
            .in3(N__8821),
            .lcout(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_10_17_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_10_17_2 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_10_17_2  (
            .in0(N__8745),
            .in1(N__7649),
            .in2(N__8484),
            .in3(N__10509),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10230),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_3_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_3_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_3_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_11_6_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_11_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8001),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10187),
            .ce(),
            .sr(N__10692));
    defparam \U712_CHIP_RAM.RASn_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_11_7_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_11_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7617),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10191),
            .ce(),
            .sr(N__10688));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_8_1 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_8_1  (
            .in0(N__11042),
            .in1(N__10862),
            .in2(N__7551),
            .in3(N__7524),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__10683));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_0  (
            .in0(N__11038),
            .in1(N__10863),
            .in2(_gnd_net_),
            .in3(N__9315),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10757),
            .sr(N__10675));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_11_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_11_9_2  (
            .in0(N__9273),
            .in1(N__11037),
            .in2(_gnd_net_),
            .in3(N__9888),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10757),
            .sr(N__10675));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_10_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_10_2  (
            .in0(N__7863),
            .in1(N__11876),
            .in2(N__9801),
            .in3(N__7984),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_11_10_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_11_10_5  (
            .in0(N__8895),
            .in1(N__8850),
            .in2(_gnd_net_),
            .in3(N__9004),
            .lcout(\U712_CHIP_RAM.N_450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_10_6  (
            .in0(N__8058),
            .in1(N__8040),
            .in2(_gnd_net_),
            .in3(N__7983),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_10_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_10_7  (
            .in0(N__11875),
            .in1(N__7985),
            .in2(N__8034),
            .in3(N__9231),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_11_4  (
            .in0(N__8025),
            .in1(N__7839),
            .in2(_gnd_net_),
            .in3(N__7982),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7857),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10198),
            .ce(N__7833),
            .sr(N__10656));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_12_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_12_1  (
            .in0(N__7812),
            .in1(N__7772),
            .in2(N__11043),
            .in3(N__7791),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10201),
            .ce(),
            .sr(N__10652));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_12_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_12_2  (
            .in0(N__7757),
            .in1(N__7737),
            .in2(_gnd_net_),
            .in3(N__7701),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_12_3 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_11_12_3  (
            .in0(N__7667),
            .in1(N__11111),
            .in2(N__7683),
            .in3(N__8381),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10201),
            .ce(),
            .sr(N__10652));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_5  (
            .in0(N__8399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8380),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.PRnW_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.PRnW_LC_11_12_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.PRnW_LC_11_12_7 .LUT_INIT=16'b1111110100110001;
    LogicCell40 \U712_REG_SM.PRnW_LC_11_12_7  (
            .in0(N__8595),
            .in1(N__8165),
            .in2(N__8532),
            .in3(N__8234),
            .lcout(PRnW_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10201),
            .ce(),
            .sr(N__10652));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_11_13_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__9468),
            .in2(_gnd_net_),
            .in3(N__8218),
            .lcout(\U712_REG_SM.N_351 ),
            .ltout(\U712_REG_SM.N_351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_11_13_2 .LUT_INIT=16'b1111111110110001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_11_13_2  (
            .in0(N__8525),
            .in1(N__8202),
            .in2(N__8169),
            .in3(N__9444),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_13_5 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_13_5  (
            .in0(N__9648),
            .in1(N__10026),
            .in2(N__10450),
            .in3(N__10059),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10207),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__11859),
            .in2(_gnd_net_),
            .in3(N__8088),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_7 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_7  (
            .in0(N__8139),
            .in1(N__8118),
            .in2(N__8091),
            .in3(N__10394),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10207),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_RNITKK4_1_LC_11_14_6.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_11_14_6.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_11_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_11_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8974),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_11_15_0  (
            .in0(N__8589),
            .in1(N__8428),
            .in2(_gnd_net_),
            .in3(N__8483),
            .lcout(\U712_REG_SM.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__10479),
            .in2(_gnd_net_),
            .in3(N__8562),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10216),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_15_3  (
            .in0(N__8429),
            .in1(N__10478),
            .in2(_gnd_net_),
            .in3(N__9501),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10216),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__8427),
            .in2(_gnd_net_),
            .in3(N__9500),
            .lcout(\U712_REG_SM.N_588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_15_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_2_LC_11_15_6  (
            .in0(N__8735),
            .in1(N__9521),
            .in2(_gnd_net_),
            .in3(N__9472),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_11_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_11_16_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_11_16_1  (
            .in0(N__8543),
            .in1(N__8524),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(\U712_REG_SM.N_395 ),
            .ltout(\U712_REG_SM.N_395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_16_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_16_2 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__8479),
            .in2(N__8451),
            .in3(N__9447),
            .lcout(),
            .ltout(\U712_REG_SM.N_439_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_11_16_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_16_3 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_11_16_3  (
            .in0(N__10504),
            .in1(N__8822),
            .in2(N__8448),
            .in3(N__8445),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10222),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_16_7 .LUT_INIT=16'b1000000010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_11_16_7  (
            .in0(N__10505),
            .in1(N__9502),
            .in2(N__8433),
            .in3(N__8439),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10222),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_17_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_11_17_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__10718),
            .in2(_gnd_net_),
            .in3(N__8761),
            .lcout(\U712_REG_SM.N_131_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_17_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_11_17_3  (
            .in0(N__10508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8724),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10227),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_17_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_11_17_7  (
            .in0(N__10507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8739),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10227),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_7_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8718),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10186),
            .ce(),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_6  (
            .in0(N__11036),
            .in1(N__9750),
            .in2(_gnd_net_),
            .in3(N__9192),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10762),
            .sr(N__10672));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_9_0  (
            .in0(N__9222),
            .in1(N__11006),
            .in2(_gnd_net_),
            .in3(N__9187),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10760),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_9_2  (
            .in0(N__9301),
            .in1(N__11014),
            .in2(_gnd_net_),
            .in3(N__10861),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10760),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_9_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_9_3  (
            .in0(N__9789),
            .in1(_gnd_net_),
            .in2(N__11034),
            .in3(N__9957),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10760),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_9_5  (
            .in0(N__11010),
            .in1(N__9887),
            .in2(_gnd_net_),
            .in3(N__9843),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10760),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_9_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_9_7  (
            .in0(N__9272),
            .in1(_gnd_net_),
            .in2(N__11035),
            .in3(N__9300),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10760),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_10_2  (
            .in0(N__9742),
            .in1(N__11001),
            .in2(_gnd_net_),
            .in3(N__9787),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10758),
            .sr(N__10653));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_10_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_10_3  (
            .in0(N__9788),
            .in1(_gnd_net_),
            .in2(N__11033),
            .in3(N__9956),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10758),
            .sr(N__10653));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_12_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_12_11_0  (
            .in0(N__9044),
            .in1(N__9068),
            .in2(N__8941),
            .in3(N__9102),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_196_i_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_196_i_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_196_i_LC_12_12_0 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \U712_BUFFERS.N_196_i_LC_12_12_0  (
            .in0(N__11277),
            .in1(N__11351),
            .in2(N__8840),
            .in3(N__11886),
            .lcout(N_196_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_12_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_12_12_1  (
            .in0(N__10351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9111),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_12_12_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_12_12_2  (
            .in0(N__8933),
            .in1(N__10348),
            .in2(N__9033),
            .in3(N__9011),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_12_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_12_3  (
            .in0(N__8781),
            .in1(N__9110),
            .in2(_gnd_net_),
            .in3(N__8931),
            .lcout(\U712_CHIP_RAM.N_492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_12_12_4 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_12_12_4  (
            .in0(N__8932),
            .in1(N__10347),
            .in2(N__9057),
            .in3(N__9010),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_12_12_5 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_12_12_5  (
            .in0(N__10346),
            .in1(N__9075),
            .in2(N__9012),
            .in3(N__8934),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_12_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__10350),
            .in2(_gnd_net_),
            .in3(N__9693),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_12_12_7  (
            .in0(N__10349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9018),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10195),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_12_13_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_12_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__9101),
            .in2(N__9090),
            .in3(N__9089),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_12_13_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_12_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__9069),
            .in2(_gnd_net_),
            .in3(N__9048),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_12_13_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_12_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__9045),
            .in2(_gnd_net_),
            .in3(N__9024),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_12_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__8888),
            .in2(_gnd_net_),
            .in3(N__9021),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_13_5 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_12_13_5  (
            .in0(N__11350),
            .in1(N__10353),
            .in2(_gnd_net_),
            .in3(N__11267),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10199),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_12_13_6 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_12_13_6  (
            .in0(N__10352),
            .in1(N__9006),
            .in2(N__8945),
            .in3(N__8901),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10199),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_14_6 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_12_14_6  (
            .in0(N__9537),
            .in1(N__9473),
            .in2(N__9531),
            .in3(N__9510),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10203),
            .ce(),
            .sr(N__10646));
    defparam \U712_REG_SM.ASn_ess_LC_12_17_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_12_17_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_12_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9445),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10217),
            .ce(N__9357),
            .sr(N__10642));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10365),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0  (
            .in0(N__9188),
            .in1(N__11015),
            .in2(_gnd_net_),
            .in3(N__9749),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(N__10765),
            .sr(N__10684));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_2  (
            .in0(N__9880),
            .in1(N__11005),
            .in2(_gnd_net_),
            .in3(N__9271),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(N__10763),
            .sr(N__10676));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_3  (
            .in0(N__9314),
            .in1(N__10994),
            .in2(_gnd_net_),
            .in3(N__9253),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10761),
            .sr(N__10667));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_3  (
            .in0(N__9221),
            .in1(N__10980),
            .in2(_gnd_net_),
            .in3(N__9168),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10756),
            .sr(N__10657));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_5  (
            .in0(N__10981),
            .in1(N__9839),
            .in2(_gnd_net_),
            .in3(N__9948),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10756),
            .sr(N__10657));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_13_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_13_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__9678),
            .in2(_gnd_net_),
            .in3(N__9672),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_13_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__9549),
            .in2(_gnd_net_),
            .in3(N__9669),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_13_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_13_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__9576),
            .in2(_gnd_net_),
            .in3(N__9666),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_13_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_13_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__9588),
            .in2(_gnd_net_),
            .in3(N__9663),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_13_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_13_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__9563),
            .in2(_gnd_net_),
            .in3(N__9660),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_13_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__10038),
            .in2(_gnd_net_),
            .in3(N__9657),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_13_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_13_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__10050),
            .in2(_gnd_net_),
            .in3(N__9654),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_13_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_13_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__9644),
            .in2(_gnd_net_),
            .in3(N__9651),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9623),
            .ce(),
            .sr(N__9600));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_13_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_13_3  (
            .in0(N__9587),
            .in1(N__9575),
            .in2(N__9564),
            .in3(N__9548),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_13_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__10049),
            .in2(_gnd_net_),
            .in3(N__10037),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_14_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10017),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10192),
            .ce(),
            .sr(N__10689));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_3  (
            .in0(N__9955),
            .in1(N__11020),
            .in2(_gnd_net_),
            .in3(N__9838),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(N__10766),
            .sr(N__10685));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_6  (
            .in0(N__9871),
            .in1(N__10982),
            .in2(_gnd_net_),
            .in3(N__9837),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10764),
            .sr(N__10677));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_11_2  (
            .in0(N__10918),
            .in1(N__9773),
            .in2(_gnd_net_),
            .in3(N__9728),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10788),
            .ce(N__10759),
            .sr(N__10668));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_14_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_14_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__10375),
            .in2(_gnd_net_),
            .in3(N__9684),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10208),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_14_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_14_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_14_12_5  (
            .in0(N__10374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10242),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10208),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_13_6  (
            .in0(N__11480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11536),
            .lcout(\U712_BYTE_ENABLE.N_331_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_412_i_LC_14_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_412_i_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_412_i_LC_14_20_1 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_BYTE_ENABLE.N_412_i_LC_14_20_1  (
            .in0(N__11711),
            .in1(N__11669),
            .in2(N__11551),
            .in3(N__11470),
            .lcout(N_412_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_9_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_9_1  (
            .in0(N__10550),
            .in1(N__11019),
            .in2(_gnd_net_),
            .in3(N__10854),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10786),
            .ce(N__10767),
            .sr(N__10690));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_10_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_15_10_5  (
            .in0(N__10551),
            .in1(N__10373),
            .in2(_gnd_net_),
            .in3(N__10527),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10202),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__10285),
            .in2(_gnd_net_),
            .in3(N__10248),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10209),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_15_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_15_12_4 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_15_12_4  (
            .in0(N__11727),
            .in1(N__11670),
            .in2(N__11904),
            .in3(N__11921),
            .lcout(\U712_BYTE_ENABLE.N_452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_15_12_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_15_12_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_15_12_7  (
            .in0(N__11126),
            .in1(N__11272),
            .in2(_gnd_net_),
            .in3(N__11189),
            .lcout(\U712_BYTE_ENABLE.N_467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_15_13_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_15_13_1 .LUT_INIT=16'b1010010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_15_13_1  (
            .in0(N__11481),
            .in1(_gnd_net_),
            .in2(N__11589),
            .in3(N__11907),
            .lcout(\U712_BYTE_ENABLE.N_455 ),
            .ltout(\U712_BYTE_ENABLE.N_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_38_i_LC_15_13_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_38_i_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_38_i_LC_15_13_2 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_BYTE_ENABLE.N_38_i_LC_15_13_2  (
            .in0(N__11725),
            .in1(N__10092),
            .in2(N__10086),
            .in3(N__11958),
            .lcout(N_38_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_15_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_15_13_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_15_13_4  (
            .in0(N__11906),
            .in1(N__11665),
            .in2(_gnd_net_),
            .in3(N__11583),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_209_i_LC_15_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_209_i_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_209_i_LC_15_13_5 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \U712_BYTE_ENABLE.N_209_i_LC_15_13_5  (
            .in0(N__11952),
            .in1(N__11724),
            .in2(N__11946),
            .in3(N__11064),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_7 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_7  (
            .in0(N__11664),
            .in1(N__11726),
            .in2(N__11922),
            .in3(N__11905),
            .lcout(\U712_BYTE_ENABLE.N_464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_15_19_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_i_LC_15_19_3 .LUT_INIT=16'b0000110111000000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_i_LC_15_19_3  (
            .in0(N__11661),
            .in1(N__11689),
            .in2(N__11582),
            .in3(N__11473),
            .lcout(N_205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_411_i_LC_15_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_411_i_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_411_i_LC_15_20_5 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_411_i_LC_15_20_5  (
            .in0(N__11713),
            .in1(N__11663),
            .in2(N__11588),
            .in3(N__11472),
            .lcout(N_411_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_15_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_15_20_7 .LUT_INIT=16'b0000011101010000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_15_20_7  (
            .in0(N__11712),
            .in1(N__11662),
            .in2(N__11587),
            .in3(N__11471),
            .lcout(N_213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_40_i_LC_16_12_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_40_i_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_40_i_LC_16_12_0 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \U712_BYTE_ENABLE.N_40_i_LC_16_12_0  (
            .in0(N__11141),
            .in1(N__11388),
            .in2(N__11198),
            .in3(N__11339),
            .lcout(N_40_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_208_i_LC_16_12_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_208_i_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_208_i_LC_16_12_3 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \U712_BYTE_ENABLE.N_208_i_LC_16_12_3  (
            .in0(N__11140),
            .in1(N__11364),
            .in2(N__11349),
            .in3(N__11190),
            .lcout(N_208_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_16_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_16_13_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_16_13_5  (
            .in0(N__11260),
            .in1(N__11194),
            .in2(_gnd_net_),
            .in3(N__11139),
            .lcout(\U712_BYTE_ENABLE.N_456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

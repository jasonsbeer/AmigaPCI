module U109_PCI_STATE_MACHINE (

    output PCICYCLEn, ADLATCH, ALATCH, PCI_DIR, AD_ENn

);

//DISABLE THE ADDRESS BUFFERS FOR NOW.

//ADDRESS DATA IS PASSED THROUGH LIVE DURING THE ADDRESS PHASE OF CPU DRIVEN CYCLES.
//FOR PCI DRIVEN DMA CYCLES, THE ADDRESS IS LATCHED DURING THE ADDRESS PHASE AND
//DRIVEN ON THE ADDRESS BUS OF THE AMIGAPCI.

assign PCICYCLEn = 1; //Disables the A <-> AD address buffers.
assign ADLATCH = 0;
assign ALATCH = 0; //WE DON'T ACTUALLY NEED THIS, BUT ITS THERE.
assign PCI_DIR = 0;
assign AD_ENn = 1;


endmodule

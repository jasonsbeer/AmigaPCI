// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 23 2024 16:31:47

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    A,
    TICK50,
    nROMEN,
    nCIACS1,
    TICK60,
    CLKCIA,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    TSn,
    nBUFEN,
    nREGSPACE,
    nRAMSPACE,
    RESETn,
    OVL,
    TACKn,
    nCIACS0,
    PORTSIZE);

    input [31:1] A;
    output TICK50;
    output nROMEN;
    output nCIACS1;
    output TICK60;
    output CLKCIA;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    input TSn;
    output nBUFEN;
    output nREGSPACE;
    output nRAMSPACE;
    input RESETn;
    input OVL;
    inout TACKn;
    output nCIACS0;
    output PORTSIZE;

    wire N__6073;
    wire N__6072;
    wire N__6071;
    wire N__6063;
    wire N__6062;
    wire N__6061;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6043;
    wire N__6042;
    wire N__6041;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6016;
    wire N__6015;
    wire N__6014;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__5998;
    wire N__5997;
    wire N__5996;
    wire N__5989;
    wire N__5988;
    wire N__5987;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5962;
    wire N__5961;
    wire N__5960;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5944;
    wire N__5943;
    wire N__5942;
    wire N__5935;
    wire N__5934;
    wire N__5933;
    wire N__5926;
    wire N__5925;
    wire N__5924;
    wire N__5917;
    wire N__5916;
    wire N__5915;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5899;
    wire N__5898;
    wire N__5897;
    wire N__5890;
    wire N__5889;
    wire N__5888;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5845;
    wire N__5844;
    wire N__5843;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5827;
    wire N__5826;
    wire N__5825;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5809;
    wire N__5808;
    wire N__5807;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5791;
    wire N__5790;
    wire N__5789;
    wire N__5782;
    wire N__5781;
    wire N__5780;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5764;
    wire N__5763;
    wire N__5762;
    wire N__5745;
    wire N__5742;
    wire N__5741;
    wire N__5740;
    wire N__5739;
    wire N__5736;
    wire N__5731;
    wire N__5728;
    wire N__5721;
    wire N__5720;
    wire N__5719;
    wire N__5718;
    wire N__5713;
    wire N__5708;
    wire N__5703;
    wire N__5700;
    wire N__5699;
    wire N__5698;
    wire N__5697;
    wire N__5692;
    wire N__5687;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5677;
    wire N__5674;
    wire N__5667;
    wire N__5662;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5648;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5627;
    wire N__5620;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5603;
    wire N__5602;
    wire N__5601;
    wire N__5600;
    wire N__5599;
    wire N__5598;
    wire N__5593;
    wire N__5588;
    wire N__5581;
    wire N__5574;
    wire N__5573;
    wire N__5572;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5482;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5476;
    wire N__5475;
    wire N__5474;
    wire N__5473;
    wire N__5472;
    wire N__5471;
    wire N__5470;
    wire N__5469;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5462;
    wire N__5459;
    wire N__5448;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5429;
    wire N__5420;
    wire N__5411;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5403;
    wire N__5400;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5366;
    wire N__5363;
    wire N__5358;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5277;
    wire N__5276;
    wire N__5275;
    wire N__5274;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5270;
    wire N__5269;
    wire N__5262;
    wire N__5255;
    wire N__5248;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5224;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5197;
    wire N__5192;
    wire N__5187;
    wire N__5178;
    wire N__5177;
    wire N__5176;
    wire N__5175;
    wire N__5174;
    wire N__5173;
    wire N__5172;
    wire N__5171;
    wire N__5166;
    wire N__5159;
    wire N__5152;
    wire N__5149;
    wire N__5142;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5122;
    wire N__5121;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4956;
    wire N__4955;
    wire N__4950;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4938;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4914;
    wire N__4911;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4899;
    wire N__4896;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4884;
    wire N__4881;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4869;
    wire N__4866;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4806;
    wire N__4803;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4773;
    wire N__4772;
    wire N__4771;
    wire N__4770;
    wire N__4769;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4746;
    wire N__4745;
    wire N__4744;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4732;
    wire N__4725;
    wire N__4724;
    wire N__4721;
    wire N__4720;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4705;
    wire N__4698;
    wire N__4697;
    wire N__4696;
    wire N__4693;
    wire N__4688;
    wire N__4683;
    wire N__4682;
    wire N__4681;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4659;
    wire N__4658;
    wire N__4657;
    wire N__4656;
    wire N__4655;
    wire N__4654;
    wire N__4653;
    wire N__4650;
    wire N__4645;
    wire N__4642;
    wire N__4633;
    wire N__4626;
    wire N__4623;
    wire N__4622;
    wire N__4621;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4607;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4591;
    wire N__4584;
    wire N__4583;
    wire N__4582;
    wire N__4579;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4567;
    wire N__4560;
    wire N__4559;
    wire N__4554;
    wire N__4551;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4526;
    wire N__4525;
    wire N__4524;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4454;
    wire N__4449;
    wire N__4448;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4300;
    wire N__4295;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4277;
    wire N__4276;
    wire N__4271;
    wire N__4268;
    wire N__4263;
    wire N__4262;
    wire N__4259;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4253;
    wire N__4246;
    wire N__4243;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4199;
    wire N__4198;
    wire N__4195;
    wire N__4190;
    wire N__4185;
    wire N__4184;
    wire N__4183;
    wire N__4178;
    wire N__4175;
    wire N__4170;
    wire N__4167;
    wire N__4166;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4158;
    wire N__4151;
    wire N__4146;
    wire N__4145;
    wire N__4142;
    wire N__4141;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4103;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4088;
    wire N__4087;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4066;
    wire N__4063;
    wire N__4056;
    wire N__4055;
    wire N__4052;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4035;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4023;
    wire N__4020;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3996;
    wire N__3995;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3987;
    wire N__3986;
    wire N__3985;
    wire N__3982;
    wire N__3981;
    wire N__3976;
    wire N__3973;
    wire N__3964;
    wire N__3961;
    wire N__3954;
    wire N__3953;
    wire N__3952;
    wire N__3951;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3945;
    wire N__3940;
    wire N__3937;
    wire N__3930;
    wire N__3921;
    wire N__3920;
    wire N__3919;
    wire N__3918;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3910;
    wire N__3909;
    wire N__3906;
    wire N__3901;
    wire N__3896;
    wire N__3891;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3816;
    wire N__3815;
    wire N__3814;
    wire N__3807;
    wire N__3804;
    wire N__3803;
    wire N__3802;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3695;
    wire N__3692;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3653;
    wire N__3652;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3641;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3612;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3546;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3534;
    wire N__3531;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3519;
    wire N__3516;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3504;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3474;
    wire N__3473;
    wire N__3472;
    wire N__3471;
    wire N__3468;
    wire N__3461;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3405;
    wire N__3402;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3309;
    wire N__3306;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3237;
    wire N__3234;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3200;
    wire N__3199;
    wire N__3198;
    wire N__3189;
    wire N__3186;
    wire N__3185;
    wire N__3184;
    wire N__3183;
    wire N__3180;
    wire N__3179;
    wire N__3174;
    wire N__3167;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3100;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3069;
    wire N__3068;
    wire N__3067;
    wire N__3064;
    wire N__3059;
    wire N__3054;
    wire N__3053;
    wire N__3052;
    wire N__3051;
    wire N__3048;
    wire N__3047;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3027;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3015;
    wire N__3012;
    wire N__3011;
    wire N__3008;
    wire N__3007;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2995;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2934;
    wire N__2931;
    wire N__2930;
    wire N__2929;
    wire N__2928;
    wire N__2925;
    wire N__2924;
    wire N__2923;
    wire N__2918;
    wire N__2915;
    wire N__2910;
    wire N__2907;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2840;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2822;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2801;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2774;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2756;
    wire N__2753;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2729;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2684;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2674;
    wire N__2671;
    wire N__2668;
    wire N__2665;
    wire N__2662;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2648;
    wire N__2647;
    wire N__2646;
    wire N__2641;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2597;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2526;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2508;
    wire N__2505;
    wire N__2504;
    wire N__2503;
    wire N__2500;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2459;
    wire N__2458;
    wire N__2455;
    wire N__2450;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2424;
    wire N__2421;
    wire N__2418;
    wire N__2415;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2397;
    wire N__2394;
    wire N__2391;
    wire N__2390;
    wire N__2389;
    wire N__2388;
    wire N__2387;
    wire N__2386;
    wire N__2385;
    wire N__2384;
    wire N__2383;
    wire N__2364;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_16;
    wire A_c_18;
    wire \U409_CIA.g0Z0Z_11 ;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.HIROM_0_cascade_ ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.HIROM_0 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire A_c_25;
    wire \U409_CIA.g0Z0Z_2_cascade_ ;
    wire A_c_30;
    wire A_c_28;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire A_c_24;
    wire A_c_26;
    wire A_c_31;
    wire A_c_27;
    wire \U409_CIA.g0Z0Z_10 ;
    wire A_c_22;
    wire A_c_21;
    wire \U409_CIA.g0Z0Z_8 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire PORTSIZE_0_i;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ;
    wire A_c_23;
    wire U409_ADDRESS_DECODE_un1_nREGSPACE_i;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_bm_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_am ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_97 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_ADDRESS_DECODE.HIROMZ0 ;
    wire U409_ADDRESS_DECODE_un1_ROMEN_0;
    wire U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_;
    wire ROMENm_i;
    wire \U409_TICK.TICK603_11_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_8 ;
    wire bfn_10_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_10_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.RESETn_c_i ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ;
    wire TSn_c;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_nCIACS1_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_nCIACS0_i;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire CIA_ENABLEm;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire CLKCIA_c;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ;
    wire U409_ADDRESS_DECODE_un1_nRAMSPACE_i;
    wire CONSTANT_ONE_NET;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_12_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_12_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire CLK6_c_g;
    wire bfn_12_9_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire CLK28_IN_c_g;
    wire TACK_EN_i;
    wire N_353_i;
    wire TACKn_in;
    wire nBUFEN_c;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__3654),
            .RESETB(N__4362),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6071),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6073),
            .DIN(N__6072),
            .DOUT(N__6071),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6073),
            .PADOUT(N__6072),
            .PADIN(N__6071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6061),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6063),
            .DIN(N__6062),
            .DOUT(N__6061),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6063),
            .PADOUT(N__6062),
            .PADIN(N__6061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6052),
            .DIN(N__6051),
            .DOUT(N__6050),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6052),
            .PADOUT(N__6051),
            .PADIN(N__6050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4323),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6043),
            .DIN(N__6042),
            .DOUT(N__6041),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6043),
            .PADOUT(N__6042),
            .PADIN(N__6041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6034),
            .DIN(N__6033),
            .DOUT(N__6032),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6034),
            .PADOUT(N__6033),
            .PADIN(N__6032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS0_obuf_iopad (
            .OE(N__6025),
            .DIN(N__6024),
            .DOUT(N__6023),
            .PACKAGEPIN(nCIACS0));
    defparam nCIACS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS0_obuf_preio (
            .PADOEN(N__6025),
            .PADOUT(N__6024),
            .PADIN(N__6023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3720),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS1_obuf_iopad (
            .OE(N__6016),
            .DIN(N__6015),
            .DOUT(N__6014),
            .PACKAGEPIN(nCIACS1));
    defparam nCIACS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS1_obuf_preio (
            .PADOEN(N__6016),
            .PADOUT(N__6015),
            .PADIN(N__6014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6007),
            .DIN(N__6006),
            .DOUT(N__6005),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6007),
            .PADOUT(N__6006),
            .PADIN(N__6005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__5998),
            .DIN(N__5997),
            .DOUT(N__5996),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__5998),
            .PADOUT(N__5997),
            .PADIN(N__5996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__5989),
            .DIN(N__5988),
            .DOUT(N__5987),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__5989),
            .PADOUT(N__5988),
            .PADIN(N__5987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__5980),
            .DIN(N__5979),
            .DOUT(N__5978),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__5980),
            .PADOUT(N__5979),
            .PADIN(N__5978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5547),
            .DIN0(TACKn_in),
            .DOUT0(N__3846),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__5971),
            .DIN(N__5970),
            .DOUT(N__5969),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__5971),
            .PADOUT(N__5970),
            .PADIN(N__5969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__5962),
            .DIN(N__5961),
            .DOUT(N__5960),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__5962),
            .PADOUT(N__5961),
            .PADIN(N__5960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__5953),
            .DIN(N__5952),
            .DOUT(N__5951),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__5953),
            .PADOUT(N__5952),
            .PADIN(N__5951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2973),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nRAMSPACE_obuf_iopad (
            .OE(N__5944),
            .DIN(N__5943),
            .DOUT(N__5942),
            .PACKAGEPIN(nRAMSPACE));
    defparam nRAMSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nRAMSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nRAMSPACE_obuf_preio (
            .PADOEN(N__5944),
            .PADOUT(N__5943),
            .PADIN(N__5942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nROMEN_obuf_iopad (
            .OE(N__5935),
            .DIN(N__5934),
            .DOUT(N__5933),
            .PACKAGEPIN(nROMEN));
    defparam nROMEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nROMEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nROMEN_obuf_preio (
            .PADOEN(N__5935),
            .PADOUT(N__5934),
            .PADIN(N__5933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3141),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__5926),
            .DIN(N__5925),
            .DOUT(N__5924),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__5926),
            .PADOUT(N__5925),
            .PADIN(N__5924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__5917),
            .DIN(N__5916),
            .DOUT(N__5915),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__5917),
            .PADOUT(N__5916),
            .PADIN(N__5915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nBUFEN_obuf_iopad (
            .OE(N__5908),
            .DIN(N__5907),
            .DOUT(N__5906),
            .PACKAGEPIN(nBUFEN));
    defparam nBUFEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nBUFEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nBUFEN_obuf_preio (
            .PADOEN(N__5908),
            .PADOUT(N__5907),
            .PADIN(N__5906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5511),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__5899),
            .DIN(N__5898),
            .DOUT(N__5897),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__5899),
            .PADOUT(N__5898),
            .PADIN(N__5897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__5890),
            .DIN(N__5889),
            .DOUT(N__5888),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__5890),
            .PADOUT(N__5889),
            .PADIN(N__5888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__5881),
            .DIN(N__5880),
            .DOUT(N__5879),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__5881),
            .PADOUT(N__5880),
            .PADIN(N__5879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__5872),
            .DIN(N__5871),
            .DOUT(N__5870),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__5872),
            .PADOUT(N__5871),
            .PADIN(N__5870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__5863),
            .DIN(N__5862),
            .DOUT(N__5861),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__5863),
            .PADOUT(N__5862),
            .PADIN(N__5861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__5854),
            .DIN(N__5853),
            .DOUT(N__5852),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__5854),
            .PADOUT(N__5853),
            .PADIN(N__5852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__5845),
            .DIN(N__5844),
            .DOUT(N__5843),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__5845),
            .PADOUT(N__5844),
            .PADIN(N__5843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nREGSPACE_obuf_iopad (
            .OE(N__5836),
            .DIN(N__5835),
            .DOUT(N__5834),
            .PACKAGEPIN(nREGSPACE));
    defparam nREGSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nREGSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nREGSPACE_obuf_preio (
            .PADOEN(N__5836),
            .PADOUT(N__5835),
            .PADIN(N__5834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__5827),
            .DIN(N__5826),
            .DOUT(N__5825),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__5827),
            .PADOUT(N__5826),
            .PADIN(N__5825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__5818),
            .DIN(N__5817),
            .DOUT(N__5816),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__5818),
            .PADOUT(N__5817),
            .PADIN(N__5816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__5809),
            .DIN(N__5808),
            .DOUT(N__5807),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__5809),
            .PADOUT(N__5808),
            .PADIN(N__5807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__5800),
            .DIN(N__5799),
            .DOUT(N__5798),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__5800),
            .PADOUT(N__5799),
            .PADIN(N__5798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__5791),
            .DIN(N__5790),
            .DOUT(N__5789),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__5791),
            .PADOUT(N__5790),
            .PADIN(N__5789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__5782),
            .DIN(N__5781),
            .DOUT(N__5780),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__5782),
            .PADOUT(N__5781),
            .PADIN(N__5780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__5773),
            .DIN(N__5772),
            .DOUT(N__5771),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__5773),
            .PADOUT(N__5772),
            .PADIN(N__5771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3282),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__5764),
            .DIN(N__5763),
            .DOUT(N__5762),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__5764),
            .PADOUT(N__5763),
            .PADIN(N__5762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1332 (
            .O(N__5745),
            .I(N__5742));
    InMux I__1331 (
            .O(N__5742),
            .I(N__5736));
    InMux I__1330 (
            .O(N__5741),
            .I(N__5731));
    InMux I__1329 (
            .O(N__5740),
            .I(N__5731));
    InMux I__1328 (
            .O(N__5739),
            .I(N__5728));
    LocalMux I__1327 (
            .O(N__5736),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1326 (
            .O(N__5731),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1325 (
            .O(N__5728),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1324 (
            .O(N__5721),
            .I(N__5713));
    InMux I__1323 (
            .O(N__5720),
            .I(N__5713));
    InMux I__1322 (
            .O(N__5719),
            .I(N__5708));
    InMux I__1321 (
            .O(N__5718),
            .I(N__5708));
    LocalMux I__1320 (
            .O(N__5713),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1319 (
            .O(N__5708),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__1318 (
            .O(N__5703),
            .I(N__5700));
    InMux I__1317 (
            .O(N__5700),
            .I(N__5692));
    InMux I__1316 (
            .O(N__5699),
            .I(N__5692));
    InMux I__1315 (
            .O(N__5698),
            .I(N__5687));
    InMux I__1314 (
            .O(N__5697),
            .I(N__5687));
    LocalMux I__1313 (
            .O(N__5692),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1312 (
            .O(N__5687),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1311 (
            .O(N__5682),
            .I(N__5674));
    InMux I__1310 (
            .O(N__5681),
            .I(N__5667));
    InMux I__1309 (
            .O(N__5680),
            .I(N__5667));
    InMux I__1308 (
            .O(N__5679),
            .I(N__5667));
    InMux I__1307 (
            .O(N__5678),
            .I(N__5662));
    InMux I__1306 (
            .O(N__5677),
            .I(N__5662));
    LocalMux I__1305 (
            .O(N__5674),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1304 (
            .O(N__5667),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1303 (
            .O(N__5662),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__1302 (
            .O(N__5655),
            .I(N__5652));
    LocalMux I__1301 (
            .O(N__5652),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    CascadeMux I__1300 (
            .O(N__5649),
            .I(N__5639));
    InMux I__1299 (
            .O(N__5648),
            .I(N__5636));
    InMux I__1298 (
            .O(N__5647),
            .I(N__5627));
    InMux I__1297 (
            .O(N__5646),
            .I(N__5627));
    InMux I__1296 (
            .O(N__5645),
            .I(N__5627));
    InMux I__1295 (
            .O(N__5644),
            .I(N__5627));
    InMux I__1294 (
            .O(N__5643),
            .I(N__5620));
    InMux I__1293 (
            .O(N__5642),
            .I(N__5620));
    InMux I__1292 (
            .O(N__5639),
            .I(N__5620));
    LocalMux I__1291 (
            .O(N__5636),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1290 (
            .O(N__5627),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1289 (
            .O(N__5620),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__1288 (
            .O(N__5613),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ));
    InMux I__1287 (
            .O(N__5610),
            .I(N__5607));
    LocalMux I__1286 (
            .O(N__5607),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    InMux I__1285 (
            .O(N__5604),
            .I(N__5593));
    InMux I__1284 (
            .O(N__5603),
            .I(N__5593));
    InMux I__1283 (
            .O(N__5602),
            .I(N__5588));
    InMux I__1282 (
            .O(N__5601),
            .I(N__5588));
    InMux I__1281 (
            .O(N__5600),
            .I(N__5581));
    InMux I__1280 (
            .O(N__5599),
            .I(N__5581));
    InMux I__1279 (
            .O(N__5598),
            .I(N__5581));
    LocalMux I__1278 (
            .O(N__5593),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1277 (
            .O(N__5588),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1276 (
            .O(N__5581),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    ClkMux I__1275 (
            .O(N__5574),
            .I(N__5565));
    ClkMux I__1274 (
            .O(N__5573),
            .I(N__5565));
    ClkMux I__1273 (
            .O(N__5572),
            .I(N__5565));
    GlobalMux I__1272 (
            .O(N__5565),
            .I(N__5562));
    gio2CtrlBuf I__1271 (
            .O(N__5562),
            .I(CLK28_IN_c_g));
    InMux I__1270 (
            .O(N__5559),
            .I(N__5556));
    LocalMux I__1269 (
            .O(N__5556),
            .I(N__5553));
    Span4Mux_v I__1268 (
            .O(N__5553),
            .I(N__5550));
    Odrv4 I__1267 (
            .O(N__5550),
            .I(TACK_EN_i));
    IoInMux I__1266 (
            .O(N__5547),
            .I(N__5544));
    LocalMux I__1265 (
            .O(N__5544),
            .I(N__5541));
    Span12Mux_s2_v I__1264 (
            .O(N__5541),
            .I(N__5538));
    Span12Mux_v I__1263 (
            .O(N__5538),
            .I(N__5535));
    Odrv12 I__1262 (
            .O(N__5535),
            .I(N_353_i));
    InMux I__1261 (
            .O(N__5532),
            .I(N__5529));
    LocalMux I__1260 (
            .O(N__5529),
            .I(N__5526));
    Span4Mux_v I__1259 (
            .O(N__5526),
            .I(N__5523));
    Sp12to4 I__1258 (
            .O(N__5523),
            .I(N__5520));
    Span12Mux_h I__1257 (
            .O(N__5520),
            .I(N__5517));
    Span12Mux_v I__1256 (
            .O(N__5517),
            .I(N__5514));
    Odrv12 I__1255 (
            .O(N__5514),
            .I(TACKn_in));
    IoInMux I__1254 (
            .O(N__5511),
            .I(N__5508));
    LocalMux I__1253 (
            .O(N__5508),
            .I(N__5505));
    Span12Mux_s9_v I__1252 (
            .O(N__5505),
            .I(N__5501));
    InMux I__1251 (
            .O(N__5504),
            .I(N__5498));
    Span12Mux_h I__1250 (
            .O(N__5501),
            .I(N__5495));
    LocalMux I__1249 (
            .O(N__5498),
            .I(N__5492));
    Odrv12 I__1248 (
            .O(N__5495),
            .I(nBUFEN_c));
    Odrv12 I__1247 (
            .O(N__5492),
            .I(nBUFEN_c));
    InMux I__1246 (
            .O(N__5487),
            .I(N__5482));
    CascadeMux I__1245 (
            .O(N__5486),
            .I(N__5476));
    CascadeMux I__1244 (
            .O(N__5485),
            .I(N__5463));
    LocalMux I__1243 (
            .O(N__5482),
            .I(N__5459));
    InMux I__1242 (
            .O(N__5481),
            .I(N__5448));
    InMux I__1241 (
            .O(N__5480),
            .I(N__5448));
    InMux I__1240 (
            .O(N__5479),
            .I(N__5448));
    InMux I__1239 (
            .O(N__5476),
            .I(N__5448));
    InMux I__1238 (
            .O(N__5475),
            .I(N__5448));
    InMux I__1237 (
            .O(N__5474),
            .I(N__5439));
    InMux I__1236 (
            .O(N__5473),
            .I(N__5439));
    InMux I__1235 (
            .O(N__5472),
            .I(N__5439));
    InMux I__1234 (
            .O(N__5471),
            .I(N__5439));
    InMux I__1233 (
            .O(N__5470),
            .I(N__5436));
    InMux I__1232 (
            .O(N__5469),
            .I(N__5433));
    InMux I__1231 (
            .O(N__5468),
            .I(N__5430));
    InMux I__1230 (
            .O(N__5467),
            .I(N__5420));
    InMux I__1229 (
            .O(N__5466),
            .I(N__5420));
    InMux I__1228 (
            .O(N__5463),
            .I(N__5420));
    InMux I__1227 (
            .O(N__5462),
            .I(N__5420));
    Span4Mux_v I__1226 (
            .O(N__5459),
            .I(N__5411));
    LocalMux I__1225 (
            .O(N__5448),
            .I(N__5411));
    LocalMux I__1224 (
            .O(N__5439),
            .I(N__5411));
    LocalMux I__1223 (
            .O(N__5436),
            .I(N__5411));
    LocalMux I__1222 (
            .O(N__5433),
            .I(N__5407));
    LocalMux I__1221 (
            .O(N__5430),
            .I(N__5404));
    InMux I__1220 (
            .O(N__5429),
            .I(N__5400));
    LocalMux I__1219 (
            .O(N__5420),
            .I(N__5395));
    Span4Mux_v I__1218 (
            .O(N__5411),
            .I(N__5395));
    InMux I__1217 (
            .O(N__5410),
            .I(N__5392));
    Span4Mux_v I__1216 (
            .O(N__5407),
            .I(N__5389));
    Span4Mux_v I__1215 (
            .O(N__5404),
            .I(N__5386));
    InMux I__1214 (
            .O(N__5403),
            .I(N__5383));
    LocalMux I__1213 (
            .O(N__5400),
            .I(N__5380));
    Span4Mux_h I__1212 (
            .O(N__5395),
            .I(N__5377));
    LocalMux I__1211 (
            .O(N__5392),
            .I(N__5374));
    Sp12to4 I__1210 (
            .O(N__5389),
            .I(N__5371));
    Span4Mux_h I__1209 (
            .O(N__5386),
            .I(N__5366));
    LocalMux I__1208 (
            .O(N__5383),
            .I(N__5366));
    Span4Mux_h I__1207 (
            .O(N__5380),
            .I(N__5363));
    Span4Mux_h I__1206 (
            .O(N__5377),
            .I(N__5358));
    Span4Mux_v I__1205 (
            .O(N__5374),
            .I(N__5358));
    Span12Mux_h I__1204 (
            .O(N__5371),
            .I(N__5351));
    Sp12to4 I__1203 (
            .O(N__5366),
            .I(N__5351));
    Sp12to4 I__1202 (
            .O(N__5363),
            .I(N__5351));
    Sp12to4 I__1201 (
            .O(N__5358),
            .I(N__5348));
    Span12Mux_v I__1200 (
            .O(N__5351),
            .I(N__5345));
    Span12Mux_h I__1199 (
            .O(N__5348),
            .I(N__5342));
    Span12Mux_h I__1198 (
            .O(N__5345),
            .I(N__5337));
    Span12Mux_v I__1197 (
            .O(N__5342),
            .I(N__5337));
    Odrv12 I__1196 (
            .O(N__5337),
            .I(RESETn_c));
    SRMux I__1195 (
            .O(N__5334),
            .I(N__5331));
    LocalMux I__1194 (
            .O(N__5331),
            .I(N__5328));
    Span4Mux_v I__1193 (
            .O(N__5328),
            .I(N__5323));
    SRMux I__1192 (
            .O(N__5327),
            .I(N__5320));
    SRMux I__1191 (
            .O(N__5326),
            .I(N__5317));
    Span4Mux_v I__1190 (
            .O(N__5323),
            .I(N__5310));
    LocalMux I__1189 (
            .O(N__5320),
            .I(N__5310));
    LocalMux I__1188 (
            .O(N__5317),
            .I(N__5310));
    Span4Mux_v I__1187 (
            .O(N__5310),
            .I(N__5307));
    Span4Mux_h I__1186 (
            .O(N__5307),
            .I(N__5304));
    Odrv4 I__1185 (
            .O(N__5304),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1184 (
            .O(N__5301),
            .I(N__5298));
    LocalMux I__1183 (
            .O(N__5298),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1182 (
            .O(N__5295),
            .I(N__5292));
    LocalMux I__1181 (
            .O(N__5292),
            .I(N__5289));
    Span4Mux_h I__1180 (
            .O(N__5289),
            .I(N__5285));
    InMux I__1179 (
            .O(N__5288),
            .I(N__5282));
    Odrv4 I__1178 (
            .O(N__5285),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1177 (
            .O(N__5282),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1176 (
            .O(N__5277),
            .I(N__5262));
    InMux I__1175 (
            .O(N__5276),
            .I(N__5262));
    InMux I__1174 (
            .O(N__5275),
            .I(N__5262));
    InMux I__1173 (
            .O(N__5274),
            .I(N__5255));
    InMux I__1172 (
            .O(N__5273),
            .I(N__5255));
    InMux I__1171 (
            .O(N__5272),
            .I(N__5255));
    InMux I__1170 (
            .O(N__5271),
            .I(N__5248));
    InMux I__1169 (
            .O(N__5270),
            .I(N__5248));
    InMux I__1168 (
            .O(N__5269),
            .I(N__5248));
    LocalMux I__1167 (
            .O(N__5262),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1166 (
            .O(N__5255),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1165 (
            .O(N__5248),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__1164 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__1163 (
            .O(N__5238),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    CascadeMux I__1162 (
            .O(N__5235),
            .I(N__5232));
    InMux I__1161 (
            .O(N__5232),
            .I(N__5224));
    CascadeMux I__1160 (
            .O(N__5231),
            .I(N__5220));
    CascadeMux I__1159 (
            .O(N__5230),
            .I(N__5217));
    CascadeMux I__1158 (
            .O(N__5229),
            .I(N__5214));
    CascadeMux I__1157 (
            .O(N__5228),
            .I(N__5211));
    CascadeMux I__1156 (
            .O(N__5227),
            .I(N__5208));
    LocalMux I__1155 (
            .O(N__5224),
            .I(N__5204));
    InMux I__1154 (
            .O(N__5223),
            .I(N__5197));
    InMux I__1153 (
            .O(N__5220),
            .I(N__5197));
    InMux I__1152 (
            .O(N__5217),
            .I(N__5197));
    InMux I__1151 (
            .O(N__5214),
            .I(N__5192));
    InMux I__1150 (
            .O(N__5211),
            .I(N__5192));
    InMux I__1149 (
            .O(N__5208),
            .I(N__5187));
    InMux I__1148 (
            .O(N__5207),
            .I(N__5187));
    Odrv4 I__1147 (
            .O(N__5204),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1146 (
            .O(N__5197),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1145 (
            .O(N__5192),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1144 (
            .O(N__5187),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__1143 (
            .O(N__5178),
            .I(N__5166));
    InMux I__1142 (
            .O(N__5177),
            .I(N__5166));
    InMux I__1141 (
            .O(N__5176),
            .I(N__5159));
    InMux I__1140 (
            .O(N__5175),
            .I(N__5159));
    InMux I__1139 (
            .O(N__5174),
            .I(N__5159));
    InMux I__1138 (
            .O(N__5173),
            .I(N__5152));
    InMux I__1137 (
            .O(N__5172),
            .I(N__5152));
    InMux I__1136 (
            .O(N__5171),
            .I(N__5152));
    LocalMux I__1135 (
            .O(N__5166),
            .I(N__5149));
    LocalMux I__1134 (
            .O(N__5159),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1133 (
            .O(N__5152),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__1132 (
            .O(N__5149),
            .I(\U409_TICK.TICK503_14 ));
    InMux I__1131 (
            .O(N__5142),
            .I(N__5138));
    InMux I__1130 (
            .O(N__5141),
            .I(N__5135));
    LocalMux I__1129 (
            .O(N__5138),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__1128 (
            .O(N__5135),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    ClkMux I__1127 (
            .O(N__5130),
            .I(N__5100));
    ClkMux I__1126 (
            .O(N__5129),
            .I(N__5100));
    ClkMux I__1125 (
            .O(N__5128),
            .I(N__5100));
    ClkMux I__1124 (
            .O(N__5127),
            .I(N__5100));
    ClkMux I__1123 (
            .O(N__5126),
            .I(N__5100));
    ClkMux I__1122 (
            .O(N__5125),
            .I(N__5100));
    ClkMux I__1121 (
            .O(N__5124),
            .I(N__5100));
    ClkMux I__1120 (
            .O(N__5123),
            .I(N__5100));
    ClkMux I__1119 (
            .O(N__5122),
            .I(N__5100));
    ClkMux I__1118 (
            .O(N__5121),
            .I(N__5100));
    GlobalMux I__1117 (
            .O(N__5100),
            .I(N__5097));
    gio2CtrlBuf I__1116 (
            .O(N__5097),
            .I(CLK6_c_g));
    InMux I__1115 (
            .O(N__5094),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1114 (
            .O(N__5091),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1113 (
            .O(N__5088),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1112 (
            .O(N__5085),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__1111 (
            .O(N__5082),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__1110 (
            .O(N__5079),
            .I(bfn_12_7_0_));
    InMux I__1109 (
            .O(N__5076),
            .I(N__5072));
    InMux I__1108 (
            .O(N__5075),
            .I(N__5069));
    LocalMux I__1107 (
            .O(N__5072),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1106 (
            .O(N__5069),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1105 (
            .O(N__5064),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    CascadeMux I__1104 (
            .O(N__5061),
            .I(N__5058));
    InMux I__1103 (
            .O(N__5058),
            .I(N__5054));
    InMux I__1102 (
            .O(N__5057),
            .I(N__5051));
    LocalMux I__1101 (
            .O(N__5054),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1100 (
            .O(N__5051),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__1099 (
            .O(N__5046),
            .I(N__5043));
    LocalMux I__1098 (
            .O(N__5043),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1097 (
            .O(N__5040),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__1096 (
            .O(N__5037),
            .I(N__5033));
    InMux I__1095 (
            .O(N__5036),
            .I(N__5030));
    LocalMux I__1094 (
            .O(N__5033),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1093 (
            .O(N__5030),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__1092 (
            .O(N__5025),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__1091 (
            .O(N__5022),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1090 (
            .O(N__5019),
            .I(N__5015));
    InMux I__1089 (
            .O(N__5018),
            .I(N__5012));
    LocalMux I__1088 (
            .O(N__5015),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1087 (
            .O(N__5012),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__1086 (
            .O(N__5007),
            .I(N__5004));
    LocalMux I__1085 (
            .O(N__5004),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1084 (
            .O(N__5001),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1083 (
            .O(N__4998),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1082 (
            .O(N__4995),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    CascadeMux I__1081 (
            .O(N__4992),
            .I(N__4988));
    InMux I__1080 (
            .O(N__4991),
            .I(N__4985));
    InMux I__1079 (
            .O(N__4988),
            .I(N__4982));
    LocalMux I__1078 (
            .O(N__4985),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__1077 (
            .O(N__4982),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    CascadeMux I__1076 (
            .O(N__4977),
            .I(N__4974));
    InMux I__1075 (
            .O(N__4974),
            .I(N__4971));
    LocalMux I__1074 (
            .O(N__4971),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1073 (
            .O(N__4968),
            .I(N__4964));
    InMux I__1072 (
            .O(N__4967),
            .I(N__4961));
    LocalMux I__1071 (
            .O(N__4964),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1070 (
            .O(N__4961),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__1069 (
            .O(N__4956),
            .I(N__4950));
    InMux I__1068 (
            .O(N__4955),
            .I(N__4950));
    LocalMux I__1067 (
            .O(N__4950),
            .I(N__4946));
    InMux I__1066 (
            .O(N__4949),
            .I(N__4943));
    Odrv4 I__1065 (
            .O(N__4946),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1064 (
            .O(N__4943),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__1063 (
            .O(N__4938),
            .I(N__4932));
    InMux I__1062 (
            .O(N__4937),
            .I(N__4927));
    InMux I__1061 (
            .O(N__4936),
            .I(N__4927));
    InMux I__1060 (
            .O(N__4935),
            .I(N__4924));
    InMux I__1059 (
            .O(N__4932),
            .I(N__4921));
    LocalMux I__1058 (
            .O(N__4927),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1057 (
            .O(N__4924),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1056 (
            .O(N__4921),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__1055 (
            .O(N__4914),
            .I(N__4911));
    LocalMux I__1054 (
            .O(N__4911),
            .I(N__4907));
    InMux I__1053 (
            .O(N__4910),
            .I(N__4904));
    Odrv4 I__1052 (
            .O(N__4907),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1051 (
            .O(N__4904),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__1050 (
            .O(N__4899),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__1049 (
            .O(N__4896),
            .I(N__4892));
    InMux I__1048 (
            .O(N__4895),
            .I(N__4889));
    LocalMux I__1047 (
            .O(N__4892),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1046 (
            .O(N__4889),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__1045 (
            .O(N__4884),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__1044 (
            .O(N__4881),
            .I(N__4877));
    InMux I__1043 (
            .O(N__4880),
            .I(N__4874));
    LocalMux I__1042 (
            .O(N__4877),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1041 (
            .O(N__4874),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__1040 (
            .O(N__4869),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__1039 (
            .O(N__4866),
            .I(N__4862));
    InMux I__1038 (
            .O(N__4865),
            .I(N__4859));
    LocalMux I__1037 (
            .O(N__4862),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1036 (
            .O(N__4859),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__1035 (
            .O(N__4854),
            .I(N__4851));
    LocalMux I__1034 (
            .O(N__4851),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1033 (
            .O(N__4848),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__1032 (
            .O(N__4845),
            .I(N__4841));
    InMux I__1031 (
            .O(N__4844),
            .I(N__4838));
    InMux I__1030 (
            .O(N__4841),
            .I(N__4835));
    LocalMux I__1029 (
            .O(N__4838),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__1028 (
            .O(N__4835),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__1027 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__1026 (
            .O(N__4827),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1025 (
            .O(N__4824),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    CascadeMux I__1024 (
            .O(N__4821),
            .I(N__4818));
    InMux I__1023 (
            .O(N__4818),
            .I(N__4814));
    InMux I__1022 (
            .O(N__4817),
            .I(N__4811));
    LocalMux I__1021 (
            .O(N__4814),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1020 (
            .O(N__4811),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__1019 (
            .O(N__4806),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__1018 (
            .O(N__4803),
            .I(N__4799));
    InMux I__1017 (
            .O(N__4802),
            .I(N__4796));
    LocalMux I__1016 (
            .O(N__4799),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1015 (
            .O(N__4796),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1014 (
            .O(N__4791),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    CascadeMux I__1013 (
            .O(N__4788),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    InMux I__1012 (
            .O(N__4785),
            .I(N__4781));
    InMux I__1011 (
            .O(N__4784),
            .I(N__4778));
    LocalMux I__1010 (
            .O(N__4781),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    LocalMux I__1009 (
            .O(N__4778),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__1008 (
            .O(N__4773),
            .I(N__4764));
    InMux I__1007 (
            .O(N__4772),
            .I(N__4764));
    InMux I__1006 (
            .O(N__4771),
            .I(N__4761));
    InMux I__1005 (
            .O(N__4770),
            .I(N__4758));
    InMux I__1004 (
            .O(N__4769),
            .I(N__4755));
    LocalMux I__1003 (
            .O(N__4764),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1002 (
            .O(N__4761),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1001 (
            .O(N__4758),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1000 (
            .O(N__4755),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__999 (
            .O(N__4746),
            .I(N__4740));
    InMux I__998 (
            .O(N__4745),
            .I(N__4737));
    InMux I__997 (
            .O(N__4744),
            .I(N__4732));
    InMux I__996 (
            .O(N__4743),
            .I(N__4732));
    LocalMux I__995 (
            .O(N__4740),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__994 (
            .O(N__4737),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__993 (
            .O(N__4732),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__992 (
            .O(N__4725),
            .I(N__4721));
    CascadeMux I__991 (
            .O(N__4724),
            .I(N__4716));
    LocalMux I__990 (
            .O(N__4721),
            .I(N__4713));
    InMux I__989 (
            .O(N__4720),
            .I(N__4710));
    InMux I__988 (
            .O(N__4719),
            .I(N__4705));
    InMux I__987 (
            .O(N__4716),
            .I(N__4705));
    Odrv4 I__986 (
            .O(N__4713),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__985 (
            .O(N__4710),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__984 (
            .O(N__4705),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__983 (
            .O(N__4698),
            .I(N__4693));
    InMux I__982 (
            .O(N__4697),
            .I(N__4688));
    InMux I__981 (
            .O(N__4696),
            .I(N__4688));
    LocalMux I__980 (
            .O(N__4693),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__979 (
            .O(N__4688),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__978 (
            .O(N__4683),
            .I(N__4677));
    InMux I__977 (
            .O(N__4682),
            .I(N__4674));
    InMux I__976 (
            .O(N__4681),
            .I(N__4671));
    InMux I__975 (
            .O(N__4680),
            .I(N__4668));
    LocalMux I__974 (
            .O(N__4677),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__973 (
            .O(N__4674),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__972 (
            .O(N__4671),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__971 (
            .O(N__4668),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__970 (
            .O(N__4659),
            .I(N__4650));
    InMux I__969 (
            .O(N__4658),
            .I(N__4645));
    InMux I__968 (
            .O(N__4657),
            .I(N__4645));
    InMux I__967 (
            .O(N__4656),
            .I(N__4642));
    InMux I__966 (
            .O(N__4655),
            .I(N__4633));
    InMux I__965 (
            .O(N__4654),
            .I(N__4633));
    InMux I__964 (
            .O(N__4653),
            .I(N__4633));
    InMux I__963 (
            .O(N__4650),
            .I(N__4633));
    LocalMux I__962 (
            .O(N__4645),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__961 (
            .O(N__4642),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__960 (
            .O(N__4633),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__959 (
            .O(N__4626),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__958 (
            .O(N__4623),
            .I(N__4616));
    InMux I__957 (
            .O(N__4622),
            .I(N__4616));
    InMux I__956 (
            .O(N__4621),
            .I(N__4613));
    LocalMux I__955 (
            .O(N__4616),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__954 (
            .O(N__4613),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__953 (
            .O(N__4608),
            .I(N__4601));
    InMux I__952 (
            .O(N__4607),
            .I(N__4598));
    InMux I__951 (
            .O(N__4606),
            .I(N__4591));
    InMux I__950 (
            .O(N__4605),
            .I(N__4591));
    InMux I__949 (
            .O(N__4604),
            .I(N__4591));
    LocalMux I__948 (
            .O(N__4601),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__947 (
            .O(N__4598),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__946 (
            .O(N__4591),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__945 (
            .O(N__4584),
            .I(N__4579));
    InMux I__944 (
            .O(N__4583),
            .I(N__4575));
    InMux I__943 (
            .O(N__4582),
            .I(N__4572));
    InMux I__942 (
            .O(N__4579),
            .I(N__4567));
    InMux I__941 (
            .O(N__4578),
            .I(N__4567));
    LocalMux I__940 (
            .O(N__4575),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__939 (
            .O(N__4572),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__938 (
            .O(N__4567),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__937 (
            .O(N__4560),
            .I(N__4554));
    InMux I__936 (
            .O(N__4559),
            .I(N__4554));
    LocalMux I__935 (
            .O(N__4554),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__934 (
            .O(N__4551),
            .I(N__4547));
    InMux I__933 (
            .O(N__4550),
            .I(N__4544));
    LocalMux I__932 (
            .O(N__4547),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__931 (
            .O(N__4544),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__930 (
            .O(N__4539),
            .I(N__4536));
    LocalMux I__929 (
            .O(N__4536),
            .I(N__4533));
    Odrv4 I__928 (
            .O(N__4533),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    CascadeMux I__927 (
            .O(N__4530),
            .I(N__4527));
    InMux I__926 (
            .O(N__4527),
            .I(N__4520));
    InMux I__925 (
            .O(N__4526),
            .I(N__4517));
    InMux I__924 (
            .O(N__4525),
            .I(N__4513));
    InMux I__923 (
            .O(N__4524),
            .I(N__4510));
    InMux I__922 (
            .O(N__4523),
            .I(N__4507));
    LocalMux I__921 (
            .O(N__4520),
            .I(N__4502));
    LocalMux I__920 (
            .O(N__4517),
            .I(N__4502));
    InMux I__919 (
            .O(N__4516),
            .I(N__4499));
    LocalMux I__918 (
            .O(N__4513),
            .I(N__4496));
    LocalMux I__917 (
            .O(N__4510),
            .I(N__4493));
    LocalMux I__916 (
            .O(N__4507),
            .I(N__4490));
    Span4Mux_v I__915 (
            .O(N__4502),
            .I(N__4485));
    LocalMux I__914 (
            .O(N__4499),
            .I(N__4485));
    Span4Mux_v I__913 (
            .O(N__4496),
            .I(N__4482));
    Span4Mux_v I__912 (
            .O(N__4493),
            .I(N__4479));
    Span4Mux_v I__911 (
            .O(N__4490),
            .I(N__4476));
    Span4Mux_h I__910 (
            .O(N__4485),
            .I(N__4472));
    Sp12to4 I__909 (
            .O(N__4482),
            .I(N__4465));
    Sp12to4 I__908 (
            .O(N__4479),
            .I(N__4465));
    Sp12to4 I__907 (
            .O(N__4476),
            .I(N__4465));
    InMux I__906 (
            .O(N__4475),
            .I(N__4462));
    Span4Mux_v I__905 (
            .O(N__4472),
            .I(N__4459));
    Span12Mux_h I__904 (
            .O(N__4465),
            .I(N__4454));
    LocalMux I__903 (
            .O(N__4462),
            .I(N__4454));
    Odrv4 I__902 (
            .O(N__4459),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv12 I__901 (
            .O(N__4454),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    InMux I__900 (
            .O(N__4449),
            .I(N__4444));
    InMux I__899 (
            .O(N__4448),
            .I(N__4441));
    InMux I__898 (
            .O(N__4447),
            .I(N__4438));
    LocalMux I__897 (
            .O(N__4444),
            .I(N__4435));
    LocalMux I__896 (
            .O(N__4441),
            .I(N__4430));
    LocalMux I__895 (
            .O(N__4438),
            .I(N__4430));
    Span4Mux_v I__894 (
            .O(N__4435),
            .I(N__4427));
    Span4Mux_v I__893 (
            .O(N__4430),
            .I(N__4424));
    Sp12to4 I__892 (
            .O(N__4427),
            .I(N__4419));
    Sp12to4 I__891 (
            .O(N__4424),
            .I(N__4419));
    Span12Mux_h I__890 (
            .O(N__4419),
            .I(N__4416));
    Span12Mux_v I__889 (
            .O(N__4416),
            .I(N__4413));
    Odrv12 I__888 (
            .O(N__4413),
            .I(OVL_c));
    InMux I__887 (
            .O(N__4410),
            .I(N__4406));
    InMux I__886 (
            .O(N__4409),
            .I(N__4403));
    LocalMux I__885 (
            .O(N__4406),
            .I(N__4399));
    LocalMux I__884 (
            .O(N__4403),
            .I(N__4396));
    InMux I__883 (
            .O(N__4402),
            .I(N__4393));
    Span12Mux_h I__882 (
            .O(N__4399),
            .I(N__4386));
    Sp12to4 I__881 (
            .O(N__4396),
            .I(N__4386));
    LocalMux I__880 (
            .O(N__4393),
            .I(N__4386));
    Odrv12 I__879 (
            .O(N__4386),
            .I(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ));
    IoInMux I__878 (
            .O(N__4383),
            .I(N__4380));
    LocalMux I__877 (
            .O(N__4380),
            .I(N__4377));
    Span4Mux_s3_v I__876 (
            .O(N__4377),
            .I(N__4374));
    Span4Mux_v I__875 (
            .O(N__4374),
            .I(N__4371));
    Span4Mux_v I__874 (
            .O(N__4371),
            .I(N__4368));
    Span4Mux_v I__873 (
            .O(N__4368),
            .I(N__4365));
    Odrv4 I__872 (
            .O(N__4365),
            .I(U409_ADDRESS_DECODE_un1_nRAMSPACE_i));
    IoInMux I__871 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__870 (
            .O(N__4359),
            .I(N__4356));
    Span4Mux_s3_v I__869 (
            .O(N__4356),
            .I(N__4353));
    Span4Mux_h I__868 (
            .O(N__4353),
            .I(N__4350));
    Odrv4 I__867 (
            .O(N__4350),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__866 (
            .O(N__4347),
            .I(\U409_CIA.N_20_cascade_ ));
    InMux I__865 (
            .O(N__4344),
            .I(N__4340));
    InMux I__864 (
            .O(N__4343),
            .I(N__4337));
    LocalMux I__863 (
            .O(N__4340),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    LocalMux I__862 (
            .O(N__4337),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    InMux I__861 (
            .O(N__4332),
            .I(N__4329));
    LocalMux I__860 (
            .O(N__4329),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__859 (
            .O(N__4326),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    IoInMux I__858 (
            .O(N__4323),
            .I(N__4320));
    LocalMux I__857 (
            .O(N__4320),
            .I(N__4317));
    Span4Mux_s1_v I__856 (
            .O(N__4317),
            .I(N__4314));
    Span4Mux_v I__855 (
            .O(N__4314),
            .I(N__4311));
    Sp12to4 I__854 (
            .O(N__4311),
            .I(N__4308));
    Span12Mux_h I__853 (
            .O(N__4308),
            .I(N__4304));
    InMux I__852 (
            .O(N__4307),
            .I(N__4301));
    Span12Mux_v I__851 (
            .O(N__4304),
            .I(N__4295));
    LocalMux I__850 (
            .O(N__4301),
            .I(N__4295));
    InMux I__849 (
            .O(N__4300),
            .I(N__4292));
    Odrv12 I__848 (
            .O(N__4295),
            .I(CLKCIA_c));
    LocalMux I__847 (
            .O(N__4292),
            .I(CLKCIA_c));
    InMux I__846 (
            .O(N__4287),
            .I(N__4284));
    LocalMux I__845 (
            .O(N__4284),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ));
    CascadeMux I__844 (
            .O(N__4281),
            .I(N__4278));
    InMux I__843 (
            .O(N__4278),
            .I(N__4271));
    InMux I__842 (
            .O(N__4277),
            .I(N__4271));
    InMux I__841 (
            .O(N__4276),
            .I(N__4268));
    LocalMux I__840 (
            .O(N__4271),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    LocalMux I__839 (
            .O(N__4268),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__838 (
            .O(N__4263),
            .I(N__4259));
    InMux I__837 (
            .O(N__4262),
            .I(N__4253));
    InMux I__836 (
            .O(N__4259),
            .I(N__4246));
    InMux I__835 (
            .O(N__4258),
            .I(N__4246));
    InMux I__834 (
            .O(N__4257),
            .I(N__4246));
    InMux I__833 (
            .O(N__4256),
            .I(N__4243));
    LocalMux I__832 (
            .O(N__4253),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__831 (
            .O(N__4246),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__830 (
            .O(N__4243),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__829 (
            .O(N__4236),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    IoInMux I__828 (
            .O(N__4233),
            .I(N__4230));
    LocalMux I__827 (
            .O(N__4230),
            .I(N__4227));
    Span4Mux_s3_v I__826 (
            .O(N__4227),
            .I(N__4224));
    Span4Mux_h I__825 (
            .O(N__4224),
            .I(N__4221));
    Sp12to4 I__824 (
            .O(N__4221),
            .I(N__4218));
    Span12Mux_v I__823 (
            .O(N__4218),
            .I(N__4214));
    InMux I__822 (
            .O(N__4217),
            .I(N__4211));
    Odrv12 I__821 (
            .O(N__4214),
            .I(TICK50_c));
    LocalMux I__820 (
            .O(N__4211),
            .I(TICK50_c));
    CascadeMux I__819 (
            .O(N__4206),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    CascadeMux I__818 (
            .O(N__4203),
            .I(\U409_CIA.N_9_cascade_ ));
    InMux I__817 (
            .O(N__4200),
            .I(N__4195));
    InMux I__816 (
            .O(N__4199),
            .I(N__4190));
    InMux I__815 (
            .O(N__4198),
            .I(N__4190));
    LocalMux I__814 (
            .O(N__4195),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__813 (
            .O(N__4190),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    InMux I__812 (
            .O(N__4185),
            .I(N__4178));
    InMux I__811 (
            .O(N__4184),
            .I(N__4178));
    InMux I__810 (
            .O(N__4183),
            .I(N__4175));
    LocalMux I__809 (
            .O(N__4178),
            .I(N__4170));
    LocalMux I__808 (
            .O(N__4175),
            .I(N__4170));
    Odrv12 I__807 (
            .O(N__4170),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__806 (
            .O(N__4167),
            .I(N__4163));
    InMux I__805 (
            .O(N__4166),
            .I(N__4158));
    InMux I__804 (
            .O(N__4163),
            .I(N__4151));
    InMux I__803 (
            .O(N__4162),
            .I(N__4151));
    InMux I__802 (
            .O(N__4161),
            .I(N__4151));
    LocalMux I__801 (
            .O(N__4158),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__800 (
            .O(N__4151),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__799 (
            .O(N__4146),
            .I(N__4142));
    InMux I__798 (
            .O(N__4145),
            .I(N__4136));
    InMux I__797 (
            .O(N__4142),
            .I(N__4136));
    CascadeMux I__796 (
            .O(N__4141),
            .I(N__4133));
    LocalMux I__795 (
            .O(N__4136),
            .I(N__4130));
    InMux I__794 (
            .O(N__4133),
            .I(N__4127));
    Span4Mux_v I__793 (
            .O(N__4130),
            .I(N__4124));
    LocalMux I__792 (
            .O(N__4127),
            .I(N__4121));
    Span4Mux_h I__791 (
            .O(N__4124),
            .I(N__4118));
    Span4Mux_v I__790 (
            .O(N__4121),
            .I(N__4115));
    Sp12to4 I__789 (
            .O(N__4118),
            .I(N__4110));
    Sp12to4 I__788 (
            .O(N__4115),
            .I(N__4110));
    Span12Mux_h I__787 (
            .O(N__4110),
            .I(N__4107));
    Odrv12 I__786 (
            .O(N__4107),
            .I(\U409_CIA.g0Z0Z_13 ));
    InMux I__785 (
            .O(N__4104),
            .I(N__4098));
    InMux I__784 (
            .O(N__4103),
            .I(N__4098));
    LocalMux I__783 (
            .O(N__4098),
            .I(N__4095));
    Odrv12 I__782 (
            .O(N__4095),
            .I(CIA_ENABLEm));
    CascadeMux I__781 (
            .O(N__4092),
            .I(N__4088));
    InMux I__780 (
            .O(N__4091),
            .I(N__4083));
    InMux I__779 (
            .O(N__4088),
            .I(N__4080));
    InMux I__778 (
            .O(N__4087),
            .I(N__4077));
    CascadeMux I__777 (
            .O(N__4086),
            .I(N__4074));
    LocalMux I__776 (
            .O(N__4083),
            .I(N__4071));
    LocalMux I__775 (
            .O(N__4080),
            .I(N__4066));
    LocalMux I__774 (
            .O(N__4077),
            .I(N__4066));
    InMux I__773 (
            .O(N__4074),
            .I(N__4063));
    Odrv4 I__772 (
            .O(N__4071),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    Odrv4 I__771 (
            .O(N__4066),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__770 (
            .O(N__4063),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    CascadeMux I__769 (
            .O(N__4056),
            .I(N__4052));
    InMux I__768 (
            .O(N__4055),
            .I(N__4048));
    InMux I__767 (
            .O(N__4052),
            .I(N__4045));
    InMux I__766 (
            .O(N__4051),
            .I(N__4042));
    LocalMux I__765 (
            .O(N__4048),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__764 (
            .O(N__4045),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__763 (
            .O(N__4042),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__762 (
            .O(N__4035),
            .I(N__4031));
    InMux I__761 (
            .O(N__4034),
            .I(N__4028));
    LocalMux I__760 (
            .O(N__4031),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__759 (
            .O(N__4028),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    CascadeMux I__758 (
            .O(N__4023),
            .I(N__4020));
    InMux I__757 (
            .O(N__4020),
            .I(N__4016));
    InMux I__756 (
            .O(N__4019),
            .I(N__4013));
    LocalMux I__755 (
            .O(N__4016),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__754 (
            .O(N__4013),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__753 (
            .O(N__4008),
            .I(N__4004));
    InMux I__752 (
            .O(N__4007),
            .I(N__4001));
    LocalMux I__751 (
            .O(N__4004),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__750 (
            .O(N__4001),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__749 (
            .O(N__3996),
            .I(N__3991));
    CascadeMux I__748 (
            .O(N__3995),
            .I(N__3988));
    CascadeMux I__747 (
            .O(N__3994),
            .I(N__3982));
    InMux I__746 (
            .O(N__3991),
            .I(N__3976));
    InMux I__745 (
            .O(N__3988),
            .I(N__3976));
    InMux I__744 (
            .O(N__3987),
            .I(N__3973));
    InMux I__743 (
            .O(N__3986),
            .I(N__3964));
    InMux I__742 (
            .O(N__3985),
            .I(N__3964));
    InMux I__741 (
            .O(N__3982),
            .I(N__3964));
    InMux I__740 (
            .O(N__3981),
            .I(N__3964));
    LocalMux I__739 (
            .O(N__3976),
            .I(N__3961));
    LocalMux I__738 (
            .O(N__3973),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__737 (
            .O(N__3964),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__736 (
            .O(N__3961),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__735 (
            .O(N__3954),
            .I(N__3945));
    InMux I__734 (
            .O(N__3953),
            .I(N__3940));
    InMux I__733 (
            .O(N__3952),
            .I(N__3940));
    InMux I__732 (
            .O(N__3951),
            .I(N__3937));
    InMux I__731 (
            .O(N__3950),
            .I(N__3930));
    InMux I__730 (
            .O(N__3949),
            .I(N__3930));
    InMux I__729 (
            .O(N__3948),
            .I(N__3930));
    LocalMux I__728 (
            .O(N__3945),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__727 (
            .O(N__3940),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__726 (
            .O(N__3937),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__725 (
            .O(N__3930),
            .I(\U409_TICK.TICK603_9 ));
    InMux I__724 (
            .O(N__3921),
            .I(N__3914));
    InMux I__723 (
            .O(N__3920),
            .I(N__3911));
    InMux I__722 (
            .O(N__3919),
            .I(N__3906));
    InMux I__721 (
            .O(N__3918),
            .I(N__3901));
    InMux I__720 (
            .O(N__3917),
            .I(N__3901));
    LocalMux I__719 (
            .O(N__3914),
            .I(N__3896));
    LocalMux I__718 (
            .O(N__3911),
            .I(N__3896));
    InMux I__717 (
            .O(N__3910),
            .I(N__3891));
    InMux I__716 (
            .O(N__3909),
            .I(N__3891));
    LocalMux I__715 (
            .O(N__3906),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__714 (
            .O(N__3901),
            .I(\U409_TICK.TICK603_14 ));
    Odrv4 I__713 (
            .O(N__3896),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__712 (
            .O(N__3891),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__711 (
            .O(N__3882),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__710 (
            .O(N__3879),
            .I(N__3876));
    LocalMux I__709 (
            .O(N__3876),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__708 (
            .O(N__3873),
            .I(N__3869));
    InMux I__707 (
            .O(N__3872),
            .I(N__3866));
    LocalMux I__706 (
            .O(N__3869),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__705 (
            .O(N__3866),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__704 (
            .O(N__3861),
            .I(N__3858));
    LocalMux I__703 (
            .O(N__3858),
            .I(N__3855));
    Odrv4 I__702 (
            .O(N__3855),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__701 (
            .O(N__3852),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    CascadeMux I__700 (
            .O(N__3849),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    IoInMux I__699 (
            .O(N__3846),
            .I(N__3843));
    LocalMux I__698 (
            .O(N__3843),
            .I(N__3840));
    IoSpan4Mux I__697 (
            .O(N__3840),
            .I(N__3837));
    Span4Mux_s3_v I__696 (
            .O(N__3837),
            .I(N__3834));
    Span4Mux_v I__695 (
            .O(N__3834),
            .I(N__3831));
    Sp12to4 I__694 (
            .O(N__3831),
            .I(N__3828));
    Span12Mux_v I__693 (
            .O(N__3828),
            .I(N__3824));
    InMux I__692 (
            .O(N__3827),
            .I(N__3821));
    Odrv12 I__691 (
            .O(N__3824),
            .I(TACK_OUTn));
    LocalMux I__690 (
            .O(N__3821),
            .I(TACK_OUTn));
    InMux I__689 (
            .O(N__3816),
            .I(N__3807));
    InMux I__688 (
            .O(N__3815),
            .I(N__3807));
    InMux I__687 (
            .O(N__3814),
            .I(N__3807));
    LocalMux I__686 (
            .O(N__3807),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__685 (
            .O(N__3804),
            .I(N__3795));
    InMux I__684 (
            .O(N__3803),
            .I(N__3795));
    InMux I__683 (
            .O(N__3802),
            .I(N__3795));
    LocalMux I__682 (
            .O(N__3795),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    CascadeMux I__681 (
            .O(N__3792),
            .I(N__3789));
    InMux I__680 (
            .O(N__3789),
            .I(N__3786));
    LocalMux I__679 (
            .O(N__3786),
            .I(N__3783));
    Odrv4 I__678 (
            .O(N__3783),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    InMux I__677 (
            .O(N__3780),
            .I(N__3777));
    LocalMux I__676 (
            .O(N__3777),
            .I(N__3774));
    Span4Mux_v I__675 (
            .O(N__3774),
            .I(N__3771));
    Sp12to4 I__674 (
            .O(N__3771),
            .I(N__3768));
    Span12Mux_h I__673 (
            .O(N__3768),
            .I(N__3765));
    Odrv12 I__672 (
            .O(N__3765),
            .I(A_c_13));
    IoInMux I__671 (
            .O(N__3762),
            .I(N__3759));
    LocalMux I__670 (
            .O(N__3759),
            .I(N__3756));
    Span4Mux_s2_h I__669 (
            .O(N__3756),
            .I(N__3753));
    Span4Mux_v I__668 (
            .O(N__3753),
            .I(N__3750));
    Span4Mux_h I__667 (
            .O(N__3750),
            .I(N__3747));
    Sp12to4 I__666 (
            .O(N__3747),
            .I(N__3744));
    Span12Mux_h I__665 (
            .O(N__3744),
            .I(N__3741));
    Odrv12 I__664 (
            .O(N__3741),
            .I(U409_ADDRESS_DECODE_un1_nCIACS1_i));
    InMux I__663 (
            .O(N__3738),
            .I(N__3735));
    LocalMux I__662 (
            .O(N__3735),
            .I(N__3732));
    Span4Mux_v I__661 (
            .O(N__3732),
            .I(N__3729));
    Sp12to4 I__660 (
            .O(N__3729),
            .I(N__3726));
    Span12Mux_h I__659 (
            .O(N__3726),
            .I(N__3723));
    Odrv12 I__658 (
            .O(N__3723),
            .I(A_c_12));
    IoInMux I__657 (
            .O(N__3720),
            .I(N__3717));
    LocalMux I__656 (
            .O(N__3717),
            .I(N__3714));
    Span4Mux_s0_h I__655 (
            .O(N__3714),
            .I(N__3711));
    Sp12to4 I__654 (
            .O(N__3711),
            .I(N__3708));
    Span12Mux_s9_v I__653 (
            .O(N__3708),
            .I(N__3705));
    Span12Mux_h I__652 (
            .O(N__3705),
            .I(N__3702));
    Odrv12 I__651 (
            .O(N__3702),
            .I(U409_ADDRESS_DECODE_un1_nCIACS0_i));
    CascadeMux I__650 (
            .O(N__3699),
            .I(N__3696));
    InMux I__649 (
            .O(N__3696),
            .I(N__3692));
    InMux I__648 (
            .O(N__3695),
            .I(N__3688));
    LocalMux I__647 (
            .O(N__3692),
            .I(N__3685));
    InMux I__646 (
            .O(N__3691),
            .I(N__3682));
    LocalMux I__645 (
            .O(N__3688),
            .I(N__3679));
    Span4Mux_h I__644 (
            .O(N__3685),
            .I(N__3674));
    LocalMux I__643 (
            .O(N__3682),
            .I(N__3674));
    Span4Mux_v I__642 (
            .O(N__3679),
            .I(N__3671));
    Span4Mux_v I__641 (
            .O(N__3674),
            .I(N__3668));
    Sp12to4 I__640 (
            .O(N__3671),
            .I(N__3663));
    Sp12to4 I__639 (
            .O(N__3668),
            .I(N__3663));
    Span12Mux_h I__638 (
            .O(N__3663),
            .I(N__3660));
    Span12Mux_v I__637 (
            .O(N__3660),
            .I(N__3657));
    Odrv12 I__636 (
            .O(N__3657),
            .I(TSn_c));
    IoInMux I__635 (
            .O(N__3654),
            .I(N__3648));
    InMux I__634 (
            .O(N__3653),
            .I(N__3645));
    CascadeMux I__633 (
            .O(N__3652),
            .I(N__3642));
    CascadeMux I__632 (
            .O(N__3651),
            .I(N__3637));
    LocalMux I__631 (
            .O(N__3648),
            .I(N__3634));
    LocalMux I__630 (
            .O(N__3645),
            .I(N__3631));
    InMux I__629 (
            .O(N__3642),
            .I(N__3628));
    InMux I__628 (
            .O(N__3641),
            .I(N__3623));
    InMux I__627 (
            .O(N__3640),
            .I(N__3623));
    InMux I__626 (
            .O(N__3637),
            .I(N__3620));
    IoSpan4Mux I__625 (
            .O(N__3634),
            .I(N__3617));
    Span4Mux_h I__624 (
            .O(N__3631),
            .I(N__3612));
    LocalMux I__623 (
            .O(N__3628),
            .I(N__3612));
    LocalMux I__622 (
            .O(N__3623),
            .I(N__3607));
    LocalMux I__621 (
            .O(N__3620),
            .I(N__3607));
    Span4Mux_s0_v I__620 (
            .O(N__3617),
            .I(N__3604));
    Span4Mux_v I__619 (
            .O(N__3612),
            .I(N__3601));
    Span4Mux_v I__618 (
            .O(N__3607),
            .I(N__3598));
    Sp12to4 I__617 (
            .O(N__3604),
            .I(N__3595));
    Span4Mux_v I__616 (
            .O(N__3601),
            .I(N__3592));
    Sp12to4 I__615 (
            .O(N__3598),
            .I(N__3589));
    Span12Mux_v I__614 (
            .O(N__3595),
            .I(N__3586));
    Sp12to4 I__613 (
            .O(N__3592),
            .I(N__3583));
    Span12Mux_h I__612 (
            .O(N__3589),
            .I(N__3580));
    Span12Mux_v I__611 (
            .O(N__3586),
            .I(N__3577));
    Span12Mux_h I__610 (
            .O(N__3583),
            .I(N__3574));
    Span12Mux_v I__609 (
            .O(N__3580),
            .I(N__3571));
    Odrv12 I__608 (
            .O(N__3577),
            .I(CLK40_IN_c));
    Odrv12 I__607 (
            .O(N__3574),
            .I(CLK40_IN_c));
    Odrv12 I__606 (
            .O(N__3571),
            .I(CLK40_IN_c));
    InMux I__605 (
            .O(N__3564),
            .I(N__3561));
    LocalMux I__604 (
            .O(N__3561),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__603 (
            .O(N__3558),
            .I(N__3554));
    InMux I__602 (
            .O(N__3557),
            .I(N__3551));
    LocalMux I__601 (
            .O(N__3554),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__600 (
            .O(N__3551),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__599 (
            .O(N__3546),
            .I(N__3542));
    InMux I__598 (
            .O(N__3545),
            .I(N__3539));
    LocalMux I__597 (
            .O(N__3542),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__596 (
            .O(N__3539),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__595 (
            .O(N__3534),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ));
    InMux I__594 (
            .O(N__3531),
            .I(N__3527));
    InMux I__593 (
            .O(N__3530),
            .I(N__3524));
    LocalMux I__592 (
            .O(N__3527),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__591 (
            .O(N__3524),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__590 (
            .O(N__3519),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__589 (
            .O(N__3516),
            .I(N__3512));
    InMux I__588 (
            .O(N__3515),
            .I(N__3509));
    LocalMux I__587 (
            .O(N__3512),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__586 (
            .O(N__3509),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__585 (
            .O(N__3504),
            .I(N__3501));
    LocalMux I__584 (
            .O(N__3501),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__583 (
            .O(N__3498),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__582 (
            .O(N__3495),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__581 (
            .O(N__3492),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__580 (
            .O(N__3489),
            .I(N__3485));
    InMux I__579 (
            .O(N__3488),
            .I(N__3482));
    LocalMux I__578 (
            .O(N__3485),
            .I(N__3479));
    LocalMux I__577 (
            .O(N__3482),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    Odrv4 I__576 (
            .O(N__3479),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__575 (
            .O(N__3474),
            .I(N__3468));
    InMux I__574 (
            .O(N__3473),
            .I(N__3461));
    InMux I__573 (
            .O(N__3472),
            .I(N__3461));
    InMux I__572 (
            .O(N__3471),
            .I(N__3461));
    LocalMux I__571 (
            .O(N__3468),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__570 (
            .O(N__3461),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    SRMux I__569 (
            .O(N__3456),
            .I(N__3453));
    LocalMux I__568 (
            .O(N__3453),
            .I(N__3450));
    Span4Mux_h I__567 (
            .O(N__3450),
            .I(N__3447));
    Odrv4 I__566 (
            .O(N__3447),
            .I(\U409_TRANSFER_ACK.RESETn_c_i ));
    CascadeMux I__565 (
            .O(N__3444),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ));
    CascadeMux I__564 (
            .O(N__3441),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__563 (
            .O(N__3438),
            .I(N__3434));
    InMux I__562 (
            .O(N__3437),
            .I(N__3431));
    LocalMux I__561 (
            .O(N__3434),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__560 (
            .O(N__3431),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__559 (
            .O(N__3426),
            .I(N__3423));
    LocalMux I__558 (
            .O(N__3423),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__557 (
            .O(N__3420),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__556 (
            .O(N__3417),
            .I(N__3413));
    InMux I__555 (
            .O(N__3416),
            .I(N__3410));
    LocalMux I__554 (
            .O(N__3413),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__553 (
            .O(N__3410),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__552 (
            .O(N__3405),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__551 (
            .O(N__3402),
            .I(N__3398));
    CascadeMux I__550 (
            .O(N__3401),
            .I(N__3395));
    InMux I__549 (
            .O(N__3398),
            .I(N__3392));
    InMux I__548 (
            .O(N__3395),
            .I(N__3389));
    LocalMux I__547 (
            .O(N__3392),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__546 (
            .O(N__3389),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__545 (
            .O(N__3384),
            .I(N__3381));
    LocalMux I__544 (
            .O(N__3381),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__543 (
            .O(N__3378),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__542 (
            .O(N__3375),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__541 (
            .O(N__3372),
            .I(N__3368));
    InMux I__540 (
            .O(N__3371),
            .I(N__3365));
    LocalMux I__539 (
            .O(N__3368),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__538 (
            .O(N__3365),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__537 (
            .O(N__3360),
            .I(N__3357));
    InMux I__536 (
            .O(N__3357),
            .I(N__3354));
    LocalMux I__535 (
            .O(N__3354),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__534 (
            .O(N__3351),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__533 (
            .O(N__3348),
            .I(N__3344));
    InMux I__532 (
            .O(N__3347),
            .I(N__3341));
    LocalMux I__531 (
            .O(N__3344),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__530 (
            .O(N__3341),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__529 (
            .O(N__3336),
            .I(N__3333));
    LocalMux I__528 (
            .O(N__3333),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__527 (
            .O(N__3330),
            .I(bfn_10_7_0_));
    InMux I__526 (
            .O(N__3327),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__525 (
            .O(N__3324),
            .I(N__3321));
    LocalMux I__524 (
            .O(N__3321),
            .I(N__3317));
    InMux I__523 (
            .O(N__3320),
            .I(N__3314));
    Odrv4 I__522 (
            .O(N__3317),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__521 (
            .O(N__3314),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__520 (
            .O(N__3309),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__519 (
            .O(N__3306),
            .I(N__3302));
    InMux I__518 (
            .O(N__3305),
            .I(N__3299));
    LocalMux I__517 (
            .O(N__3302),
            .I(N__3296));
    LocalMux I__516 (
            .O(N__3299),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    Odrv4 I__515 (
            .O(N__3296),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__514 (
            .O(N__3291),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    CascadeMux I__513 (
            .O(N__3288),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    CascadeMux I__512 (
            .O(N__3285),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    IoInMux I__511 (
            .O(N__3282),
            .I(N__3279));
    LocalMux I__510 (
            .O(N__3279),
            .I(N__3276));
    Span4Mux_s2_v I__509 (
            .O(N__3276),
            .I(N__3273));
    Span4Mux_v I__508 (
            .O(N__3273),
            .I(N__3270));
    Span4Mux_v I__507 (
            .O(N__3270),
            .I(N__3267));
    Span4Mux_h I__506 (
            .O(N__3267),
            .I(N__3263));
    InMux I__505 (
            .O(N__3266),
            .I(N__3260));
    Odrv4 I__504 (
            .O(N__3263),
            .I(TICK60_c));
    LocalMux I__503 (
            .O(N__3260),
            .I(TICK60_c));
    InMux I__502 (
            .O(N__3255),
            .I(N__3252));
    LocalMux I__501 (
            .O(N__3252),
            .I(\U409_TICK.TICK603_8 ));
    InMux I__500 (
            .O(N__3249),
            .I(N__3245));
    InMux I__499 (
            .O(N__3248),
            .I(N__3242));
    LocalMux I__498 (
            .O(N__3245),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__497 (
            .O(N__3242),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__496 (
            .O(N__3237),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__495 (
            .O(N__3234),
            .I(N__3230));
    InMux I__494 (
            .O(N__3233),
            .I(N__3227));
    LocalMux I__493 (
            .O(N__3230),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__492 (
            .O(N__3227),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__491 (
            .O(N__3222),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    CascadeMux I__490 (
            .O(N__3219),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ));
    InMux I__489 (
            .O(N__3216),
            .I(N__3213));
    LocalMux I__488 (
            .O(N__3213),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ));
    InMux I__487 (
            .O(N__3210),
            .I(N__3207));
    LocalMux I__486 (
            .O(N__3207),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ));
    CascadeMux I__485 (
            .O(N__3204),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ));
    InMux I__484 (
            .O(N__3201),
            .I(N__3189));
    InMux I__483 (
            .O(N__3200),
            .I(N__3189));
    InMux I__482 (
            .O(N__3199),
            .I(N__3189));
    InMux I__481 (
            .O(N__3198),
            .I(N__3189));
    LocalMux I__480 (
            .O(N__3189),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__479 (
            .O(N__3186),
            .I(N__3180));
    InMux I__478 (
            .O(N__3185),
            .I(N__3174));
    InMux I__477 (
            .O(N__3184),
            .I(N__3174));
    InMux I__476 (
            .O(N__3183),
            .I(N__3167));
    InMux I__475 (
            .O(N__3180),
            .I(N__3167));
    InMux I__474 (
            .O(N__3179),
            .I(N__3167));
    LocalMux I__473 (
            .O(N__3174),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__472 (
            .O(N__3167),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__471 (
            .O(N__3162),
            .I(N__3159));
    LocalMux I__470 (
            .O(N__3159),
            .I(N__3156));
    Span12Mux_h I__469 (
            .O(N__3156),
            .I(N__3153));
    Odrv12 I__468 (
            .O(N__3153),
            .I(\U409_ADDRESS_DECODE.HIROMZ0 ));
    InMux I__467 (
            .O(N__3150),
            .I(N__3147));
    LocalMux I__466 (
            .O(N__3147),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    CascadeMux I__465 (
            .O(N__3144),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_));
    IoInMux I__464 (
            .O(N__3141),
            .I(N__3138));
    LocalMux I__463 (
            .O(N__3138),
            .I(N__3135));
    Span4Mux_s0_v I__462 (
            .O(N__3135),
            .I(N__3132));
    Span4Mux_v I__461 (
            .O(N__3132),
            .I(N__3129));
    Sp12to4 I__460 (
            .O(N__3129),
            .I(N__3126));
    Span12Mux_h I__459 (
            .O(N__3126),
            .I(N__3123));
    Odrv12 I__458 (
            .O(N__3123),
            .I(ROMENm_i));
    CascadeMux I__457 (
            .O(N__3120),
            .I(\U409_TICK.TICK603_11_cascade_ ));
    CascadeMux I__456 (
            .O(N__3117),
            .I(\U409_TRANSFER_ACK.m9_bm_cascade_ ));
    InMux I__455 (
            .O(N__3114),
            .I(N__3111));
    LocalMux I__454 (
            .O(N__3111),
            .I(\U409_TRANSFER_ACK.N_4 ));
    CascadeMux I__453 (
            .O(N__3108),
            .I(N__3104));
    CascadeMux I__452 (
            .O(N__3107),
            .I(N__3101));
    InMux I__451 (
            .O(N__3104),
            .I(N__3093));
    InMux I__450 (
            .O(N__3101),
            .I(N__3093));
    InMux I__449 (
            .O(N__3100),
            .I(N__3093));
    LocalMux I__448 (
            .O(N__3093),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__447 (
            .O(N__3090),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    InMux I__446 (
            .O(N__3087),
            .I(N__3084));
    LocalMux I__445 (
            .O(N__3084),
            .I(\U409_TRANSFER_ACK.m9_am ));
    InMux I__444 (
            .O(N__3081),
            .I(N__3077));
    InMux I__443 (
            .O(N__3080),
            .I(N__3074));
    LocalMux I__442 (
            .O(N__3077),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__441 (
            .O(N__3074),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__440 (
            .O(N__3069),
            .I(N__3064));
    InMux I__439 (
            .O(N__3068),
            .I(N__3059));
    InMux I__438 (
            .O(N__3067),
            .I(N__3059));
    LocalMux I__437 (
            .O(N__3064),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__436 (
            .O(N__3059),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__435 (
            .O(N__3054),
            .I(N__3048));
    InMux I__434 (
            .O(N__3053),
            .I(N__3040));
    InMux I__433 (
            .O(N__3052),
            .I(N__3040));
    InMux I__432 (
            .O(N__3051),
            .I(N__3040));
    LocalMux I__431 (
            .O(N__3048),
            .I(N__3037));
    InMux I__430 (
            .O(N__3047),
            .I(N__3034));
    LocalMux I__429 (
            .O(N__3040),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    Odrv4 I__428 (
            .O(N__3037),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__427 (
            .O(N__3034),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__426 (
            .O(N__3027),
            .I(N__3023));
    InMux I__425 (
            .O(N__3026),
            .I(N__3020));
    LocalMux I__424 (
            .O(N__3023),
            .I(\U409_TRANSFER_ACK.N_97 ));
    LocalMux I__423 (
            .O(N__3020),
            .I(\U409_TRANSFER_ACK.N_97 ));
    CascadeMux I__422 (
            .O(N__3015),
            .I(N__3012));
    InMux I__421 (
            .O(N__3012),
            .I(N__3008));
    InMux I__420 (
            .O(N__3011),
            .I(N__3003));
    LocalMux I__419 (
            .O(N__3008),
            .I(N__3000));
    InMux I__418 (
            .O(N__3007),
            .I(N__2995));
    InMux I__417 (
            .O(N__3006),
            .I(N__2995));
    LocalMux I__416 (
            .O(N__3003),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    Odrv4 I__415 (
            .O(N__3000),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__414 (
            .O(N__2995),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__413 (
            .O(N__2988),
            .I(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ));
    CascadeMux I__412 (
            .O(N__2985),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ));
    InMux I__411 (
            .O(N__2982),
            .I(N__2979));
    LocalMux I__410 (
            .O(N__2979),
            .I(N__2976));
    Odrv12 I__409 (
            .O(N__2976),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    IoInMux I__408 (
            .O(N__2973),
            .I(N__2970));
    LocalMux I__407 (
            .O(N__2970),
            .I(N__2967));
    IoSpan4Mux I__406 (
            .O(N__2967),
            .I(N__2964));
    Span4Mux_s0_v I__405 (
            .O(N__2964),
            .I(N__2961));
    Span4Mux_v I__404 (
            .O(N__2961),
            .I(N__2958));
    Sp12to4 I__403 (
            .O(N__2958),
            .I(N__2955));
    Odrv12 I__402 (
            .O(N__2955),
            .I(PORTSIZE_0_i));
    InMux I__401 (
            .O(N__2952),
            .I(N__2949));
    LocalMux I__400 (
            .O(N__2949),
            .I(N__2946));
    Span4Mux_v I__399 (
            .O(N__2946),
            .I(N__2942));
    InMux I__398 (
            .O(N__2945),
            .I(N__2939));
    Sp12to4 I__397 (
            .O(N__2942),
            .I(N__2934));
    LocalMux I__396 (
            .O(N__2939),
            .I(N__2934));
    Odrv12 I__395 (
            .O(N__2934),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    CascadeMux I__394 (
            .O(N__2931),
            .I(N__2925));
    InMux I__393 (
            .O(N__2930),
            .I(N__2918));
    InMux I__392 (
            .O(N__2929),
            .I(N__2918));
    InMux I__391 (
            .O(N__2928),
            .I(N__2915));
    InMux I__390 (
            .O(N__2925),
            .I(N__2910));
    InMux I__389 (
            .O(N__2924),
            .I(N__2910));
    InMux I__388 (
            .O(N__2923),
            .I(N__2907));
    LocalMux I__387 (
            .O(N__2918),
            .I(N__2902));
    LocalMux I__386 (
            .O(N__2915),
            .I(N__2902));
    LocalMux I__385 (
            .O(N__2910),
            .I(N__2899));
    LocalMux I__384 (
            .O(N__2907),
            .I(N__2896));
    Span4Mux_v I__383 (
            .O(N__2902),
            .I(N__2893));
    Span4Mux_v I__382 (
            .O(N__2899),
            .I(N__2890));
    Span4Mux_v I__381 (
            .O(N__2896),
            .I(N__2887));
    Sp12to4 I__380 (
            .O(N__2893),
            .I(N__2884));
    Span4Mux_h I__379 (
            .O(N__2890),
            .I(N__2881));
    Span4Mux_h I__378 (
            .O(N__2887),
            .I(N__2878));
    Odrv12 I__377 (
            .O(N__2884),
            .I(A_c_23));
    Odrv4 I__376 (
            .O(N__2881),
            .I(A_c_23));
    Odrv4 I__375 (
            .O(N__2878),
            .I(A_c_23));
    IoInMux I__374 (
            .O(N__2871),
            .I(N__2868));
    LocalMux I__373 (
            .O(N__2868),
            .I(N__2865));
    IoSpan4Mux I__372 (
            .O(N__2865),
            .I(N__2862));
    IoSpan4Mux I__371 (
            .O(N__2862),
            .I(N__2859));
    Span4Mux_s2_v I__370 (
            .O(N__2859),
            .I(N__2856));
    Sp12to4 I__369 (
            .O(N__2856),
            .I(N__2853));
    Span12Mux_v I__368 (
            .O(N__2853),
            .I(N__2850));
    Odrv12 I__367 (
            .O(N__2850),
            .I(U409_ADDRESS_DECODE_un1_nREGSPACE_i));
    CascadeMux I__366 (
            .O(N__2847),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    CascadeMux I__365 (
            .O(N__2844),
            .I(\U409_CIA.g0Z0Z_2_cascade_ ));
    InMux I__364 (
            .O(N__2841),
            .I(N__2835));
    InMux I__363 (
            .O(N__2840),
            .I(N__2835));
    LocalMux I__362 (
            .O(N__2835),
            .I(N__2832));
    Span4Mux_v I__361 (
            .O(N__2832),
            .I(N__2829));
    Span4Mux_h I__360 (
            .O(N__2829),
            .I(N__2826));
    Odrv4 I__359 (
            .O(N__2826),
            .I(A_c_30));
    InMux I__358 (
            .O(N__2823),
            .I(N__2817));
    InMux I__357 (
            .O(N__2822),
            .I(N__2817));
    LocalMux I__356 (
            .O(N__2817),
            .I(N__2814));
    Span4Mux_v I__355 (
            .O(N__2814),
            .I(N__2811));
    Span4Mux_v I__354 (
            .O(N__2811),
            .I(N__2808));
    Sp12to4 I__353 (
            .O(N__2808),
            .I(N__2805));
    Odrv12 I__352 (
            .O(N__2805),
            .I(A_c_28));
    InMux I__351 (
            .O(N__2802),
            .I(N__2796));
    InMux I__350 (
            .O(N__2801),
            .I(N__2796));
    LocalMux I__349 (
            .O(N__2796),
            .I(N__2793));
    Span4Mux_h I__348 (
            .O(N__2793),
            .I(N__2790));
    Span4Mux_v I__347 (
            .O(N__2790),
            .I(N__2787));
    Odrv4 I__346 (
            .O(N__2787),
            .I(A_c_29));
    CascadeMux I__345 (
            .O(N__2784),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ));
    InMux I__344 (
            .O(N__2781),
            .I(N__2778));
    LocalMux I__343 (
            .O(N__2778),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    InMux I__342 (
            .O(N__2775),
            .I(N__2769));
    InMux I__341 (
            .O(N__2774),
            .I(N__2769));
    LocalMux I__340 (
            .O(N__2769),
            .I(N__2766));
    Span4Mux_h I__339 (
            .O(N__2766),
            .I(N__2763));
    Span4Mux_v I__338 (
            .O(N__2763),
            .I(N__2760));
    Odrv4 I__337 (
            .O(N__2760),
            .I(A_c_24));
    CascadeMux I__336 (
            .O(N__2757),
            .I(N__2753));
    InMux I__335 (
            .O(N__2756),
            .I(N__2748));
    InMux I__334 (
            .O(N__2753),
            .I(N__2748));
    LocalMux I__333 (
            .O(N__2748),
            .I(N__2745));
    Span4Mux_v I__332 (
            .O(N__2745),
            .I(N__2742));
    Span4Mux_v I__331 (
            .O(N__2742),
            .I(N__2739));
    Sp12to4 I__330 (
            .O(N__2739),
            .I(N__2736));
    Odrv12 I__329 (
            .O(N__2736),
            .I(A_c_26));
    CascadeMux I__328 (
            .O(N__2733),
            .I(N__2730));
    InMux I__327 (
            .O(N__2730),
            .I(N__2724));
    InMux I__326 (
            .O(N__2729),
            .I(N__2724));
    LocalMux I__325 (
            .O(N__2724),
            .I(N__2721));
    Span4Mux_v I__324 (
            .O(N__2721),
            .I(N__2718));
    Sp12to4 I__323 (
            .O(N__2718),
            .I(N__2715));
    Odrv12 I__322 (
            .O(N__2715),
            .I(A_c_31));
    InMux I__321 (
            .O(N__2712),
            .I(N__2708));
    InMux I__320 (
            .O(N__2711),
            .I(N__2705));
    LocalMux I__319 (
            .O(N__2708),
            .I(N__2700));
    LocalMux I__318 (
            .O(N__2705),
            .I(N__2700));
    Span4Mux_v I__317 (
            .O(N__2700),
            .I(N__2697));
    Span4Mux_h I__316 (
            .O(N__2697),
            .I(N__2694));
    Odrv4 I__315 (
            .O(N__2694),
            .I(A_c_27));
    InMux I__314 (
            .O(N__2691),
            .I(N__2688));
    LocalMux I__313 (
            .O(N__2688),
            .I(\U409_CIA.g0Z0Z_10 ));
    InMux I__312 (
            .O(N__2685),
            .I(N__2674));
    InMux I__311 (
            .O(N__2684),
            .I(N__2674));
    InMux I__310 (
            .O(N__2683),
            .I(N__2674));
    InMux I__309 (
            .O(N__2682),
            .I(N__2671));
    InMux I__308 (
            .O(N__2681),
            .I(N__2668));
    LocalMux I__307 (
            .O(N__2674),
            .I(N__2665));
    LocalMux I__306 (
            .O(N__2671),
            .I(N__2662));
    LocalMux I__305 (
            .O(N__2668),
            .I(N__2655));
    Sp12to4 I__304 (
            .O(N__2665),
            .I(N__2655));
    Sp12to4 I__303 (
            .O(N__2662),
            .I(N__2655));
    Span12Mux_v I__302 (
            .O(N__2655),
            .I(N__2652));
    Odrv12 I__301 (
            .O(N__2652),
            .I(A_c_22));
    InMux I__300 (
            .O(N__2649),
            .I(N__2641));
    InMux I__299 (
            .O(N__2648),
            .I(N__2641));
    InMux I__298 (
            .O(N__2647),
            .I(N__2636));
    InMux I__297 (
            .O(N__2646),
            .I(N__2636));
    LocalMux I__296 (
            .O(N__2641),
            .I(N__2633));
    LocalMux I__295 (
            .O(N__2636),
            .I(N__2630));
    Span4Mux_v I__294 (
            .O(N__2633),
            .I(N__2627));
    Span12Mux_v I__293 (
            .O(N__2630),
            .I(N__2624));
    Span4Mux_h I__292 (
            .O(N__2627),
            .I(N__2621));
    Odrv12 I__291 (
            .O(N__2624),
            .I(A_c_21));
    Odrv4 I__290 (
            .O(N__2621),
            .I(A_c_21));
    CascadeMux I__289 (
            .O(N__2616),
            .I(N__2613));
    InMux I__288 (
            .O(N__2613),
            .I(N__2610));
    LocalMux I__287 (
            .O(N__2610),
            .I(N__2607));
    Span4Mux_v I__286 (
            .O(N__2607),
            .I(N__2604));
    Odrv4 I__285 (
            .O(N__2604),
            .I(\U409_CIA.g0Z0Z_8 ));
    CascadeMux I__284 (
            .O(N__2601),
            .I(N__2598));
    InMux I__283 (
            .O(N__2598),
            .I(N__2592));
    InMux I__282 (
            .O(N__2597),
            .I(N__2592));
    LocalMux I__281 (
            .O(N__2592),
            .I(N__2589));
    Span4Mux_v I__280 (
            .O(N__2589),
            .I(N__2586));
    Span4Mux_h I__279 (
            .O(N__2586),
            .I(N__2583));
    Span4Mux_v I__278 (
            .O(N__2583),
            .I(N__2580));
    Odrv4 I__277 (
            .O(N__2580),
            .I(A_c_16));
    CascadeMux I__276 (
            .O(N__2577),
            .I(N__2573));
    InMux I__275 (
            .O(N__2576),
            .I(N__2570));
    InMux I__274 (
            .O(N__2573),
            .I(N__2567));
    LocalMux I__273 (
            .O(N__2570),
            .I(N__2564));
    LocalMux I__272 (
            .O(N__2567),
            .I(N__2561));
    Span4Mux_v I__271 (
            .O(N__2564),
            .I(N__2556));
    Span4Mux_v I__270 (
            .O(N__2561),
            .I(N__2556));
    Span4Mux_h I__269 (
            .O(N__2556),
            .I(N__2553));
    Span4Mux_v I__268 (
            .O(N__2553),
            .I(N__2550));
    Span4Mux_v I__267 (
            .O(N__2550),
            .I(N__2547));
    Odrv4 I__266 (
            .O(N__2547),
            .I(A_c_18));
    InMux I__265 (
            .O(N__2544),
            .I(N__2541));
    LocalMux I__264 (
            .O(N__2541),
            .I(\U409_CIA.g0Z0Z_11 ));
    InMux I__263 (
            .O(N__2538),
            .I(N__2534));
    InMux I__262 (
            .O(N__2537),
            .I(N__2531));
    LocalMux I__261 (
            .O(N__2534),
            .I(N__2526));
    LocalMux I__260 (
            .O(N__2531),
            .I(N__2526));
    Sp12to4 I__259 (
            .O(N__2526),
            .I(N__2523));
    Span12Mux_v I__258 (
            .O(N__2523),
            .I(N__2520));
    Odrv12 I__257 (
            .O(N__2520),
            .I(A_c_17));
    CascadeMux I__256 (
            .O(N__2517),
            .I(\U409_ADDRESS_DECODE.HIROM_0_cascade_ ));
    InMux I__255 (
            .O(N__2514),
            .I(N__2511));
    LocalMux I__254 (
            .O(N__2511),
            .I(N__2508));
    Span4Mux_v I__253 (
            .O(N__2508),
            .I(N__2505));
    Span4Mux_v I__252 (
            .O(N__2505),
            .I(N__2500));
    InMux I__251 (
            .O(N__2504),
            .I(N__2495));
    InMux I__250 (
            .O(N__2503),
            .I(N__2495));
    Sp12to4 I__249 (
            .O(N__2500),
            .I(N__2492));
    LocalMux I__248 (
            .O(N__2495),
            .I(N__2489));
    Span12Mux_s3_h I__247 (
            .O(N__2492),
            .I(N__2484));
    Span12Mux_h I__246 (
            .O(N__2489),
            .I(N__2484));
    Span12Mux_v I__245 (
            .O(N__2484),
            .I(N__2481));
    Odrv12 I__244 (
            .O(N__2481),
            .I(A_c_19));
    CascadeMux I__243 (
            .O(N__2478),
            .I(N__2475));
    InMux I__242 (
            .O(N__2475),
            .I(N__2472));
    LocalMux I__241 (
            .O(N__2472),
            .I(\U409_ADDRESS_DECODE.HIROM_0 ));
    InMux I__240 (
            .O(N__2469),
            .I(N__2466));
    LocalMux I__239 (
            .O(N__2466),
            .I(N__2463));
    Span4Mux_h I__238 (
            .O(N__2463),
            .I(N__2460));
    Span4Mux_v I__237 (
            .O(N__2460),
            .I(N__2455));
    InMux I__236 (
            .O(N__2459),
            .I(N__2450));
    InMux I__235 (
            .O(N__2458),
            .I(N__2450));
    Sp12to4 I__234 (
            .O(N__2455),
            .I(N__2445));
    LocalMux I__233 (
            .O(N__2450),
            .I(N__2445));
    Odrv12 I__232 (
            .O(N__2445),
            .I(A_c_20));
    CascadeMux I__231 (
            .O(N__2442),
            .I(N__2439));
    InMux I__230 (
            .O(N__2439),
            .I(N__2436));
    LocalMux I__229 (
            .O(N__2436),
            .I(N__2432));
    InMux I__228 (
            .O(N__2435),
            .I(N__2429));
    Sp12to4 I__227 (
            .O(N__2432),
            .I(N__2424));
    LocalMux I__226 (
            .O(N__2429),
            .I(N__2424));
    Odrv12 I__225 (
            .O(N__2424),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    InMux I__224 (
            .O(N__2421),
            .I(N__2418));
    LocalMux I__223 (
            .O(N__2418),
            .I(N__2415));
    Span4Mux_v I__222 (
            .O(N__2415),
            .I(N__2411));
    InMux I__221 (
            .O(N__2414),
            .I(N__2408));
    Span4Mux_v I__220 (
            .O(N__2411),
            .I(N__2405));
    LocalMux I__219 (
            .O(N__2408),
            .I(N__2402));
    Span4Mux_v I__218 (
            .O(N__2405),
            .I(N__2397));
    Span4Mux_v I__217 (
            .O(N__2402),
            .I(N__2397));
    Span4Mux_h I__216 (
            .O(N__2397),
            .I(N__2394));
    Odrv4 I__215 (
            .O(N__2394),
            .I(A_c_25));
    ClkMux I__214 (
            .O(N__2391),
            .I(N__2364));
    ClkMux I__213 (
            .O(N__2390),
            .I(N__2364));
    ClkMux I__212 (
            .O(N__2389),
            .I(N__2364));
    ClkMux I__211 (
            .O(N__2388),
            .I(N__2364));
    ClkMux I__210 (
            .O(N__2387),
            .I(N__2364));
    ClkMux I__209 (
            .O(N__2386),
            .I(N__2364));
    ClkMux I__208 (
            .O(N__2385),
            .I(N__2364));
    ClkMux I__207 (
            .O(N__2384),
            .I(N__2364));
    ClkMux I__206 (
            .O(N__2383),
            .I(N__2364));
    GlobalMux I__205 (
            .O(N__2364),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2389));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2386));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__2390));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2388));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .I(N__2385));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2383));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2391));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2387));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__2384));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_7_0  (
            .in0(N__2597),
            .in1(N__2503),
            .in2(N__2577),
            .in3(N__2537),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_7_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_7_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_7_2  (
            .in0(N__2421),
            .in1(N__2504),
            .in2(N__2601),
            .in3(N__2576),
            .lcout(\U409_CIA.g0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_1_8_4 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_1_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_1_8_4  (
            .in0(N__2544),
            .in1(N__2469),
            .in2(N__2616),
            .in3(N__2538),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__2648),
            .in2(_gnd_net_),
            .in3(N__2458),
            .lcout(\U409_ADDRESS_DECODE.HIROM_0 ),
            .ltout(\U409_ADDRESS_DECODE.HIROM_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_1_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_1_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_1_12_2  (
            .in0(N__2923),
            .in1(N__2684),
            .in2(N__2517),
            .in3(N__2514),
            .lcout(\U409_ADDRESS_DECODE.HIROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_5  (
            .in0(N__2683),
            .in1(N__4475),
            .in2(N__2478),
            .in3(N__2435),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_12_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_12_7  (
            .in0(N__2685),
            .in1(N__2459),
            .in2(N__2442),
            .in3(N__2649),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0  (
            .in0(N__2414),
            .in1(N__2711),
            .in2(N__2757),
            .in3(N__2774),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_17_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_17_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.g0_2_LC_1_17_1  (
            .in0(N__2802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2841),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_17_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_17_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_CIA.g0_13_LC_1_17_2  (
            .in0(N__2823),
            .in1(N__2691),
            .in2(N__2844),
            .in3(N__2682),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_3  (
            .in0(N__2729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2840),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_4  (
            .in0(N__2822),
            .in1(N__2801),
            .in2(N__2784),
            .in3(N__2781),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_17_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_17_5  (
            .in0(N__2775),
            .in1(N__2756),
            .in2(N__2733),
            .in3(N__2712),
            .lcout(\U409_CIA.g0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_2_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_2_12_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_2_12_0  (
            .in0(N__2681),
            .in1(N__2924),
            .in2(_gnd_net_),
            .in3(N__2646),
            .lcout(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_2_12_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_2_12_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_CIA.g0_8_LC_2_12_5  (
            .in0(N__2647),
            .in1(_gnd_net_),
            .in2(N__2931),
            .in3(N__5469),
            .lcout(\U409_CIA.g0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_12_2  (
            .in0(N__2930),
            .in1(N__2945),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_3  (
            .in0(N__5468),
            .in1(N__2929),
            .in2(N__2985),
            .in3(N__2982),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_7_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_7_13_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_7_13_5  (
            .in0(N__2952),
            .in1(N__2928),
            .in2(_gnd_net_),
            .in3(N__4516),
            .lcout(U409_ADDRESS_DECODE_un1_nREGSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_9_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_9_6_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_9_6_1  (
            .in0(N__3953),
            .in1(N__3918),
            .in2(N__3996),
            .in3(N__3336),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_9_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_9_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_9_6_7  (
            .in0(N__3952),
            .in1(N__3917),
            .in2(N__3995),
            .in3(N__3504),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_7_7  (
            .in0(N__5429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_2  (
            .in0(N__5470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3474),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_9_0 .LUT_INIT=16'b0000010100110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_9_0  (
            .in0(N__3473),
            .in1(N__3114),
            .in2(N__3108),
            .in3(N__3051),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_9_1 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_9_1  (
            .in0(N__3052),
            .in1(N__5472),
            .in2(N__2847),
            .in3(N__3011),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_9_9_2  (
            .in0(N__5474),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3068),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_9_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_9_9_3  (
            .in0(N__4307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5473),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_9_4 .LUT_INIT=16'b0000010000110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_9_4  (
            .in0(N__3472),
            .in1(N__3007),
            .in2(N__3107),
            .in3(N__3027),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_9_5 .LUT_INIT=16'b0000100001001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_9_5  (
            .in0(N__3053),
            .in1(N__5471),
            .in2(N__3117),
            .in3(N__3087),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__3080),
            .in2(_gnd_net_),
            .in3(N__3067),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_9_7 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_9_7  (
            .in0(N__3006),
            .in1(N__3100),
            .in2(N__3090),
            .in3(N__3471),
            .lcout(\U409_TRANSFER_ACK.m9_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_10_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_10_4  (
            .in0(N__3047),
            .in1(N__3081),
            .in2(N__3651),
            .in3(N__3069),
            .lcout(\U409_TRANSFER_ACK.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_11_0 .LUT_INIT=16'b0001101100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_11_0  (
            .in0(N__3054),
            .in1(N__3026),
            .in2(N__3015),
            .in3(N__3546),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_11_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__5475),
            .in2(N__2988),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_11_2 .LUT_INIT=16'b0111000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_11_2  (
            .in0(N__3184),
            .in1(N__3200),
            .in2(N__5486),
            .in3(N__3216),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_11_3  (
            .in0(N__3150),
            .in1(N__5480),
            .in2(N__4530),
            .in3(N__3691),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_11_4  (
            .in0(N__3640),
            .in1(N__3179),
            .in2(N__3219),
            .in3(N__3198),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_11_5 .LUT_INIT=16'b1010000110100101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_11_5  (
            .in0(N__3199),
            .in1(N__3210),
            .in2(N__3186),
            .in3(N__3641),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_11_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_11_6  (
            .in0(N__5481),
            .in1(N__3183),
            .in2(N__3204),
            .in3(N__3531),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_11_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_11_7  (
            .in0(N__3201),
            .in1(N__5479),
            .in2(_gnd_net_),
            .in3(N__3185),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_9_12_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ROMEN_LC_9_12_1  (
            .in0(N__4449),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__3162),
            .lcout(U409_ADDRESS_DECODE_un1_ROMEN_0),
            .ltout(U409_ADDRESS_DECODE_un1_ROMEN_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_12_2 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_9_12_2  (
            .in0(N__4526),
            .in1(_gnd_net_),
            .in2(N__3144),
            .in3(N__5487),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_0  (
            .in0(N__3306),
            .in1(N__3249),
            .in2(N__4056),
            .in3(N__3489),
            .lcout(),
            .ltout(\U409_TICK.TICK603_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_1  (
            .in0(N__3255),
            .in1(N__3324),
            .in2(N__3120),
            .in3(N__3234),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_10_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_10_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_10_5_2  (
            .in0(N__3981),
            .in1(N__3948),
            .in2(N__3288),
            .in3(N__3426),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_3  (
            .in0(N__3348),
            .in1(N__3372),
            .in2(N__3402),
            .in3(N__3516),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_10_5_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_10_5_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_10_5_4  (
            .in0(N__3985),
            .in1(N__3920),
            .in2(N__3285),
            .in3(N__3266),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_10_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_10_5_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_10_5_5  (
            .in0(N__3950),
            .in1(N__3910),
            .in2(N__3360),
            .in3(N__3986),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_10_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_10_5_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_10_5_6  (
            .in0(N__3909),
            .in1(N__3949),
            .in2(N__3994),
            .in3(N__3384),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_7  (
            .in0(N__3417),
            .in1(N__3438),
            .in2(_gnd_net_),
            .in3(N__4087),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__4051),
            .in2(N__4086),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__3248),
            .in2(_gnd_net_),
            .in3(N__3237),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__3233),
            .in2(_gnd_net_),
            .in3(N__3222),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__3437),
            .in2(_gnd_net_),
            .in3(N__3420),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__3416),
            .in2(_gnd_net_),
            .in3(N__3405),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3401),
            .in3(N__3378),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__4019),
            .in2(_gnd_net_),
            .in3(N__3375),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__3371),
            .in2(_gnd_net_),
            .in3(N__3351),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__3347),
            .in2(_gnd_net_),
            .in3(N__3330),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__4007),
            .in2(_gnd_net_),
            .in3(N__3327),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__5130),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__3320),
            .in2(_gnd_net_),
            .in3(N__3309),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__5130),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__3305),
            .in2(_gnd_net_),
            .in3(N__3291),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__5130),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__4034),
            .in2(_gnd_net_),
            .in3(N__3519),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__5130),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__3515),
            .in2(_gnd_net_),
            .in3(N__3498),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__3872),
            .in2(_gnd_net_),
            .in3(N__3495),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__3488),
            .in2(_gnd_net_),
            .in3(N__3492),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5130),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_8_1 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_8_1  (
            .in0(N__4200),
            .in1(N__4183),
            .in2(N__4141),
            .in3(N__4166),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__3456));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_0  (
            .in0(N__4276),
            .in1(N__4720),
            .in2(_gnd_net_),
            .in3(N__4771),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_1 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__4682),
            .in2(N__3444),
            .in3(N__4256),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__5334));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_5 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_5  (
            .in0(N__3653),
            .in1(N__4784),
            .in2(N__3699),
            .in3(N__4621),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_6 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__4287),
            .in2(N__3441),
            .in3(N__4746),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__5334));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0  (
            .in0(N__4623),
            .in1(N__3695),
            .in2(N__3652),
            .in3(N__4657),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1  (
            .in0(N__3558),
            .in1(N__4622),
            .in2(_gnd_net_),
            .in3(N__4785),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_2  (
            .in0(N__4277),
            .in1(N__4772),
            .in2(_gnd_net_),
            .in3(N__4257),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_3  (
            .in0(N__4658),
            .in1(N__4583),
            .in2(_gnd_net_),
            .in3(N__4608),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_4 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_4  (
            .in0(N__4725),
            .in1(N__4773),
            .in2(N__4281),
            .in3(N__4258),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_10_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_10_5  (
            .in0(N__4698),
            .in1(N__3564),
            .in2(N__4263),
            .in3(N__4683),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5327));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_11_0  (
            .in0(N__5462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4551),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2  (
            .in0(N__3557),
            .in1(N__3545),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_11_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_11_3  (
            .in0(N__3802),
            .in1(N__3814),
            .in2(N__3534),
            .in3(N__3530),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_11_4 .LUT_INIT=16'b0100111001001100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_10_11_4  (
            .in0(N__5467),
            .in1(N__3827),
            .in2(N__3849),
            .in3(N__3804),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_11_5 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_11_5  (
            .in0(N__3803),
            .in1(N__3815),
            .in2(_gnd_net_),
            .in3(N__5466),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_11_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_11_6  (
            .in0(N__3816),
            .in1(_gnd_net_),
            .in2(N__5485),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_12_5 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_12_5  (
            .in0(N__4448),
            .in1(N__4524),
            .in2(N__3792),
            .in3(N__4409),
            .lcout(nBUFEN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_11_4_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_11_4_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_11_4_2  (
            .in0(N__4104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3780),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_11_4_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_11_4_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__4103),
            .in2(_gnd_net_),
            .in3(N__3738),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_11_5_6 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_11_5_6  (
            .in0(N__3951),
            .in1(N__3921),
            .in2(N__4092),
            .in3(N__3987),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_11_6_0  (
            .in0(N__5171),
            .in1(N__5273),
            .in2(N__5235),
            .in3(N__4854),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_11_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_11_6_1  (
            .in0(N__4956),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4937),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_2  (
            .in0(N__4914),
            .in1(N__4803),
            .in2(N__4992),
            .in3(N__4955),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_11_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_11_6_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_11_6_3  (
            .in0(N__5274),
            .in1(N__5173),
            .in2(N__5229),
            .in3(N__4830),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_11_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_11_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__4091),
            .in2(_gnd_net_),
            .in3(N__4055),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_11_6_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_11_6_5  (
            .in0(N__5272),
            .in1(N__5172),
            .in2(N__5228),
            .in3(N__4936),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6  (
            .in0(N__4035),
            .in1(N__3873),
            .in2(N__4023),
            .in3(N__4008),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_11_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_11_6_7  (
            .in0(N__3954),
            .in1(N__3919),
            .in2(N__3882),
            .in3(N__3879),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_11_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_11_7_0  (
            .in0(N__5177),
            .in1(N__5269),
            .in2(N__5227),
            .in3(N__5046),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_1  (
            .in0(N__4866),
            .in1(N__4896),
            .in2(_gnd_net_),
            .in3(N__4935),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_2  (
            .in0(N__3861),
            .in1(N__5037),
            .in2(N__3852),
            .in3(N__5076),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_11_7_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_11_7_3  (
            .in0(N__5271),
            .in1(N__5207),
            .in2(N__4236),
            .in3(N__4217),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_5  (
            .in0(N__5019),
            .in1(N__4881),
            .in2(N__4821),
            .in3(N__4968),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6  (
            .in0(N__5295),
            .in1(N__5142),
            .in2(N__5061),
            .in3(N__4844),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_11_7_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_11_7_7  (
            .in0(N__5270),
            .in1(N__5178),
            .in2(N__4206),
            .in3(N__5007),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5127),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_11_8_0  (
            .in0(N__5603),
            .in1(N__5648),
            .in2(_gnd_net_),
            .in3(N__5682),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_11_8_1 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_11_8_1  (
            .in0(N__4161),
            .in1(N__5604),
            .in2(N__4203),
            .in3(N__4344),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5574),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_11_8_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_11_8_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_11_8_4  (
            .in0(N__4184),
            .in1(N__4162),
            .in2(N__4146),
            .in3(N__4198),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5574),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_8_7 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_8_7  (
            .in0(N__4199),
            .in1(N__4185),
            .in2(N__4167),
            .in3(N__4145),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5645),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5573),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_1  (
            .in0(N__5697),
            .in1(N__5718),
            .in2(_gnd_net_),
            .in3(N__5739),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__5647),
            .in2(_gnd_net_),
            .in3(N__5680),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5573),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_11_9_3  (
            .in0(N__5698),
            .in1(N__5602),
            .in2(N__5745),
            .in3(N__5719),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_11_9_4  (
            .in0(N__5601),
            .in1(N__5644),
            .in2(_gnd_net_),
            .in3(N__5679),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__4300),
            .in2(N__4347),
            .in3(N__4343),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_11_9_6  (
            .in0(N__4332),
            .in1(N__5646),
            .in2(N__4326),
            .in3(N__5681),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5573),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_9_7  (
            .in0(N__4656),
            .in1(N__4582),
            .in2(_gnd_net_),
            .in3(N__4607),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_10_0  (
            .in0(N__4605),
            .in1(N__4745),
            .in2(N__4584),
            .in3(N__4654),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_2  (
            .in0(N__4606),
            .in1(N__4655),
            .in2(_gnd_net_),
            .in3(N__4262),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5326));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_10_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_10_3  (
            .in0(N__4680),
            .in1(N__4744),
            .in2(N__4659),
            .in3(N__4696),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_10_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_10_4  (
            .in0(N__4770),
            .in1(N__4719),
            .in2(N__4788),
            .in3(N__4559),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_10_5  (
            .in0(N__4769),
            .in1(N__4743),
            .in2(N__4724),
            .in3(N__4697),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_10_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_10_6  (
            .in0(N__4681),
            .in1(N__4653),
            .in2(N__4626),
            .in3(N__4560),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_10_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__4604),
            .in2(_gnd_net_),
            .in3(N__4578),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_11_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__5403),
            .in2(_gnd_net_),
            .in3(N__4550),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__4539),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_12_1 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_12_1  (
            .in0(N__4525),
            .in1(N__4447),
            .in2(_gnd_net_),
            .in3(N__4410),
            .lcout(U409_ADDRESS_DECODE_un1_nRAMSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__4949),
            .in2(N__4938),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__4910),
            .in2(_gnd_net_),
            .in3(N__4899),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__4895),
            .in2(_gnd_net_),
            .in3(N__4884),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__4880),
            .in2(_gnd_net_),
            .in3(N__4869),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__4865),
            .in2(_gnd_net_),
            .in3(N__4848),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4845),
            .in3(N__4824),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__4817),
            .in2(_gnd_net_),
            .in3(N__4806),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__4802),
            .in2(_gnd_net_),
            .in3(N__4791),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__5141),
            .in2(_gnd_net_),
            .in3(N__5079),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__5075),
            .in2(_gnd_net_),
            .in3(N__5064),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__5057),
            .in2(_gnd_net_),
            .in3(N__5040),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__5036),
            .in2(_gnd_net_),
            .in3(N__5025),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__5288),
            .in2(_gnd_net_),
            .in3(N__5022),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__5018),
            .in2(_gnd_net_),
            .in3(N__5001),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__4967),
            .in2(_gnd_net_),
            .in3(N__4998),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__4991),
            .in2(_gnd_net_),
            .in3(N__4995),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_12_8_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_12_8_2  (
            .in0(N__5174),
            .in1(N__5276),
            .in2(N__4977),
            .in3(N__5223),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_12_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_12_8_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_12_8_3  (
            .in0(N__5275),
            .in1(N__5175),
            .in2(N__5230),
            .in3(N__5301),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_12_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_12_8_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_12_8_7  (
            .in0(N__5277),
            .in1(N__5241),
            .in2(N__5231),
            .in3(N__5176),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__5677),
            .in2(N__5649),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__5740),
            .in2(_gnd_net_),
            .in3(N__5094),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__5572),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__5598),
            .in2(_gnd_net_),
            .in3(N__5091),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__5699),
            .in2(_gnd_net_),
            .in3(N__5088),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__5572),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__5720),
            .in2(_gnd_net_),
            .in3(N__5085),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5  (
            .in0(N__5600),
            .in1(N__5642),
            .in2(N__5082),
            .in3(N__5655),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5572),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6  (
            .in0(N__5741),
            .in1(N__5721),
            .in2(N__5703),
            .in3(N__5678),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .LUT_INIT=16'b0001010110101010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7  (
            .in0(N__5599),
            .in1(N__5643),
            .in2(N__5613),
            .in3(N__5610),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5572),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_14_12_6.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_14_12_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_iobuf_RNO_LC_14_12_6 (
            .in0(N__5559),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_353_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_17_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_17_12_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_17_12_6  (
            .in0(N__5532),
            .in1(N__5504),
            .in2(_gnd_net_),
            .in3(N__5410),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 25 2025 11:06:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    A,
    TICK50,
    nROMEN,
    nCIACS1,
    TICK60,
    CLKCIA,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    TSn,
    nBUFEN,
    nREGSPACE,
    nRAMSPACE,
    RESETn,
    OVL,
    TACKn,
    nCIACS0,
    PORTSIZE);

    input [1:0] TT;
    input [31:1] A;
    output TICK50;
    output nROMEN;
    output nCIACS1;
    output TICK60;
    output CLKCIA;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    input TSn;
    output nBUFEN;
    output nREGSPACE;
    output nRAMSPACE;
    input RESETn;
    input OVL;
    inout TACKn;
    output nCIACS0;
    output PORTSIZE;

    wire N__6284;
    wire N__6283;
    wire N__6282;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6263;
    wire N__6262;
    wire N__6261;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6236;
    wire N__6235;
    wire N__6234;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6218;
    wire N__6217;
    wire N__6216;
    wire N__6209;
    wire N__6208;
    wire N__6207;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6191;
    wire N__6190;
    wire N__6189;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6155;
    wire N__6154;
    wire N__6153;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6119;
    wire N__6118;
    wire N__6117;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6101;
    wire N__6100;
    wire N__6099;
    wire N__6092;
    wire N__6091;
    wire N__6090;
    wire N__6083;
    wire N__6082;
    wire N__6081;
    wire N__6074;
    wire N__6073;
    wire N__6072;
    wire N__6065;
    wire N__6064;
    wire N__6063;
    wire N__6056;
    wire N__6055;
    wire N__6054;
    wire N__6047;
    wire N__6046;
    wire N__6045;
    wire N__6038;
    wire N__6037;
    wire N__6036;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6020;
    wire N__6019;
    wire N__6018;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5993;
    wire N__5992;
    wire N__5991;
    wire N__5984;
    wire N__5983;
    wire N__5982;
    wire N__5975;
    wire N__5974;
    wire N__5973;
    wire N__5966;
    wire N__5965;
    wire N__5964;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5929;
    wire N__5926;
    wire N__5925;
    wire N__5924;
    wire N__5917;
    wire N__5914;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5857;
    wire N__5856;
    wire N__5853;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5821;
    wire N__5818;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5804;
    wire N__5799;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5771;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5745;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5723;
    wire N__5718;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5637;
    wire N__5634;
    wire N__5633;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5613;
    wire N__5612;
    wire N__5607;
    wire N__5604;
    wire N__5599;
    wire N__5598;
    wire N__5597;
    wire N__5596;
    wire N__5589;
    wire N__5586;
    wire N__5581;
    wire N__5580;
    wire N__5579;
    wire N__5576;
    wire N__5575;
    wire N__5570;
    wire N__5565;
    wire N__5560;
    wire N__5559;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5494;
    wire N__5491;
    wire N__5490;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5473;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5461;
    wire N__5458;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5446;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5431;
    wire N__5428;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5416;
    wire N__5413;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5383;
    wire N__5380;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5323;
    wire N__5322;
    wire N__5321;
    wire N__5320;
    wire N__5319;
    wire N__5318;
    wire N__5317;
    wire N__5316;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5260;
    wire N__5257;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5224;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5188;
    wire N__5185;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5127;
    wire N__5120;
    wire N__5117;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5034;
    wire N__5033;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5018;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__5001;
    wire N__4996;
    wire N__4993;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4969;
    wire N__4966;
    wire N__4965;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4923;
    wire N__4920;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4910;
    wire N__4905;
    wire N__4900;
    wire N__4899;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4875;
    wire N__4874;
    wire N__4869;
    wire N__4866;
    wire N__4861;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4855;
    wire N__4848;
    wire N__4845;
    wire N__4840;
    wire N__4839;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4790;
    wire N__4787;
    wire N__4780;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4765;
    wire N__4758;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4735;
    wire N__4734;
    wire N__4729;
    wire N__4724;
    wire N__4721;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4707;
    wire N__4706;
    wire N__4701;
    wire N__4698;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4686;
    wire N__4685;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4673;
    wire N__4666;
    wire N__4665;
    wire N__4664;
    wire N__4663;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4639;
    wire N__4636;
    wire N__4635;
    wire N__4630;
    wire N__4627;
    wire N__4626;
    wire N__4625;
    wire N__4624;
    wire N__4623;
    wire N__4620;
    wire N__4611;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4589;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4536;
    wire N__4527;
    wire N__4522;
    wire N__4521;
    wire N__4518;
    wire N__4517;
    wire N__4516;
    wire N__4515;
    wire N__4514;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4496;
    wire N__4489;
    wire N__4488;
    wire N__4487;
    wire N__4486;
    wire N__4485;
    wire N__4484;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4472;
    wire N__4461;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4449;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4420;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4395;
    wire N__4394;
    wire N__4391;
    wire N__4390;
    wire N__4387;
    wire N__4386;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4368;
    wire N__4367;
    wire N__4364;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4290;
    wire N__4289;
    wire N__4286;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4268;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4253;
    wire N__4248;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4236;
    wire N__4235;
    wire N__4232;
    wire N__4227;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4209;
    wire N__4208;
    wire N__4205;
    wire N__4200;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4179;
    wire N__4178;
    wire N__4173;
    wire N__4170;
    wire N__4165;
    wire N__4162;
    wire N__4161;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4139;
    wire N__4134;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4108;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4095;
    wire N__4094;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4078;
    wire N__4075;
    wire N__4068;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4041;
    wire N__4036;
    wire N__4033;
    wire N__4032;
    wire N__4031;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4023;
    wire N__4022;
    wire N__4019;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3946;
    wire N__3945;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3861;
    wire N__3858;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3843;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3808;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3757;
    wire N__3754;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3742;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3706;
    wire N__3705;
    wire N__3704;
    wire N__3703;
    wire N__3702;
    wire N__3701;
    wire N__3700;
    wire N__3699;
    wire N__3690;
    wire N__3681;
    wire N__3676;
    wire N__3675;
    wire N__3674;
    wire N__3673;
    wire N__3672;
    wire N__3671;
    wire N__3668;
    wire N__3667;
    wire N__3666;
    wire N__3655;
    wire N__3652;
    wire N__3647;
    wire N__3644;
    wire N__3637;
    wire N__3636;
    wire N__3635;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3609;
    wire N__3606;
    wire N__3599;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3550;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3523;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3511;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3501;
    wire N__3496;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3466;
    wire N__3463;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3414;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3398;
    wire N__3395;
    wire N__3388;
    wire N__3387;
    wire N__3386;
    wire N__3381;
    wire N__3378;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3339;
    wire N__3338;
    wire N__3337;
    wire N__3332;
    wire N__3327;
    wire N__3322;
    wire N__3321;
    wire N__3320;
    wire N__3317;
    wire N__3316;
    wire N__3311;
    wire N__3306;
    wire N__3301;
    wire N__3300;
    wire N__3297;
    wire N__3296;
    wire N__3295;
    wire N__3292;
    wire N__3287;
    wire N__3284;
    wire N__3277;
    wire N__3276;
    wire N__3275;
    wire N__3274;
    wire N__3273;
    wire N__3272;
    wire N__3269;
    wire N__3262;
    wire N__3257;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3234;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3230;
    wire N__3229;
    wire N__3228;
    wire N__3225;
    wire N__3220;
    wire N__3217;
    wire N__3212;
    wire N__3205;
    wire N__3196;
    wire N__3195;
    wire N__3194;
    wire N__3193;
    wire N__3192;
    wire N__3191;
    wire N__3190;
    wire N__3187;
    wire N__3180;
    wire N__3173;
    wire N__3166;
    wire N__3163;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3048;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2949;
    wire N__2948;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2931;
    wire N__2930;
    wire N__2927;
    wire N__2922;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2901;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2884;
    wire N__2881;
    wire N__2880;
    wire N__2877;
    wire N__2876;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2853;
    wire N__2848;
    wire N__2845;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2833;
    wire N__2830;
    wire N__2829;
    wire N__2826;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2800;
    wire N__2799;
    wire N__2798;
    wire N__2795;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2753;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2700;
    wire N__2699;
    wire N__2696;
    wire N__2691;
    wire N__2686;
    wire N__2683;
    wire N__2682;
    wire N__2679;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2667;
    wire N__2662;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2649;
    wire N__2648;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2604;
    wire N__2603;
    wire N__2600;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2553;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2529;
    wire N__2526;
    wire N__2521;
    wire N__2518;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2505;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2473;
    wire N__2472;
    wire N__2471;
    wire N__2470;
    wire N__2469;
    wire N__2468;
    wire N__2467;
    wire N__2466;
    wire N__2465;
    wire N__2446;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_18;
    wire A_c_17;
    wire A_c_16;
    wire \U409_CIA.g0Z0Z_8_cascade_ ;
    wire \U409_CIA.g0Z0Z_11 ;
    wire A_c_25;
    wire A_c_24;
    wire A_c_26;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire TT_c_0;
    wire A_c_31;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ;
    wire \U409_CIA.g0Z0Z_10 ;
    wire \U409_CIA.g0Z0Z_2_cascade_ ;
    wire A_c_29;
    wire A_c_28;
    wire A_c_27;
    wire A_c_30;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_3 ;
    wire TT_c_1;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire PORTSIZE_0_i;
    wire bfn_8_8_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_8_9_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire bfn_8_13_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_nREGSPACE_i;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_nCIACS1_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_nCIACS0_i;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire U409_ADDRESS_DECODE_un1_nRAMSPACE_i;
    wire CLK28_IN_c_g;
    wire CIA_ENABLEm;
    wire A_c_22;
    wire A_c_23;
    wire A_c_21;
    wire AUTOVECTORm;
    wire ROMENm_i;
    wire \U409_ADDRESS_DECODE.LOWROMZ0 ;
    wire \U409_ADDRESS_DECODE.HIROMZ0 ;
    wire ROMENm;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ;
    wire \U409_TRANSFER_ACK.m9_am_cascade_ ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ;
    wire \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0 ;
    wire OVL_c;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.N_107 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_107_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_bm ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire CLKCIA_c;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire CONSTANT_ONE_NET;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_12_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_12_7_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire CLK6_c_g;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire RESETn_c_i;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire TACK_EN_i;
    wire N_373_i;
    wire RESETn_c;
    wire nBUFEN_c;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__5110),
            .RESETB(N__4891),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6282),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6284),
            .DIN(N__6283),
            .DOUT(N__6282),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6284),
            .PADOUT(N__6283),
            .PADIN(N__6282),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6272),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6274),
            .DIN(N__6273),
            .DOUT(N__6272),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6274),
            .PADOUT(N__6273),
            .PADIN(N__6272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__6263),
            .DIN(N__6262),
            .DOUT(N__6261),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__6263),
            .PADOUT(N__6262),
            .PADIN(N__6261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6254),
            .DIN(N__6253),
            .DOUT(N__6252),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6254),
            .PADOUT(N__6253),
            .PADIN(N__6252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4948),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6245),
            .DIN(N__6244),
            .DOUT(N__6243),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6245),
            .PADOUT(N__6244),
            .PADIN(N__6243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6236),
            .DIN(N__6235),
            .DOUT(N__6234),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6236),
            .PADOUT(N__6235),
            .PADIN(N__6234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS0_obuf_iopad (
            .OE(N__6227),
            .DIN(N__6226),
            .DOUT(N__6225),
            .PACKAGEPIN(nCIACS0));
    defparam nCIACS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS0_obuf_preio (
            .PADOEN(N__6227),
            .PADOUT(N__6226),
            .PADIN(N__6225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS1_obuf_iopad (
            .OE(N__6218),
            .DIN(N__6217),
            .DOUT(N__6216),
            .PACKAGEPIN(nCIACS1));
    defparam nCIACS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS1_obuf_preio (
            .PADOEN(N__6218),
            .PADOUT(N__6217),
            .PADIN(N__6216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3109),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6209),
            .DIN(N__6208),
            .DOUT(N__6207),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6209),
            .PADOUT(N__6208),
            .PADIN(N__6207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6200),
            .DIN(N__6199),
            .DOUT(N__6198),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6200),
            .PADOUT(N__6199),
            .PADIN(N__6198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6191),
            .DIN(N__6190),
            .DOUT(N__6189),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6191),
            .PADOUT(N__6190),
            .PADIN(N__6189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__6182),
            .DIN(N__6181),
            .DOUT(N__6180),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__6182),
            .PADOUT(N__6181),
            .PADIN(N__6180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5878),
            .DIN0(TACKn_in),
            .DOUT0(N__5515),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6173),
            .DIN(N__6172),
            .DOUT(N__6171),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6173),
            .PADOUT(N__6172),
            .PADIN(N__6171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__6164),
            .DIN(N__6163),
            .DOUT(N__6162),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__6164),
            .PADOUT(N__6163),
            .PADIN(N__6162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6155),
            .DIN(N__6154),
            .DOUT(N__6153),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6155),
            .PADOUT(N__6154),
            .PADIN(N__6153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__6146),
            .DIN(N__6145),
            .DOUT(N__6144),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__6146),
            .PADOUT(N__6145),
            .PADIN(N__6144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nRAMSPACE_obuf_iopad (
            .OE(N__6137),
            .DIN(N__6136),
            .DOUT(N__6135),
            .PACKAGEPIN(nRAMSPACE));
    defparam nRAMSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nRAMSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nRAMSPACE_obuf_preio (
            .PADOEN(N__6137),
            .PADOUT(N__6136),
            .PADIN(N__6135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nROMEN_obuf_iopad (
            .OE(N__6128),
            .DIN(N__6127),
            .DOUT(N__6126),
            .PACKAGEPIN(nROMEN));
    defparam nROMEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nROMEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nROMEN_obuf_preio (
            .PADOEN(N__6128),
            .PADOUT(N__6127),
            .PADIN(N__6126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6119),
            .DIN(N__6118),
            .DOUT(N__6117),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6119),
            .PADOUT(N__6118),
            .PADIN(N__6117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6110),
            .DIN(N__6109),
            .DOUT(N__6108),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6110),
            .PADOUT(N__6109),
            .PADIN(N__6108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nBUFEN_obuf_iopad (
            .OE(N__6101),
            .DIN(N__6100),
            .DOUT(N__6099),
            .PACKAGEPIN(nBUFEN));
    defparam nBUFEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nBUFEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nBUFEN_obuf_preio (
            .PADOEN(N__6101),
            .PADOUT(N__6100),
            .PADIN(N__6099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5713),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6092),
            .DIN(N__6091),
            .DOUT(N__6090),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6092),
            .PADOUT(N__6091),
            .PADIN(N__6090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6083),
            .DIN(N__6082),
            .DOUT(N__6081),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6083),
            .PADOUT(N__6082),
            .PADIN(N__6081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6074),
            .DIN(N__6073),
            .DOUT(N__6072),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6074),
            .PADOUT(N__6073),
            .PADIN(N__6072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__6065),
            .DIN(N__6064),
            .DOUT(N__6063),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__6065),
            .PADOUT(N__6064),
            .PADIN(N__6063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6056),
            .DIN(N__6055),
            .DOUT(N__6054),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6056),
            .PADOUT(N__6055),
            .PADIN(N__6054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6047),
            .DIN(N__6046),
            .DOUT(N__6045),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6047),
            .PADOUT(N__6046),
            .PADIN(N__6045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6038),
            .DIN(N__6037),
            .DOUT(N__6036),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6038),
            .PADOUT(N__6037),
            .PADIN(N__6036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nREGSPACE_obuf_iopad (
            .OE(N__6029),
            .DIN(N__6028),
            .DOUT(N__6027),
            .PACKAGEPIN(nREGSPACE));
    defparam nREGSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nREGSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nREGSPACE_obuf_preio (
            .PADOEN(N__6029),
            .PADOUT(N__6028),
            .PADIN(N__6027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__6020),
            .DIN(N__6019),
            .DOUT(N__6018),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__6020),
            .PADOUT(N__6019),
            .PADIN(N__6018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3448),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6011),
            .DIN(N__6010),
            .DOUT(N__6009),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6011),
            .PADOUT(N__6010),
            .PADIN(N__6009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6002),
            .DIN(N__6001),
            .DOUT(N__6000),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6002),
            .PADOUT(N__6001),
            .PADIN(N__6000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__5993),
            .DIN(N__5992),
            .DOUT(N__5991),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__5993),
            .PADOUT(N__5992),
            .PADIN(N__5991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__5984),
            .DIN(N__5983),
            .DOUT(N__5982),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__5984),
            .PADOUT(N__5983),
            .PADIN(N__5982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__5975),
            .DIN(N__5974),
            .DOUT(N__5973),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__5975),
            .PADOUT(N__5974),
            .PADIN(N__5973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__5966),
            .DIN(N__5965),
            .DOUT(N__5964),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__5966),
            .PADOUT(N__5965),
            .PADIN(N__5964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4576),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__5957),
            .DIN(N__5956),
            .DOUT(N__5955),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__5957),
            .PADOUT(N__5956),
            .PADIN(N__5955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1376 (
            .O(N__5938),
            .I(N__5929));
    InMux I__1375 (
            .O(N__5937),
            .I(N__5929));
    InMux I__1374 (
            .O(N__5936),
            .I(N__5929));
    LocalMux I__1373 (
            .O(N__5929),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1372 (
            .O(N__5926),
            .I(N__5917));
    InMux I__1371 (
            .O(N__5925),
            .I(N__5917));
    InMux I__1370 (
            .O(N__5924),
            .I(N__5917));
    LocalMux I__1369 (
            .O(N__5917),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1368 (
            .O(N__5914),
            .I(N__5910));
    InMux I__1367 (
            .O(N__5913),
            .I(N__5907));
    LocalMux I__1366 (
            .O(N__5910),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__1365 (
            .O(N__5907),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__1364 (
            .O(N__5902),
            .I(N__5899));
    LocalMux I__1363 (
            .O(N__5899),
            .I(N__5896));
    Span4Mux_h I__1362 (
            .O(N__5896),
            .I(N__5893));
    Odrv4 I__1361 (
            .O(N__5893),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    InMux I__1360 (
            .O(N__5890),
            .I(N__5887));
    LocalMux I__1359 (
            .O(N__5887),
            .I(N__5884));
    Span4Mux_v I__1358 (
            .O(N__5884),
            .I(N__5881));
    Odrv4 I__1357 (
            .O(N__5881),
            .I(TACK_EN_i));
    IoInMux I__1356 (
            .O(N__5878),
            .I(N__5875));
    LocalMux I__1355 (
            .O(N__5875),
            .I(N__5872));
    Span4Mux_s0_v I__1354 (
            .O(N__5872),
            .I(N__5869));
    Sp12to4 I__1353 (
            .O(N__5869),
            .I(N__5866));
    Span12Mux_h I__1352 (
            .O(N__5866),
            .I(N__5863));
    Odrv12 I__1351 (
            .O(N__5863),
            .I(N_373_i));
    InMux I__1350 (
            .O(N__5860),
            .I(N__5853));
    InMux I__1349 (
            .O(N__5859),
            .I(N__5848));
    InMux I__1348 (
            .O(N__5858),
            .I(N__5848));
    InMux I__1347 (
            .O(N__5857),
            .I(N__5845));
    InMux I__1346 (
            .O(N__5856),
            .I(N__5842));
    LocalMux I__1345 (
            .O(N__5853),
            .I(N__5835));
    LocalMux I__1344 (
            .O(N__5848),
            .I(N__5832));
    LocalMux I__1343 (
            .O(N__5845),
            .I(N__5829));
    LocalMux I__1342 (
            .O(N__5842),
            .I(N__5826));
    InMux I__1341 (
            .O(N__5841),
            .I(N__5821));
    InMux I__1340 (
            .O(N__5840),
            .I(N__5821));
    CascadeMux I__1339 (
            .O(N__5839),
            .I(N__5818));
    InMux I__1338 (
            .O(N__5838),
            .I(N__5814));
    Span4Mux_v I__1337 (
            .O(N__5835),
            .I(N__5811));
    Span4Mux_v I__1336 (
            .O(N__5832),
            .I(N__5808));
    Span4Mux_v I__1335 (
            .O(N__5829),
            .I(N__5805));
    Span4Mux_v I__1334 (
            .O(N__5826),
            .I(N__5799));
    LocalMux I__1333 (
            .O(N__5821),
            .I(N__5799));
    InMux I__1332 (
            .O(N__5818),
            .I(N__5794));
    InMux I__1331 (
            .O(N__5817),
            .I(N__5794));
    LocalMux I__1330 (
            .O(N__5814),
            .I(N__5789));
    Sp12to4 I__1329 (
            .O(N__5811),
            .I(N__5785));
    Span4Mux_h I__1328 (
            .O(N__5808),
            .I(N__5782));
    Sp12to4 I__1327 (
            .O(N__5805),
            .I(N__5779));
    InMux I__1326 (
            .O(N__5804),
            .I(N__5776));
    Span4Mux_h I__1325 (
            .O(N__5799),
            .I(N__5771));
    LocalMux I__1324 (
            .O(N__5794),
            .I(N__5771));
    InMux I__1323 (
            .O(N__5793),
            .I(N__5766));
    InMux I__1322 (
            .O(N__5792),
            .I(N__5766));
    Span4Mux_v I__1321 (
            .O(N__5789),
            .I(N__5763));
    InMux I__1320 (
            .O(N__5788),
            .I(N__5760));
    Span12Mux_h I__1319 (
            .O(N__5785),
            .I(N__5757));
    Sp12to4 I__1318 (
            .O(N__5782),
            .I(N__5754));
    Span12Mux_h I__1317 (
            .O(N__5779),
            .I(N__5745));
    LocalMux I__1316 (
            .O(N__5776),
            .I(N__5745));
    Sp12to4 I__1315 (
            .O(N__5771),
            .I(N__5745));
    LocalMux I__1314 (
            .O(N__5766),
            .I(N__5745));
    Sp12to4 I__1313 (
            .O(N__5763),
            .I(N__5740));
    LocalMux I__1312 (
            .O(N__5760),
            .I(N__5740));
    Span12Mux_v I__1311 (
            .O(N__5757),
            .I(N__5737));
    Span12Mux_h I__1310 (
            .O(N__5754),
            .I(N__5734));
    Span12Mux_v I__1309 (
            .O(N__5745),
            .I(N__5731));
    Span12Mux_h I__1308 (
            .O(N__5740),
            .I(N__5728));
    Span12Mux_h I__1307 (
            .O(N__5737),
            .I(N__5723));
    Span12Mux_v I__1306 (
            .O(N__5734),
            .I(N__5723));
    Span12Mux_h I__1305 (
            .O(N__5731),
            .I(N__5718));
    Span12Mux_v I__1304 (
            .O(N__5728),
            .I(N__5718));
    Odrv12 I__1303 (
            .O(N__5723),
            .I(RESETn_c));
    Odrv12 I__1302 (
            .O(N__5718),
            .I(RESETn_c));
    IoInMux I__1301 (
            .O(N__5713),
            .I(N__5710));
    LocalMux I__1300 (
            .O(N__5710),
            .I(N__5707));
    Span12Mux_s10_v I__1299 (
            .O(N__5707),
            .I(N__5703));
    InMux I__1298 (
            .O(N__5706),
            .I(N__5700));
    Span12Mux_h I__1297 (
            .O(N__5703),
            .I(N__5697));
    LocalMux I__1296 (
            .O(N__5700),
            .I(N__5694));
    Odrv12 I__1295 (
            .O(N__5697),
            .I(nBUFEN_c));
    Odrv12 I__1294 (
            .O(N__5694),
            .I(nBUFEN_c));
    InMux I__1293 (
            .O(N__5689),
            .I(N__5686));
    LocalMux I__1292 (
            .O(N__5686),
            .I(N__5683));
    Span4Mux_h I__1291 (
            .O(N__5683),
            .I(N__5680));
    Span4Mux_h I__1290 (
            .O(N__5680),
            .I(N__5677));
    Sp12to4 I__1289 (
            .O(N__5677),
            .I(N__5674));
    Span12Mux_v I__1288 (
            .O(N__5674),
            .I(N__5671));
    Odrv12 I__1287 (
            .O(N__5671),
            .I(TACKn_in));
    SRMux I__1286 (
            .O(N__5668),
            .I(N__5665));
    LocalMux I__1285 (
            .O(N__5665),
            .I(N__5661));
    SRMux I__1284 (
            .O(N__5664),
            .I(N__5658));
    Span4Mux_v I__1283 (
            .O(N__5661),
            .I(N__5655));
    LocalMux I__1282 (
            .O(N__5658),
            .I(N__5652));
    Sp12to4 I__1281 (
            .O(N__5655),
            .I(N__5647));
    Span12Mux_v I__1280 (
            .O(N__5652),
            .I(N__5647));
    Odrv12 I__1279 (
            .O(N__5647),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1278 (
            .O(N__5644),
            .I(N__5641));
    LocalMux I__1277 (
            .O(N__5641),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ));
    CascadeMux I__1276 (
            .O(N__5638),
            .I(N__5634));
    InMux I__1275 (
            .O(N__5637),
            .I(N__5626));
    InMux I__1274 (
            .O(N__5634),
            .I(N__5626));
    InMux I__1273 (
            .O(N__5633),
            .I(N__5626));
    LocalMux I__1272 (
            .O(N__5626),
            .I(N__5623));
    Span4Mux_v I__1271 (
            .O(N__5623),
            .I(N__5620));
    Span4Mux_v I__1270 (
            .O(N__5620),
            .I(N__5617));
    Odrv4 I__1269 (
            .O(N__5617),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    InMux I__1268 (
            .O(N__5614),
            .I(N__5607));
    InMux I__1267 (
            .O(N__5613),
            .I(N__5607));
    InMux I__1266 (
            .O(N__5612),
            .I(N__5604));
    LocalMux I__1265 (
            .O(N__5607),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1264 (
            .O(N__5604),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1263 (
            .O(N__5599),
            .I(N__5589));
    InMux I__1262 (
            .O(N__5598),
            .I(N__5589));
    InMux I__1261 (
            .O(N__5597),
            .I(N__5589));
    InMux I__1260 (
            .O(N__5596),
            .I(N__5586));
    LocalMux I__1259 (
            .O(N__5589),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1258 (
            .O(N__5586),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1257 (
            .O(N__5581),
            .I(N__5576));
    InMux I__1256 (
            .O(N__5580),
            .I(N__5570));
    InMux I__1255 (
            .O(N__5579),
            .I(N__5570));
    InMux I__1254 (
            .O(N__5576),
            .I(N__5565));
    InMux I__1253 (
            .O(N__5575),
            .I(N__5565));
    LocalMux I__1252 (
            .O(N__5570),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1251 (
            .O(N__5565),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    SRMux I__1250 (
            .O(N__5560),
            .I(N__5555));
    SRMux I__1249 (
            .O(N__5559),
            .I(N__5552));
    SRMux I__1248 (
            .O(N__5558),
            .I(N__5549));
    LocalMux I__1247 (
            .O(N__5555),
            .I(N__5545));
    LocalMux I__1246 (
            .O(N__5552),
            .I(N__5542));
    LocalMux I__1245 (
            .O(N__5549),
            .I(N__5539));
    SRMux I__1244 (
            .O(N__5548),
            .I(N__5536));
    Span4Mux_v I__1243 (
            .O(N__5545),
            .I(N__5533));
    Span4Mux_v I__1242 (
            .O(N__5542),
            .I(N__5530));
    Span4Mux_h I__1241 (
            .O(N__5539),
            .I(N__5527));
    LocalMux I__1240 (
            .O(N__5536),
            .I(N__5524));
    Odrv4 I__1239 (
            .O(N__5533),
            .I(RESETn_c_i));
    Odrv4 I__1238 (
            .O(N__5530),
            .I(RESETn_c_i));
    Odrv4 I__1237 (
            .O(N__5527),
            .I(RESETn_c_i));
    Odrv12 I__1236 (
            .O(N__5524),
            .I(RESETn_c_i));
    IoInMux I__1235 (
            .O(N__5515),
            .I(N__5512));
    LocalMux I__1234 (
            .O(N__5512),
            .I(N__5509));
    Span12Mux_s7_v I__1233 (
            .O(N__5509),
            .I(N__5506));
    Span12Mux_h I__1232 (
            .O(N__5506),
            .I(N__5502));
    InMux I__1231 (
            .O(N__5505),
            .I(N__5499));
    Odrv12 I__1230 (
            .O(N__5502),
            .I(TACK_OUTn));
    LocalMux I__1229 (
            .O(N__5499),
            .I(TACK_OUTn));
    CascadeMux I__1228 (
            .O(N__5494),
            .I(N__5491));
    InMux I__1227 (
            .O(N__5491),
            .I(N__5486));
    InMux I__1226 (
            .O(N__5490),
            .I(N__5483));
    InMux I__1225 (
            .O(N__5489),
            .I(N__5480));
    LocalMux I__1224 (
            .O(N__5486),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1223 (
            .O(N__5483),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1222 (
            .O(N__5480),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1221 (
            .O(N__5473),
            .I(N__5469));
    InMux I__1220 (
            .O(N__5472),
            .I(N__5466));
    LocalMux I__1219 (
            .O(N__5469),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1218 (
            .O(N__5466),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__1217 (
            .O(N__5461),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ));
    InMux I__1216 (
            .O(N__5458),
            .I(N__5454));
    InMux I__1215 (
            .O(N__5457),
            .I(N__5451));
    LocalMux I__1214 (
            .O(N__5454),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1213 (
            .O(N__5451),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__1212 (
            .O(N__5446),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    InMux I__1211 (
            .O(N__5443),
            .I(N__5439));
    InMux I__1210 (
            .O(N__5442),
            .I(N__5436));
    LocalMux I__1209 (
            .O(N__5439),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1208 (
            .O(N__5436),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__1207 (
            .O(N__5431),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1206 (
            .O(N__5428),
            .I(N__5424));
    InMux I__1205 (
            .O(N__5427),
            .I(N__5421));
    LocalMux I__1204 (
            .O(N__5424),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1203 (
            .O(N__5421),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__1202 (
            .O(N__5416),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1201 (
            .O(N__5413),
            .I(N__5409));
    InMux I__1200 (
            .O(N__5412),
            .I(N__5406));
    LocalMux I__1199 (
            .O(N__5409),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1198 (
            .O(N__5406),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1197 (
            .O(N__5401),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    CascadeMux I__1196 (
            .O(N__5398),
            .I(N__5395));
    InMux I__1195 (
            .O(N__5395),
            .I(N__5391));
    InMux I__1194 (
            .O(N__5394),
            .I(N__5388));
    LocalMux I__1193 (
            .O(N__5391),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1192 (
            .O(N__5388),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1191 (
            .O(N__5383),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1190 (
            .O(N__5380),
            .I(N__5376));
    InMux I__1189 (
            .O(N__5379),
            .I(N__5373));
    LocalMux I__1188 (
            .O(N__5376),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__1187 (
            .O(N__5373),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__1186 (
            .O(N__5368),
            .I(N__5365));
    LocalMux I__1185 (
            .O(N__5365),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__1184 (
            .O(N__5362),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1183 (
            .O(N__5359),
            .I(N__5355));
    InMux I__1182 (
            .O(N__5358),
            .I(N__5352));
    LocalMux I__1181 (
            .O(N__5355),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1180 (
            .O(N__5352),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1179 (
            .O(N__5347),
            .I(N__5344));
    LocalMux I__1178 (
            .O(N__5344),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1177 (
            .O(N__5341),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1176 (
            .O(N__5338),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1175 (
            .O(N__5335),
            .I(N__5331));
    InMux I__1174 (
            .O(N__5334),
            .I(N__5328));
    LocalMux I__1173 (
            .O(N__5331),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1172 (
            .O(N__5328),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    ClkMux I__1171 (
            .O(N__5323),
            .I(N__5299));
    ClkMux I__1170 (
            .O(N__5322),
            .I(N__5299));
    ClkMux I__1169 (
            .O(N__5321),
            .I(N__5299));
    ClkMux I__1168 (
            .O(N__5320),
            .I(N__5299));
    ClkMux I__1167 (
            .O(N__5319),
            .I(N__5299));
    ClkMux I__1166 (
            .O(N__5318),
            .I(N__5299));
    ClkMux I__1165 (
            .O(N__5317),
            .I(N__5299));
    ClkMux I__1164 (
            .O(N__5316),
            .I(N__5299));
    GlobalMux I__1163 (
            .O(N__5299),
            .I(N__5296));
    gio2CtrlBuf I__1162 (
            .O(N__5296),
            .I(CLK6_c_g));
    CascadeMux I__1161 (
            .O(N__5293),
            .I(N__5290));
    InMux I__1160 (
            .O(N__5290),
            .I(N__5286));
    InMux I__1159 (
            .O(N__5289),
            .I(N__5283));
    LocalMux I__1158 (
            .O(N__5286),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1157 (
            .O(N__5283),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__1156 (
            .O(N__5278),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1155 (
            .O(N__5275),
            .I(N__5272));
    LocalMux I__1154 (
            .O(N__5272),
            .I(N__5268));
    InMux I__1153 (
            .O(N__5271),
            .I(N__5265));
    Odrv4 I__1152 (
            .O(N__5268),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1151 (
            .O(N__5265),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__1150 (
            .O(N__5260),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1149 (
            .O(N__5257),
            .I(N__5253));
    InMux I__1148 (
            .O(N__5256),
            .I(N__5250));
    LocalMux I__1147 (
            .O(N__5253),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__1146 (
            .O(N__5250),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__1145 (
            .O(N__5245),
            .I(N__5242));
    LocalMux I__1144 (
            .O(N__5242),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1143 (
            .O(N__5239),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1142 (
            .O(N__5236),
            .I(N__5232));
    InMux I__1141 (
            .O(N__5235),
            .I(N__5229));
    LocalMux I__1140 (
            .O(N__5232),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1139 (
            .O(N__5229),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1138 (
            .O(N__5224),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1137 (
            .O(N__5221),
            .I(N__5217));
    InMux I__1136 (
            .O(N__5220),
            .I(N__5214));
    LocalMux I__1135 (
            .O(N__5217),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__1134 (
            .O(N__5214),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__1133 (
            .O(N__5209),
            .I(N__5206));
    LocalMux I__1132 (
            .O(N__5206),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1131 (
            .O(N__5203),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__1130 (
            .O(N__5200),
            .I(N__5196));
    InMux I__1129 (
            .O(N__5199),
            .I(N__5193));
    LocalMux I__1128 (
            .O(N__5196),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1127 (
            .O(N__5193),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__1126 (
            .O(N__5188),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__1125 (
            .O(N__5185),
            .I(N__5181));
    InMux I__1124 (
            .O(N__5184),
            .I(N__5178));
    LocalMux I__1123 (
            .O(N__5181),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__1122 (
            .O(N__5178),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__1121 (
            .O(N__5173),
            .I(N__5170));
    InMux I__1120 (
            .O(N__5170),
            .I(N__5167));
    LocalMux I__1119 (
            .O(N__5167),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1118 (
            .O(N__5164),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    CascadeMux I__1117 (
            .O(N__5161),
            .I(N__5158));
    InMux I__1116 (
            .O(N__5158),
            .I(N__5154));
    InMux I__1115 (
            .O(N__5157),
            .I(N__5151));
    LocalMux I__1114 (
            .O(N__5154),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__1113 (
            .O(N__5151),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__1112 (
            .O(N__5146),
            .I(N__5143));
    InMux I__1111 (
            .O(N__5143),
            .I(N__5140));
    LocalMux I__1110 (
            .O(N__5140),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__1109 (
            .O(N__5137),
            .I(bfn_12_7_0_));
    InMux I__1108 (
            .O(N__5134),
            .I(N__5127));
    InMux I__1107 (
            .O(N__5133),
            .I(N__5120));
    InMux I__1106 (
            .O(N__5132),
            .I(N__5120));
    InMux I__1105 (
            .O(N__5131),
            .I(N__5120));
    InMux I__1104 (
            .O(N__5130),
            .I(N__5117));
    LocalMux I__1103 (
            .O(N__5127),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1102 (
            .O(N__5120),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1101 (
            .O(N__5117),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    IoInMux I__1100 (
            .O(N__5110),
            .I(N__5107));
    LocalMux I__1099 (
            .O(N__5107),
            .I(N__5104));
    IoSpan4Mux I__1098 (
            .O(N__5104),
            .I(N__5097));
    InMux I__1097 (
            .O(N__5103),
            .I(N__5094));
    InMux I__1096 (
            .O(N__5102),
            .I(N__5091));
    CascadeMux I__1095 (
            .O(N__5101),
            .I(N__5088));
    InMux I__1094 (
            .O(N__5100),
            .I(N__5085));
    Span4Mux_s0_v I__1093 (
            .O(N__5097),
            .I(N__5082));
    LocalMux I__1092 (
            .O(N__5094),
            .I(N__5077));
    LocalMux I__1091 (
            .O(N__5091),
            .I(N__5077));
    InMux I__1090 (
            .O(N__5088),
            .I(N__5074));
    LocalMux I__1089 (
            .O(N__5085),
            .I(N__5071));
    Sp12to4 I__1088 (
            .O(N__5082),
            .I(N__5068));
    Span4Mux_h I__1087 (
            .O(N__5077),
            .I(N__5063));
    LocalMux I__1086 (
            .O(N__5074),
            .I(N__5063));
    Span4Mux_h I__1085 (
            .O(N__5071),
            .I(N__5060));
    Span12Mux_v I__1084 (
            .O(N__5068),
            .I(N__5055));
    Sp12to4 I__1083 (
            .O(N__5063),
            .I(N__5055));
    Sp12to4 I__1082 (
            .O(N__5060),
            .I(N__5052));
    Span12Mux_v I__1081 (
            .O(N__5055),
            .I(N__5049));
    Odrv12 I__1080 (
            .O(N__5052),
            .I(CLK40_IN_c));
    Odrv12 I__1079 (
            .O(N__5049),
            .I(CLK40_IN_c));
    CascadeMux I__1078 (
            .O(N__5044),
            .I(N__5041));
    InMux I__1077 (
            .O(N__5041),
            .I(N__5038));
    LocalMux I__1076 (
            .O(N__5038),
            .I(\U409_TRANSFER_ACK.N_107 ));
    CascadeMux I__1075 (
            .O(N__5035),
            .I(N__5029));
    InMux I__1074 (
            .O(N__5034),
            .I(N__5026));
    InMux I__1073 (
            .O(N__5033),
            .I(N__5023));
    InMux I__1072 (
            .O(N__5032),
            .I(N__5018));
    InMux I__1071 (
            .O(N__5029),
            .I(N__5018));
    LocalMux I__1070 (
            .O(N__5026),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1069 (
            .O(N__5023),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1068 (
            .O(N__5018),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__1067 (
            .O(N__5011),
            .I(\U409_TRANSFER_ACK.N_107_cascade_ ));
    InMux I__1066 (
            .O(N__5008),
            .I(N__5005));
    LocalMux I__1065 (
            .O(N__5005),
            .I(\U409_TRANSFER_ACK.m9_bm ));
    InMux I__1064 (
            .O(N__5002),
            .I(N__4996));
    InMux I__1063 (
            .O(N__5001),
            .I(N__4996));
    LocalMux I__1062 (
            .O(N__4996),
            .I(\U409_TRANSFER_ACK.N_4 ));
    InMux I__1061 (
            .O(N__4993),
            .I(N__4987));
    InMux I__1060 (
            .O(N__4992),
            .I(N__4984));
    InMux I__1059 (
            .O(N__4991),
            .I(N__4981));
    InMux I__1058 (
            .O(N__4990),
            .I(N__4978));
    LocalMux I__1057 (
            .O(N__4987),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1056 (
            .O(N__4984),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1055 (
            .O(N__4981),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1054 (
            .O(N__4978),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__1053 (
            .O(N__4969),
            .I(N__4966));
    InMux I__1052 (
            .O(N__4966),
            .I(N__4960));
    InMux I__1051 (
            .O(N__4965),
            .I(N__4960));
    LocalMux I__1050 (
            .O(N__4960),
            .I(N__4956));
    InMux I__1049 (
            .O(N__4959),
            .I(N__4953));
    Odrv4 I__1048 (
            .O(N__4956),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__1047 (
            .O(N__4953),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    IoInMux I__1046 (
            .O(N__4948),
            .I(N__4945));
    LocalMux I__1045 (
            .O(N__4945),
            .I(N__4942));
    IoSpan4Mux I__1044 (
            .O(N__4942),
            .I(N__4939));
    Span4Mux_s1_v I__1043 (
            .O(N__4939),
            .I(N__4936));
    Sp12to4 I__1042 (
            .O(N__4936),
            .I(N__4932));
    InMux I__1041 (
            .O(N__4935),
            .I(N__4929));
    Span12Mux_v I__1040 (
            .O(N__4932),
            .I(N__4923));
    LocalMux I__1039 (
            .O(N__4929),
            .I(N__4923));
    InMux I__1038 (
            .O(N__4928),
            .I(N__4920));
    Odrv12 I__1037 (
            .O(N__4923),
            .I(CLKCIA_c));
    LocalMux I__1036 (
            .O(N__4920),
            .I(CLKCIA_c));
    InMux I__1035 (
            .O(N__4915),
            .I(N__4910));
    InMux I__1034 (
            .O(N__4914),
            .I(N__4905));
    InMux I__1033 (
            .O(N__4913),
            .I(N__4905));
    LocalMux I__1032 (
            .O(N__4910),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1031 (
            .O(N__4905),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1030 (
            .O(N__4900),
            .I(N__4894));
    InMux I__1029 (
            .O(N__4899),
            .I(N__4894));
    LocalMux I__1028 (
            .O(N__4894),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    IoInMux I__1027 (
            .O(N__4891),
            .I(N__4888));
    LocalMux I__1026 (
            .O(N__4888),
            .I(N__4885));
    Span4Mux_s2_v I__1025 (
            .O(N__4885),
            .I(N__4882));
    Span4Mux_v I__1024 (
            .O(N__4882),
            .I(N__4879));
    Odrv4 I__1023 (
            .O(N__4879),
            .I(CONSTANT_ONE_NET));
    InMux I__1022 (
            .O(N__4876),
            .I(N__4869));
    InMux I__1021 (
            .O(N__4875),
            .I(N__4869));
    InMux I__1020 (
            .O(N__4874),
            .I(N__4866));
    LocalMux I__1019 (
            .O(N__4869),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1018 (
            .O(N__4866),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__1017 (
            .O(N__4861),
            .I(N__4855));
    InMux I__1016 (
            .O(N__4860),
            .I(N__4848));
    InMux I__1015 (
            .O(N__4859),
            .I(N__4848));
    InMux I__1014 (
            .O(N__4858),
            .I(N__4848));
    InMux I__1013 (
            .O(N__4855),
            .I(N__4845));
    LocalMux I__1012 (
            .O(N__4848),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1011 (
            .O(N__4845),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__1010 (
            .O(N__4840),
            .I(N__4835));
    InMux I__1009 (
            .O(N__4839),
            .I(N__4832));
    InMux I__1008 (
            .O(N__4838),
            .I(N__4829));
    LocalMux I__1007 (
            .O(N__4835),
            .I(N__4826));
    LocalMux I__1006 (
            .O(N__4832),
            .I(N__4821));
    LocalMux I__1005 (
            .O(N__4829),
            .I(N__4821));
    Span4Mux_v I__1004 (
            .O(N__4826),
            .I(N__4818));
    Span12Mux_h I__1003 (
            .O(N__4821),
            .I(N__4815));
    Sp12to4 I__1002 (
            .O(N__4818),
            .I(N__4812));
    Span12Mux_v I__1001 (
            .O(N__4815),
            .I(N__4809));
    Span12Mux_h I__1000 (
            .O(N__4812),
            .I(N__4806));
    Odrv12 I__999 (
            .O(N__4809),
            .I(TSn_c));
    Odrv12 I__998 (
            .O(N__4806),
            .I(TSn_c));
    InMux I__997 (
            .O(N__4801),
            .I(N__4795));
    InMux I__996 (
            .O(N__4800),
            .I(N__4790));
    InMux I__995 (
            .O(N__4799),
            .I(N__4790));
    InMux I__994 (
            .O(N__4798),
            .I(N__4787));
    LocalMux I__993 (
            .O(N__4795),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__992 (
            .O(N__4790),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__991 (
            .O(N__4787),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__990 (
            .O(N__4780),
            .I(N__4775));
    CascadeMux I__989 (
            .O(N__4779),
            .I(N__4769));
    CascadeMux I__988 (
            .O(N__4778),
            .I(N__4766));
    InMux I__987 (
            .O(N__4775),
            .I(N__4758));
    InMux I__986 (
            .O(N__4774),
            .I(N__4758));
    InMux I__985 (
            .O(N__4773),
            .I(N__4758));
    InMux I__984 (
            .O(N__4772),
            .I(N__4753));
    InMux I__983 (
            .O(N__4769),
            .I(N__4753));
    InMux I__982 (
            .O(N__4766),
            .I(N__4750));
    InMux I__981 (
            .O(N__4765),
            .I(N__4747));
    LocalMux I__980 (
            .O(N__4758),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__979 (
            .O(N__4753),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__978 (
            .O(N__4750),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__977 (
            .O(N__4747),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__976 (
            .O(N__4738),
            .I(N__4729));
    InMux I__975 (
            .O(N__4737),
            .I(N__4729));
    InMux I__974 (
            .O(N__4736),
            .I(N__4724));
    InMux I__973 (
            .O(N__4735),
            .I(N__4724));
    InMux I__972 (
            .O(N__4734),
            .I(N__4721));
    LocalMux I__971 (
            .O(N__4729),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__970 (
            .O(N__4724),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__969 (
            .O(N__4721),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__968 (
            .O(N__4714),
            .I(N__4711));
    LocalMux I__967 (
            .O(N__4711),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__966 (
            .O(N__4708),
            .I(N__4701));
    InMux I__965 (
            .O(N__4707),
            .I(N__4701));
    InMux I__964 (
            .O(N__4706),
            .I(N__4698));
    LocalMux I__963 (
            .O(N__4701),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__962 (
            .O(N__4698),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__961 (
            .O(N__4693),
            .I(N__4690));
    LocalMux I__960 (
            .O(N__4690),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ));
    InMux I__959 (
            .O(N__4687),
            .I(N__4681));
    InMux I__958 (
            .O(N__4686),
            .I(N__4678));
    InMux I__957 (
            .O(N__4685),
            .I(N__4673));
    InMux I__956 (
            .O(N__4684),
            .I(N__4673));
    LocalMux I__955 (
            .O(N__4681),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__954 (
            .O(N__4678),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__953 (
            .O(N__4673),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__952 (
            .O(N__4666),
            .I(N__4657));
    InMux I__951 (
            .O(N__4665),
            .I(N__4657));
    InMux I__950 (
            .O(N__4664),
            .I(N__4654));
    InMux I__949 (
            .O(N__4663),
            .I(N__4651));
    InMux I__948 (
            .O(N__4662),
            .I(N__4648));
    LocalMux I__947 (
            .O(N__4657),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__946 (
            .O(N__4654),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__945 (
            .O(N__4651),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__944 (
            .O(N__4648),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__943 (
            .O(N__4639),
            .I(N__4636));
    InMux I__942 (
            .O(N__4636),
            .I(N__4630));
    InMux I__941 (
            .O(N__4635),
            .I(N__4630));
    LocalMux I__940 (
            .O(N__4630),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    InMux I__939 (
            .O(N__4627),
            .I(N__4620));
    InMux I__938 (
            .O(N__4626),
            .I(N__4611));
    InMux I__937 (
            .O(N__4625),
            .I(N__4611));
    InMux I__936 (
            .O(N__4624),
            .I(N__4611));
    InMux I__935 (
            .O(N__4623),
            .I(N__4611));
    LocalMux I__934 (
            .O(N__4620),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__933 (
            .O(N__4611),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__932 (
            .O(N__4606),
            .I(N__4600));
    InMux I__931 (
            .O(N__4605),
            .I(N__4597));
    InMux I__930 (
            .O(N__4604),
            .I(N__4594));
    InMux I__929 (
            .O(N__4603),
            .I(N__4589));
    InMux I__928 (
            .O(N__4600),
            .I(N__4589));
    LocalMux I__927 (
            .O(N__4597),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__926 (
            .O(N__4594),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__925 (
            .O(N__4589),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    CascadeMux I__924 (
            .O(N__4582),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__923 (
            .O(N__4579),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    IoInMux I__922 (
            .O(N__4576),
            .I(N__4573));
    LocalMux I__921 (
            .O(N__4573),
            .I(N__4570));
    Span4Mux_s0_v I__920 (
            .O(N__4570),
            .I(N__4567));
    Sp12to4 I__919 (
            .O(N__4567),
            .I(N__4564));
    Span12Mux_h I__918 (
            .O(N__4564),
            .I(N__4561));
    Span12Mux_v I__917 (
            .O(N__4561),
            .I(N__4557));
    InMux I__916 (
            .O(N__4560),
            .I(N__4554));
    Odrv12 I__915 (
            .O(N__4557),
            .I(TICK60_c));
    LocalMux I__914 (
            .O(N__4554),
            .I(TICK60_c));
    InMux I__913 (
            .O(N__4549),
            .I(N__4536));
    InMux I__912 (
            .O(N__4548),
            .I(N__4536));
    InMux I__911 (
            .O(N__4547),
            .I(N__4536));
    InMux I__910 (
            .O(N__4546),
            .I(N__4527));
    InMux I__909 (
            .O(N__4545),
            .I(N__4527));
    InMux I__908 (
            .O(N__4544),
            .I(N__4527));
    InMux I__907 (
            .O(N__4543),
            .I(N__4527));
    LocalMux I__906 (
            .O(N__4536),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__905 (
            .O(N__4527),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__904 (
            .O(N__4522),
            .I(N__4518));
    InMux I__903 (
            .O(N__4521),
            .I(N__4510));
    InMux I__902 (
            .O(N__4518),
            .I(N__4507));
    InMux I__901 (
            .O(N__4517),
            .I(N__4496));
    InMux I__900 (
            .O(N__4516),
            .I(N__4496));
    InMux I__899 (
            .O(N__4515),
            .I(N__4496));
    InMux I__898 (
            .O(N__4514),
            .I(N__4496));
    InMux I__897 (
            .O(N__4513),
            .I(N__4496));
    LocalMux I__896 (
            .O(N__4510),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__895 (
            .O(N__4507),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__894 (
            .O(N__4496),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__893 (
            .O(N__4489),
            .I(N__4480));
    CascadeMux I__892 (
            .O(N__4488),
            .I(N__4477));
    InMux I__891 (
            .O(N__4487),
            .I(N__4472));
    InMux I__890 (
            .O(N__4486),
            .I(N__4472));
    InMux I__889 (
            .O(N__4485),
            .I(N__4461));
    InMux I__888 (
            .O(N__4484),
            .I(N__4461));
    InMux I__887 (
            .O(N__4483),
            .I(N__4461));
    InMux I__886 (
            .O(N__4480),
            .I(N__4461));
    InMux I__885 (
            .O(N__4477),
            .I(N__4461));
    LocalMux I__884 (
            .O(N__4472),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__883 (
            .O(N__4461),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__882 (
            .O(N__4456),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ));
    CascadeMux I__881 (
            .O(N__4453),
            .I(N__4450));
    InMux I__880 (
            .O(N__4450),
            .I(N__4444));
    InMux I__879 (
            .O(N__4449),
            .I(N__4444));
    LocalMux I__878 (
            .O(N__4444),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__877 (
            .O(N__4441),
            .I(N__4438));
    LocalMux I__876 (
            .O(N__4438),
            .I(N__4434));
    CascadeMux I__875 (
            .O(N__4437),
            .I(N__4431));
    Span4Mux_v I__874 (
            .O(N__4434),
            .I(N__4428));
    InMux I__873 (
            .O(N__4431),
            .I(N__4425));
    Odrv4 I__872 (
            .O(N__4428),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    LocalMux I__871 (
            .O(N__4425),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    InMux I__870 (
            .O(N__4420),
            .I(N__4416));
    InMux I__869 (
            .O(N__4419),
            .I(N__4413));
    LocalMux I__868 (
            .O(N__4416),
            .I(N__4410));
    LocalMux I__867 (
            .O(N__4413),
            .I(N__4407));
    Odrv4 I__866 (
            .O(N__4410),
            .I(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ));
    Odrv4 I__865 (
            .O(N__4407),
            .I(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ));
    CascadeMux I__864 (
            .O(N__4402),
            .I(N__4399));
    InMux I__863 (
            .O(N__4399),
            .I(N__4396));
    LocalMux I__862 (
            .O(N__4396),
            .I(N__4391));
    InMux I__861 (
            .O(N__4395),
            .I(N__4387));
    InMux I__860 (
            .O(N__4394),
            .I(N__4382));
    Span4Mux_v I__859 (
            .O(N__4391),
            .I(N__4379));
    InMux I__858 (
            .O(N__4390),
            .I(N__4376));
    LocalMux I__857 (
            .O(N__4387),
            .I(N__4373));
    InMux I__856 (
            .O(N__4386),
            .I(N__4368));
    InMux I__855 (
            .O(N__4385),
            .I(N__4368));
    LocalMux I__854 (
            .O(N__4382),
            .I(N__4364));
    Sp12to4 I__853 (
            .O(N__4379),
            .I(N__4359));
    LocalMux I__852 (
            .O(N__4376),
            .I(N__4359));
    Span4Mux_v I__851 (
            .O(N__4373),
            .I(N__4356));
    LocalMux I__850 (
            .O(N__4368),
            .I(N__4353));
    InMux I__849 (
            .O(N__4367),
            .I(N__4350));
    Span12Mux_v I__848 (
            .O(N__4364),
            .I(N__4347));
    Span12Mux_h I__847 (
            .O(N__4359),
            .I(N__4344));
    Span4Mux_h I__846 (
            .O(N__4356),
            .I(N__4341));
    Span4Mux_h I__845 (
            .O(N__4353),
            .I(N__4338));
    LocalMux I__844 (
            .O(N__4350),
            .I(N__4335));
    Odrv12 I__843 (
            .O(N__4347),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv12 I__842 (
            .O(N__4344),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__841 (
            .O(N__4341),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__840 (
            .O(N__4338),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__839 (
            .O(N__4335),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    InMux I__838 (
            .O(N__4324),
            .I(N__4321));
    LocalMux I__837 (
            .O(N__4321),
            .I(N__4318));
    Span4Mux_v I__836 (
            .O(N__4318),
            .I(N__4313));
    InMux I__835 (
            .O(N__4317),
            .I(N__4310));
    InMux I__834 (
            .O(N__4316),
            .I(N__4307));
    Sp12to4 I__833 (
            .O(N__4313),
            .I(N__4300));
    LocalMux I__832 (
            .O(N__4310),
            .I(N__4300));
    LocalMux I__831 (
            .O(N__4307),
            .I(N__4300));
    Span12Mux_h I__830 (
            .O(N__4300),
            .I(N__4297));
    Span12Mux_v I__829 (
            .O(N__4297),
            .I(N__4294));
    Odrv12 I__828 (
            .O(N__4294),
            .I(OVL_c));
    InMux I__827 (
            .O(N__4291),
            .I(N__4286));
    CascadeMux I__826 (
            .O(N__4290),
            .I(N__4282));
    CascadeMux I__825 (
            .O(N__4289),
            .I(N__4279));
    LocalMux I__824 (
            .O(N__4286),
            .I(N__4276));
    InMux I__823 (
            .O(N__4285),
            .I(N__4273));
    InMux I__822 (
            .O(N__4282),
            .I(N__4268));
    InMux I__821 (
            .O(N__4279),
            .I(N__4268));
    Odrv4 I__820 (
            .O(N__4276),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__819 (
            .O(N__4273),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__818 (
            .O(N__4268),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__817 (
            .O(N__4261),
            .I(N__4258));
    LocalMux I__816 (
            .O(N__4258),
            .I(N__4253));
    InMux I__815 (
            .O(N__4257),
            .I(N__4248));
    InMux I__814 (
            .O(N__4256),
            .I(N__4248));
    Sp12to4 I__813 (
            .O(N__4253),
            .I(N__4243));
    LocalMux I__812 (
            .O(N__4248),
            .I(N__4243));
    Odrv12 I__811 (
            .O(N__4243),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__810 (
            .O(N__4240),
            .I(N__4237));
    InMux I__809 (
            .O(N__4237),
            .I(N__4232));
    InMux I__808 (
            .O(N__4236),
            .I(N__4227));
    InMux I__807 (
            .O(N__4235),
            .I(N__4227));
    LocalMux I__806 (
            .O(N__4232),
            .I(N__4222));
    LocalMux I__805 (
            .O(N__4227),
            .I(N__4222));
    Span4Mux_h I__804 (
            .O(N__4222),
            .I(N__4219));
    Span4Mux_v I__803 (
            .O(N__4219),
            .I(N__4216));
    Span4Mux_h I__802 (
            .O(N__4216),
            .I(N__4213));
    Odrv4 I__801 (
            .O(N__4213),
            .I(\U409_CIA.g0Z0Z_13 ));
    InMux I__800 (
            .O(N__4210),
            .I(N__4205));
    InMux I__799 (
            .O(N__4209),
            .I(N__4200));
    InMux I__798 (
            .O(N__4208),
            .I(N__4200));
    LocalMux I__797 (
            .O(N__4205),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__796 (
            .O(N__4200),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    CascadeMux I__795 (
            .O(N__4195),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    CascadeMux I__794 (
            .O(N__4192),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__793 (
            .O(N__4189),
            .I(N__4186));
    LocalMux I__792 (
            .O(N__4186),
            .I(\U409_TICK.TICK603_11 ));
    CascadeMux I__791 (
            .O(N__4183),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__790 (
            .O(N__4180),
            .I(N__4173));
    InMux I__789 (
            .O(N__4179),
            .I(N__4173));
    InMux I__788 (
            .O(N__4178),
            .I(N__4170));
    LocalMux I__787 (
            .O(N__4173),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__786 (
            .O(N__4170),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__785 (
            .O(N__4165),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    InMux I__784 (
            .O(N__4162),
            .I(N__4156));
    InMux I__783 (
            .O(N__4161),
            .I(N__4156));
    LocalMux I__782 (
            .O(N__4156),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__781 (
            .O(N__4153),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ));
    CascadeMux I__780 (
            .O(N__4150),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__779 (
            .O(N__4147),
            .I(N__4139));
    InMux I__778 (
            .O(N__4146),
            .I(N__4139));
    InMux I__777 (
            .O(N__4145),
            .I(N__4134));
    InMux I__776 (
            .O(N__4144),
            .I(N__4134));
    LocalMux I__775 (
            .O(N__4139),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__774 (
            .O(N__4134),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__773 (
            .O(N__4129),
            .I(\U409_TRANSFER_ACK.m9_am_cascade_ ));
    CascadeMux I__772 (
            .O(N__4126),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    InMux I__771 (
            .O(N__4123),
            .I(N__4120));
    LocalMux I__770 (
            .O(N__4120),
            .I(N__4116));
    InMux I__769 (
            .O(N__4119),
            .I(N__4113));
    Span12Mux_h I__768 (
            .O(N__4116),
            .I(N__4108));
    LocalMux I__767 (
            .O(N__4113),
            .I(N__4108));
    Odrv12 I__766 (
            .O(N__4108),
            .I(CIA_ENABLEm));
    InMux I__765 (
            .O(N__4105),
            .I(N__4099));
    InMux I__764 (
            .O(N__4104),
            .I(N__4096));
    InMux I__763 (
            .O(N__4103),
            .I(N__4089));
    InMux I__762 (
            .O(N__4102),
            .I(N__4089));
    LocalMux I__761 (
            .O(N__4099),
            .I(N__4086));
    LocalMux I__760 (
            .O(N__4096),
            .I(N__4083));
    InMux I__759 (
            .O(N__4095),
            .I(N__4078));
    InMux I__758 (
            .O(N__4094),
            .I(N__4078));
    LocalMux I__757 (
            .O(N__4089),
            .I(N__4075));
    Span4Mux_v I__756 (
            .O(N__4086),
            .I(N__4068));
    Span4Mux_h I__755 (
            .O(N__4083),
            .I(N__4068));
    LocalMux I__754 (
            .O(N__4078),
            .I(N__4068));
    Sp12to4 I__753 (
            .O(N__4075),
            .I(N__4064));
    Span4Mux_v I__752 (
            .O(N__4068),
            .I(N__4061));
    InMux I__751 (
            .O(N__4067),
            .I(N__4058));
    Span12Mux_v I__750 (
            .O(N__4064),
            .I(N__4055));
    Span4Mux_v I__749 (
            .O(N__4061),
            .I(N__4052));
    LocalMux I__748 (
            .O(N__4058),
            .I(N__4049));
    Span12Mux_h I__747 (
            .O(N__4055),
            .I(N__4046));
    Sp12to4 I__746 (
            .O(N__4052),
            .I(N__4041));
    Span12Mux_v I__745 (
            .O(N__4049),
            .I(N__4041));
    Odrv12 I__744 (
            .O(N__4046),
            .I(A_c_22));
    Odrv12 I__743 (
            .O(N__4041),
            .I(A_c_22));
    CascadeMux I__742 (
            .O(N__4036),
            .I(N__4033));
    InMux I__741 (
            .O(N__4033),
            .I(N__4023));
    InMux I__740 (
            .O(N__4032),
            .I(N__4023));
    InMux I__739 (
            .O(N__4031),
            .I(N__4019));
    InMux I__738 (
            .O(N__4030),
            .I(N__4014));
    InMux I__737 (
            .O(N__4029),
            .I(N__4014));
    InMux I__736 (
            .O(N__4028),
            .I(N__4011));
    LocalMux I__735 (
            .O(N__4023),
            .I(N__4008));
    InMux I__734 (
            .O(N__4022),
            .I(N__4005));
    LocalMux I__733 (
            .O(N__4019),
            .I(N__4002));
    LocalMux I__732 (
            .O(N__4014),
            .I(N__3998));
    LocalMux I__731 (
            .O(N__4011),
            .I(N__3995));
    Span4Mux_v I__730 (
            .O(N__4008),
            .I(N__3992));
    LocalMux I__729 (
            .O(N__4005),
            .I(N__3989));
    Span4Mux_v I__728 (
            .O(N__4002),
            .I(N__3986));
    InMux I__727 (
            .O(N__4001),
            .I(N__3983));
    Sp12to4 I__726 (
            .O(N__3998),
            .I(N__3980));
    Span4Mux_v I__725 (
            .O(N__3995),
            .I(N__3977));
    Sp12to4 I__724 (
            .O(N__3992),
            .I(N__3968));
    Span12Mux_v I__723 (
            .O(N__3989),
            .I(N__3968));
    Sp12to4 I__722 (
            .O(N__3986),
            .I(N__3968));
    LocalMux I__721 (
            .O(N__3983),
            .I(N__3968));
    Span12Mux_v I__720 (
            .O(N__3980),
            .I(N__3965));
    Span4Mux_h I__719 (
            .O(N__3977),
            .I(N__3962));
    Odrv12 I__718 (
            .O(N__3968),
            .I(A_c_23));
    Odrv12 I__717 (
            .O(N__3965),
            .I(A_c_23));
    Odrv4 I__716 (
            .O(N__3962),
            .I(A_c_23));
    CascadeMux I__715 (
            .O(N__3955),
            .I(N__3951));
    InMux I__714 (
            .O(N__3954),
            .I(N__3946));
    InMux I__713 (
            .O(N__3951),
            .I(N__3946));
    LocalMux I__712 (
            .O(N__3946),
            .I(N__3940));
    CascadeMux I__711 (
            .O(N__3945),
            .I(N__3937));
    InMux I__710 (
            .O(N__3944),
            .I(N__3932));
    InMux I__709 (
            .O(N__3943),
            .I(N__3932));
    Span4Mux_v I__708 (
            .O(N__3940),
            .I(N__3929));
    InMux I__707 (
            .O(N__3937),
            .I(N__3926));
    LocalMux I__706 (
            .O(N__3932),
            .I(N__3923));
    Span4Mux_h I__705 (
            .O(N__3929),
            .I(N__3920));
    LocalMux I__704 (
            .O(N__3926),
            .I(N__3917));
    Span4Mux_v I__703 (
            .O(N__3923),
            .I(N__3914));
    Span4Mux_h I__702 (
            .O(N__3920),
            .I(N__3909));
    Span4Mux_v I__701 (
            .O(N__3917),
            .I(N__3909));
    Span4Mux_h I__700 (
            .O(N__3914),
            .I(N__3906));
    Span4Mux_h I__699 (
            .O(N__3909),
            .I(N__3903));
    Odrv4 I__698 (
            .O(N__3906),
            .I(A_c_21));
    Odrv4 I__697 (
            .O(N__3903),
            .I(A_c_21));
    InMux I__696 (
            .O(N__3898),
            .I(N__3895));
    LocalMux I__695 (
            .O(N__3895),
            .I(N__3892));
    Span4Mux_h I__694 (
            .O(N__3892),
            .I(N__3889));
    Span4Mux_h I__693 (
            .O(N__3889),
            .I(N__3886));
    Odrv4 I__692 (
            .O(N__3886),
            .I(AUTOVECTORm));
    IoInMux I__691 (
            .O(N__3883),
            .I(N__3880));
    LocalMux I__690 (
            .O(N__3880),
            .I(N__3877));
    IoSpan4Mux I__689 (
            .O(N__3877),
            .I(N__3874));
    Span4Mux_s2_v I__688 (
            .O(N__3874),
            .I(N__3871));
    Span4Mux_v I__687 (
            .O(N__3871),
            .I(N__3868));
    Span4Mux_v I__686 (
            .O(N__3868),
            .I(N__3865));
    Odrv4 I__685 (
            .O(N__3865),
            .I(ROMENm_i));
    CascadeMux I__684 (
            .O(N__3862),
            .I(N__3858));
    InMux I__683 (
            .O(N__3861),
            .I(N__3853));
    InMux I__682 (
            .O(N__3858),
            .I(N__3853));
    LocalMux I__681 (
            .O(N__3853),
            .I(N__3850));
    Odrv4 I__680 (
            .O(N__3850),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0 ));
    CascadeMux I__679 (
            .O(N__3847),
            .I(N__3844));
    InMux I__678 (
            .O(N__3844),
            .I(N__3838));
    InMux I__677 (
            .O(N__3843),
            .I(N__3838));
    LocalMux I__676 (
            .O(N__3838),
            .I(N__3835));
    Span4Mux_h I__675 (
            .O(N__3835),
            .I(N__3832));
    Odrv4 I__674 (
            .O(N__3832),
            .I(\U409_ADDRESS_DECODE.HIROMZ0 ));
    CascadeMux I__673 (
            .O(N__3829),
            .I(N__3826));
    InMux I__672 (
            .O(N__3826),
            .I(N__3823));
    LocalMux I__671 (
            .O(N__3823),
            .I(ROMENm));
    InMux I__670 (
            .O(N__3820),
            .I(N__3816));
    InMux I__669 (
            .O(N__3819),
            .I(N__3813));
    LocalMux I__668 (
            .O(N__3816),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__667 (
            .O(N__3813),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__666 (
            .O(N__3808),
            .I(N__3804));
    InMux I__665 (
            .O(N__3807),
            .I(N__3801));
    LocalMux I__664 (
            .O(N__3804),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__663 (
            .O(N__3801),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__662 (
            .O(N__3796),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__661 (
            .O(N__3793),
            .I(N__3790));
    LocalMux I__660 (
            .O(N__3790),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__659 (
            .O(N__3787),
            .I(N__3783));
    InMux I__658 (
            .O(N__3786),
            .I(N__3780));
    LocalMux I__657 (
            .O(N__3783),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__656 (
            .O(N__3780),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__655 (
            .O(N__3775),
            .I(N__3772));
    LocalMux I__654 (
            .O(N__3772),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__653 (
            .O(N__3769),
            .I(N__3765));
    InMux I__652 (
            .O(N__3768),
            .I(N__3762));
    LocalMux I__651 (
            .O(N__3765),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__650 (
            .O(N__3762),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__649 (
            .O(N__3757),
            .I(N__3754));
    InMux I__648 (
            .O(N__3754),
            .I(N__3750));
    InMux I__647 (
            .O(N__3753),
            .I(N__3747));
    LocalMux I__646 (
            .O(N__3750),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__645 (
            .O(N__3747),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__644 (
            .O(N__3742),
            .I(N__3738));
    InMux I__643 (
            .O(N__3741),
            .I(N__3735));
    LocalMux I__642 (
            .O(N__3738),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__641 (
            .O(N__3735),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__640 (
            .O(N__3730),
            .I(N__3727));
    LocalMux I__639 (
            .O(N__3727),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    CascadeMux I__638 (
            .O(N__3724),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__637 (
            .O(N__3721),
            .I(N__3718));
    InMux I__636 (
            .O(N__3718),
            .I(N__3714));
    InMux I__635 (
            .O(N__3717),
            .I(N__3711));
    LocalMux I__634 (
            .O(N__3714),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__633 (
            .O(N__3711),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__632 (
            .O(N__3706),
            .I(N__3690));
    InMux I__631 (
            .O(N__3705),
            .I(N__3690));
    InMux I__630 (
            .O(N__3704),
            .I(N__3690));
    InMux I__629 (
            .O(N__3703),
            .I(N__3690));
    InMux I__628 (
            .O(N__3702),
            .I(N__3681));
    InMux I__627 (
            .O(N__3701),
            .I(N__3681));
    InMux I__626 (
            .O(N__3700),
            .I(N__3681));
    InMux I__625 (
            .O(N__3699),
            .I(N__3681));
    LocalMux I__624 (
            .O(N__3690),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__623 (
            .O(N__3681),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__622 (
            .O(N__3676),
            .I(N__3668));
    InMux I__621 (
            .O(N__3675),
            .I(N__3655));
    InMux I__620 (
            .O(N__3674),
            .I(N__3655));
    InMux I__619 (
            .O(N__3673),
            .I(N__3655));
    InMux I__618 (
            .O(N__3672),
            .I(N__3655));
    InMux I__617 (
            .O(N__3671),
            .I(N__3655));
    InMux I__616 (
            .O(N__3668),
            .I(N__3652));
    InMux I__615 (
            .O(N__3667),
            .I(N__3647));
    InMux I__614 (
            .O(N__3666),
            .I(N__3647));
    LocalMux I__613 (
            .O(N__3655),
            .I(N__3644));
    LocalMux I__612 (
            .O(N__3652),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__611 (
            .O(N__3647),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__610 (
            .O(N__3644),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__609 (
            .O(N__3637),
            .I(N__3628));
    CascadeMux I__608 (
            .O(N__3636),
            .I(N__3625));
    CascadeMux I__607 (
            .O(N__3635),
            .I(N__3621));
    CascadeMux I__606 (
            .O(N__3634),
            .I(N__3618));
    InMux I__605 (
            .O(N__3633),
            .I(N__3609));
    InMux I__604 (
            .O(N__3632),
            .I(N__3609));
    InMux I__603 (
            .O(N__3631),
            .I(N__3609));
    InMux I__602 (
            .O(N__3628),
            .I(N__3609));
    InMux I__601 (
            .O(N__3625),
            .I(N__3606));
    InMux I__600 (
            .O(N__3624),
            .I(N__3599));
    InMux I__599 (
            .O(N__3621),
            .I(N__3599));
    InMux I__598 (
            .O(N__3618),
            .I(N__3599));
    LocalMux I__597 (
            .O(N__3609),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__596 (
            .O(N__3606),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__595 (
            .O(N__3599),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__594 (
            .O(N__3592),
            .I(N__3589));
    LocalMux I__593 (
            .O(N__3589),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__592 (
            .O(N__3586),
            .I(N__3582));
    InMux I__591 (
            .O(N__3585),
            .I(N__3579));
    LocalMux I__590 (
            .O(N__3582),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__589 (
            .O(N__3579),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    IoInMux I__588 (
            .O(N__3574),
            .I(N__3571));
    LocalMux I__587 (
            .O(N__3571),
            .I(N__3568));
    IoSpan4Mux I__586 (
            .O(N__3568),
            .I(N__3565));
    Span4Mux_s2_v I__585 (
            .O(N__3565),
            .I(N__3562));
    Sp12to4 I__584 (
            .O(N__3562),
            .I(N__3559));
    Span12Mux_s11_v I__583 (
            .O(N__3559),
            .I(N__3556));
    Odrv12 I__582 (
            .O(N__3556),
            .I(U409_ADDRESS_DECODE_un1_nRAMSPACE_i));
    ClkMux I__581 (
            .O(N__3553),
            .I(N__3541));
    ClkMux I__580 (
            .O(N__3552),
            .I(N__3541));
    ClkMux I__579 (
            .O(N__3551),
            .I(N__3541));
    ClkMux I__578 (
            .O(N__3550),
            .I(N__3541));
    GlobalMux I__577 (
            .O(N__3541),
            .I(N__3538));
    gio2CtrlBuf I__576 (
            .O(N__3538),
            .I(CLK28_IN_c_g));
    InMux I__575 (
            .O(N__3535),
            .I(N__3531));
    InMux I__574 (
            .O(N__3534),
            .I(N__3528));
    LocalMux I__573 (
            .O(N__3531),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__572 (
            .O(N__3528),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__571 (
            .O(N__3523),
            .I(N__3519));
    InMux I__570 (
            .O(N__3522),
            .I(N__3516));
    LocalMux I__569 (
            .O(N__3519),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__568 (
            .O(N__3516),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    CascadeMux I__567 (
            .O(N__3511),
            .I(N__3507));
    InMux I__566 (
            .O(N__3510),
            .I(N__3504));
    InMux I__565 (
            .O(N__3507),
            .I(N__3501));
    LocalMux I__564 (
            .O(N__3504),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__563 (
            .O(N__3501),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__562 (
            .O(N__3496),
            .I(N__3492));
    InMux I__561 (
            .O(N__3495),
            .I(N__3489));
    LocalMux I__560 (
            .O(N__3492),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__559 (
            .O(N__3489),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__558 (
            .O(N__3484),
            .I(N__3481));
    LocalMux I__557 (
            .O(N__3481),
            .I(\U409_TICK.TICK503_11 ));
    InMux I__556 (
            .O(N__3478),
            .I(N__3474));
    InMux I__555 (
            .O(N__3477),
            .I(N__3471));
    LocalMux I__554 (
            .O(N__3474),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__553 (
            .O(N__3471),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__552 (
            .O(N__3466),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__551 (
            .O(N__3463),
            .I(N__3459));
    InMux I__550 (
            .O(N__3462),
            .I(N__3456));
    LocalMux I__549 (
            .O(N__3459),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__548 (
            .O(N__3456),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    CascadeMux I__547 (
            .O(N__3451),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    IoInMux I__546 (
            .O(N__3448),
            .I(N__3445));
    LocalMux I__545 (
            .O(N__3445),
            .I(N__3442));
    Span4Mux_s1_v I__544 (
            .O(N__3442),
            .I(N__3439));
    Sp12to4 I__543 (
            .O(N__3439),
            .I(N__3436));
    Span12Mux_h I__542 (
            .O(N__3436),
            .I(N__3433));
    Span12Mux_v I__541 (
            .O(N__3433),
            .I(N__3429));
    InMux I__540 (
            .O(N__3432),
            .I(N__3426));
    Odrv12 I__539 (
            .O(N__3429),
            .I(TICK50_c));
    LocalMux I__538 (
            .O(N__3426),
            .I(TICK50_c));
    InMux I__537 (
            .O(N__3421),
            .I(N__3418));
    LocalMux I__536 (
            .O(N__3418),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    CascadeMux I__535 (
            .O(N__3415),
            .I(N__3411));
    CascadeMux I__534 (
            .O(N__3414),
            .I(N__3406));
    InMux I__533 (
            .O(N__3411),
            .I(N__3403));
    InMux I__532 (
            .O(N__3410),
            .I(N__3398));
    InMux I__531 (
            .O(N__3409),
            .I(N__3398));
    InMux I__530 (
            .O(N__3406),
            .I(N__3395));
    LocalMux I__529 (
            .O(N__3403),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__528 (
            .O(N__3398),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__527 (
            .O(N__3395),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__526 (
            .O(N__3388),
            .I(N__3381));
    InMux I__525 (
            .O(N__3387),
            .I(N__3381));
    InMux I__524 (
            .O(N__3386),
            .I(N__3378));
    LocalMux I__523 (
            .O(N__3381),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__522 (
            .O(N__3378),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__521 (
            .O(N__3373),
            .I(N__3370));
    LocalMux I__520 (
            .O(N__3370),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__519 (
            .O(N__3367),
            .I(N__3363));
    InMux I__518 (
            .O(N__3366),
            .I(N__3360));
    LocalMux I__517 (
            .O(N__3363),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__516 (
            .O(N__3360),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__515 (
            .O(N__3355),
            .I(N__3352));
    LocalMux I__514 (
            .O(N__3352),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__513 (
            .O(N__3349),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__512 (
            .O(N__3346),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__511 (
            .O(N__3343),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__510 (
            .O(N__3340),
            .I(N__3332));
    InMux I__509 (
            .O(N__3339),
            .I(N__3332));
    InMux I__508 (
            .O(N__3338),
            .I(N__3327));
    InMux I__507 (
            .O(N__3337),
            .I(N__3327));
    LocalMux I__506 (
            .O(N__3332),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__505 (
            .O(N__3327),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__504 (
            .O(N__3322),
            .I(N__3317));
    InMux I__503 (
            .O(N__3321),
            .I(N__3311));
    InMux I__502 (
            .O(N__3320),
            .I(N__3311));
    InMux I__501 (
            .O(N__3317),
            .I(N__3306));
    InMux I__500 (
            .O(N__3316),
            .I(N__3306));
    LocalMux I__499 (
            .O(N__3311),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__498 (
            .O(N__3306),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__497 (
            .O(N__3301),
            .I(N__3297));
    InMux I__496 (
            .O(N__3300),
            .I(N__3292));
    InMux I__495 (
            .O(N__3297),
            .I(N__3287));
    InMux I__494 (
            .O(N__3296),
            .I(N__3287));
    InMux I__493 (
            .O(N__3295),
            .I(N__3284));
    LocalMux I__492 (
            .O(N__3292),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__491 (
            .O(N__3287),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__490 (
            .O(N__3284),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__489 (
            .O(N__3277),
            .I(N__3269));
    InMux I__488 (
            .O(N__3276),
            .I(N__3262));
    InMux I__487 (
            .O(N__3275),
            .I(N__3262));
    InMux I__486 (
            .O(N__3274),
            .I(N__3262));
    InMux I__485 (
            .O(N__3273),
            .I(N__3257));
    InMux I__484 (
            .O(N__3272),
            .I(N__3257));
    LocalMux I__483 (
            .O(N__3269),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__482 (
            .O(N__3262),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__481 (
            .O(N__3257),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__480 (
            .O(N__3250),
            .I(N__3247));
    LocalMux I__479 (
            .O(N__3247),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    InMux I__478 (
            .O(N__3244),
            .I(N__3241));
    LocalMux I__477 (
            .O(N__3241),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__476 (
            .O(N__3238),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ));
    CascadeMux I__475 (
            .O(N__3235),
            .I(N__3225));
    InMux I__474 (
            .O(N__3234),
            .I(N__3220));
    InMux I__473 (
            .O(N__3233),
            .I(N__3220));
    InMux I__472 (
            .O(N__3232),
            .I(N__3217));
    InMux I__471 (
            .O(N__3231),
            .I(N__3212));
    InMux I__470 (
            .O(N__3230),
            .I(N__3212));
    InMux I__469 (
            .O(N__3229),
            .I(N__3205));
    InMux I__468 (
            .O(N__3228),
            .I(N__3205));
    InMux I__467 (
            .O(N__3225),
            .I(N__3205));
    LocalMux I__466 (
            .O(N__3220),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__465 (
            .O(N__3217),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__464 (
            .O(N__3212),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__463 (
            .O(N__3205),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__462 (
            .O(N__3196),
            .I(N__3187));
    InMux I__461 (
            .O(N__3195),
            .I(N__3180));
    InMux I__460 (
            .O(N__3194),
            .I(N__3180));
    InMux I__459 (
            .O(N__3193),
            .I(N__3180));
    InMux I__458 (
            .O(N__3192),
            .I(N__3173));
    InMux I__457 (
            .O(N__3191),
            .I(N__3173));
    InMux I__456 (
            .O(N__3190),
            .I(N__3173));
    LocalMux I__455 (
            .O(N__3187),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__454 (
            .O(N__3180),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__453 (
            .O(N__3173),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__452 (
            .O(N__3166),
            .I(N__3163));
    LocalMux I__451 (
            .O(N__3163),
            .I(N__3159));
    InMux I__450 (
            .O(N__3162),
            .I(N__3156));
    Span12Mux_v I__449 (
            .O(N__3159),
            .I(N__3151));
    LocalMux I__448 (
            .O(N__3156),
            .I(N__3151));
    Odrv12 I__447 (
            .O(N__3151),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    IoInMux I__446 (
            .O(N__3148),
            .I(N__3145));
    LocalMux I__445 (
            .O(N__3145),
            .I(N__3142));
    IoSpan4Mux I__444 (
            .O(N__3142),
            .I(N__3139));
    Span4Mux_s3_v I__443 (
            .O(N__3139),
            .I(N__3136));
    Sp12to4 I__442 (
            .O(N__3136),
            .I(N__3133));
    Span12Mux_s11_v I__441 (
            .O(N__3133),
            .I(N__3130));
    Odrv12 I__440 (
            .O(N__3130),
            .I(U409_ADDRESS_DECODE_un1_nREGSPACE_i));
    InMux I__439 (
            .O(N__3127),
            .I(N__3124));
    LocalMux I__438 (
            .O(N__3124),
            .I(N__3121));
    Span4Mux_v I__437 (
            .O(N__3121),
            .I(N__3118));
    Sp12to4 I__436 (
            .O(N__3118),
            .I(N__3115));
    Span12Mux_h I__435 (
            .O(N__3115),
            .I(N__3112));
    Odrv12 I__434 (
            .O(N__3112),
            .I(A_c_13));
    IoInMux I__433 (
            .O(N__3109),
            .I(N__3106));
    LocalMux I__432 (
            .O(N__3106),
            .I(N__3103));
    Span4Mux_s1_h I__431 (
            .O(N__3103),
            .I(N__3100));
    Sp12to4 I__430 (
            .O(N__3100),
            .I(N__3097));
    Span12Mux_s9_v I__429 (
            .O(N__3097),
            .I(N__3094));
    Span12Mux_h I__428 (
            .O(N__3094),
            .I(N__3091));
    Odrv12 I__427 (
            .O(N__3091),
            .I(U409_ADDRESS_DECODE_un1_nCIACS1_i));
    InMux I__426 (
            .O(N__3088),
            .I(N__3085));
    LocalMux I__425 (
            .O(N__3085),
            .I(N__3082));
    Span12Mux_h I__424 (
            .O(N__3082),
            .I(N__3079));
    Odrv12 I__423 (
            .O(N__3079),
            .I(A_c_12));
    IoInMux I__422 (
            .O(N__3076),
            .I(N__3073));
    LocalMux I__421 (
            .O(N__3073),
            .I(N__3070));
    Span4Mux_s1_h I__420 (
            .O(N__3070),
            .I(N__3067));
    Sp12to4 I__419 (
            .O(N__3067),
            .I(N__3064));
    Span12Mux_s10_v I__418 (
            .O(N__3064),
            .I(N__3061));
    Span12Mux_h I__417 (
            .O(N__3061),
            .I(N__3058));
    Odrv12 I__416 (
            .O(N__3058),
            .I(U409_ADDRESS_DECODE_un1_nCIACS0_i));
    CascadeMux I__415 (
            .O(N__3055),
            .I(\U409_CIA.N_9_cascade_ ));
    CascadeMux I__414 (
            .O(N__3052),
            .I(\U409_CIA.N_20_cascade_ ));
    InMux I__413 (
            .O(N__3049),
            .I(N__3043));
    InMux I__412 (
            .O(N__3048),
            .I(N__3043));
    LocalMux I__411 (
            .O(N__3043),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    InMux I__410 (
            .O(N__3040),
            .I(N__3037));
    LocalMux I__409 (
            .O(N__3037),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__408 (
            .O(N__3034),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    InMux I__407 (
            .O(N__3031),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__406 (
            .O(N__3028),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__405 (
            .O(N__3025),
            .I(bfn_8_9_0_));
    InMux I__404 (
            .O(N__3022),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__403 (
            .O(N__3019),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__402 (
            .O(N__3016),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__401 (
            .O(N__3013),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__400 (
            .O(N__3010),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__399 (
            .O(N__3007),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__398 (
            .O(N__3004),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__397 (
            .O(N__3001),
            .I(N__2998));
    LocalMux I__396 (
            .O(N__2998),
            .I(N__2995));
    Span4Mux_h I__395 (
            .O(N__2995),
            .I(N__2992));
    Odrv4 I__394 (
            .O(N__2992),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    IoInMux I__393 (
            .O(N__2989),
            .I(N__2986));
    LocalMux I__392 (
            .O(N__2986),
            .I(N__2983));
    IoSpan4Mux I__391 (
            .O(N__2983),
            .I(N__2980));
    Sp12to4 I__390 (
            .O(N__2980),
            .I(N__2977));
    Span12Mux_v I__389 (
            .O(N__2977),
            .I(N__2974));
    Odrv12 I__388 (
            .O(N__2974),
            .I(PORTSIZE_0_i));
    InMux I__387 (
            .O(N__2971),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__386 (
            .O(N__2968),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__385 (
            .O(N__2965),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__384 (
            .O(N__2962),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__383 (
            .O(N__2959),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__382 (
            .O(N__2956),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__381 (
            .O(N__2953),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__380 (
            .O(N__2950),
            .I(N__2941));
    InMux I__379 (
            .O(N__2949),
            .I(N__2941));
    InMux I__378 (
            .O(N__2948),
            .I(N__2941));
    LocalMux I__377 (
            .O(N__2941),
            .I(N__2938));
    Span12Mux_v I__376 (
            .O(N__2938),
            .I(N__2935));
    Odrv12 I__375 (
            .O(N__2935),
            .I(A_c_29));
    InMux I__374 (
            .O(N__2932),
            .I(N__2927));
    InMux I__373 (
            .O(N__2931),
            .I(N__2922));
    InMux I__372 (
            .O(N__2930),
            .I(N__2922));
    LocalMux I__371 (
            .O(N__2927),
            .I(N__2917));
    LocalMux I__370 (
            .O(N__2922),
            .I(N__2917));
    Span4Mux_h I__369 (
            .O(N__2917),
            .I(N__2914));
    Span4Mux_v I__368 (
            .O(N__2914),
            .I(N__2911));
    Span4Mux_v I__367 (
            .O(N__2911),
            .I(N__2908));
    Odrv4 I__366 (
            .O(N__2908),
            .I(A_c_28));
    CascadeMux I__365 (
            .O(N__2905),
            .I(N__2902));
    InMux I__364 (
            .O(N__2902),
            .I(N__2897));
    InMux I__363 (
            .O(N__2901),
            .I(N__2894));
    InMux I__362 (
            .O(N__2900),
            .I(N__2891));
    LocalMux I__361 (
            .O(N__2897),
            .I(N__2884));
    LocalMux I__360 (
            .O(N__2894),
            .I(N__2884));
    LocalMux I__359 (
            .O(N__2891),
            .I(N__2884));
    Odrv12 I__358 (
            .O(N__2884),
            .I(A_c_27));
    CascadeMux I__357 (
            .O(N__2881),
            .I(N__2877));
    InMux I__356 (
            .O(N__2880),
            .I(N__2869));
    InMux I__355 (
            .O(N__2877),
            .I(N__2869));
    InMux I__354 (
            .O(N__2876),
            .I(N__2869));
    LocalMux I__353 (
            .O(N__2869),
            .I(N__2866));
    Span12Mux_v I__352 (
            .O(N__2866),
            .I(N__2863));
    Odrv12 I__351 (
            .O(N__2863),
            .I(A_c_30));
    InMux I__350 (
            .O(N__2860),
            .I(N__2857));
    LocalMux I__349 (
            .O(N__2857),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ));
    InMux I__348 (
            .O(N__2854),
            .I(N__2848));
    InMux I__347 (
            .O(N__2853),
            .I(N__2848));
    LocalMux I__346 (
            .O(N__2848),
            .I(N__2845));
    Span4Mux_v I__345 (
            .O(N__2845),
            .I(N__2841));
    InMux I__344 (
            .O(N__2844),
            .I(N__2838));
    Sp12to4 I__343 (
            .O(N__2841),
            .I(N__2833));
    LocalMux I__342 (
            .O(N__2838),
            .I(N__2833));
    Odrv12 I__341 (
            .O(N__2833),
            .I(A_c_20));
    CascadeMux I__340 (
            .O(N__2830),
            .I(N__2826));
    InMux I__339 (
            .O(N__2829),
            .I(N__2822));
    InMux I__338 (
            .O(N__2826),
            .I(N__2819));
    InMux I__337 (
            .O(N__2825),
            .I(N__2816));
    LocalMux I__336 (
            .O(N__2822),
            .I(N__2811));
    LocalMux I__335 (
            .O(N__2819),
            .I(N__2811));
    LocalMux I__334 (
            .O(N__2816),
            .I(N__2808));
    Span4Mux_v I__333 (
            .O(N__2811),
            .I(N__2805));
    Odrv12 I__332 (
            .O(N__2808),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    Odrv4 I__331 (
            .O(N__2805),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    InMux I__330 (
            .O(N__2800),
            .I(N__2795));
    InMux I__329 (
            .O(N__2799),
            .I(N__2790));
    InMux I__328 (
            .O(N__2798),
            .I(N__2790));
    LocalMux I__327 (
            .O(N__2795),
            .I(N__2787));
    LocalMux I__326 (
            .O(N__2790),
            .I(N__2784));
    Span4Mux_v I__325 (
            .O(N__2787),
            .I(N__2781));
    Span4Mux_v I__324 (
            .O(N__2784),
            .I(N__2778));
    Span4Mux_h I__323 (
            .O(N__2781),
            .I(N__2775));
    Sp12to4 I__322 (
            .O(N__2778),
            .I(N__2772));
    Sp12to4 I__321 (
            .O(N__2775),
            .I(N__2767));
    Span12Mux_s3_h I__320 (
            .O(N__2772),
            .I(N__2767));
    Span12Mux_v I__319 (
            .O(N__2767),
            .I(N__2764));
    Odrv12 I__318 (
            .O(N__2764),
            .I(A_c_19));
    CascadeMux I__317 (
            .O(N__2761),
            .I(N__2757));
    CascadeMux I__316 (
            .O(N__2760),
            .I(N__2754));
    InMux I__315 (
            .O(N__2757),
            .I(N__2748));
    InMux I__314 (
            .O(N__2754),
            .I(N__2748));
    CascadeMux I__313 (
            .O(N__2753),
            .I(N__2745));
    LocalMux I__312 (
            .O(N__2748),
            .I(N__2742));
    InMux I__311 (
            .O(N__2745),
            .I(N__2739));
    Odrv4 I__310 (
            .O(N__2742),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_3 ));
    LocalMux I__309 (
            .O(N__2739),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_3 ));
    InMux I__308 (
            .O(N__2734),
            .I(N__2731));
    LocalMux I__307 (
            .O(N__2731),
            .I(N__2728));
    Span4Mux_v I__306 (
            .O(N__2728),
            .I(N__2725));
    Span4Mux_v I__305 (
            .O(N__2725),
            .I(N__2722));
    IoSpan4Mux I__304 (
            .O(N__2722),
            .I(N__2719));
    Odrv4 I__303 (
            .O(N__2719),
            .I(TT_c_1));
    InMux I__302 (
            .O(N__2716),
            .I(N__2713));
    LocalMux I__301 (
            .O(N__2713),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ));
    InMux I__300 (
            .O(N__2710),
            .I(N__2707));
    LocalMux I__299 (
            .O(N__2707),
            .I(N__2704));
    Span4Mux_h I__298 (
            .O(N__2704),
            .I(N__2701));
    Span4Mux_v I__297 (
            .O(N__2701),
            .I(N__2696));
    InMux I__296 (
            .O(N__2700),
            .I(N__2691));
    InMux I__295 (
            .O(N__2699),
            .I(N__2691));
    Sp12to4 I__294 (
            .O(N__2696),
            .I(N__2686));
    LocalMux I__293 (
            .O(N__2691),
            .I(N__2686));
    Odrv12 I__292 (
            .O(N__2686),
            .I(A_c_25));
    CascadeMux I__291 (
            .O(N__2683),
            .I(N__2679));
    CascadeMux I__290 (
            .O(N__2682),
            .I(N__2675));
    InMux I__289 (
            .O(N__2679),
            .I(N__2672));
    InMux I__288 (
            .O(N__2678),
            .I(N__2667));
    InMux I__287 (
            .O(N__2675),
            .I(N__2667));
    LocalMux I__286 (
            .O(N__2672),
            .I(N__2662));
    LocalMux I__285 (
            .O(N__2667),
            .I(N__2662));
    Span4Mux_v I__284 (
            .O(N__2662),
            .I(N__2659));
    Span4Mux_v I__283 (
            .O(N__2659),
            .I(N__2656));
    Sp12to4 I__282 (
            .O(N__2656),
            .I(N__2653));
    Odrv12 I__281 (
            .O(N__2653),
            .I(A_c_24));
    InMux I__280 (
            .O(N__2650),
            .I(N__2641));
    InMux I__279 (
            .O(N__2649),
            .I(N__2641));
    InMux I__278 (
            .O(N__2648),
            .I(N__2641));
    LocalMux I__277 (
            .O(N__2641),
            .I(N__2638));
    Span4Mux_v I__276 (
            .O(N__2638),
            .I(N__2635));
    Span4Mux_v I__275 (
            .O(N__2635),
            .I(N__2632));
    Span4Mux_h I__274 (
            .O(N__2632),
            .I(N__2629));
    Odrv4 I__273 (
            .O(N__2629),
            .I(A_c_26));
    CascadeMux I__272 (
            .O(N__2626),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ));
    InMux I__271 (
            .O(N__2623),
            .I(N__2620));
    LocalMux I__270 (
            .O(N__2620),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    InMux I__269 (
            .O(N__2617),
            .I(N__2614));
    LocalMux I__268 (
            .O(N__2614),
            .I(N__2611));
    Span12Mux_v I__267 (
            .O(N__2611),
            .I(N__2608));
    Odrv12 I__266 (
            .O(N__2608),
            .I(TT_c_0));
    CascadeMux I__265 (
            .O(N__2605),
            .I(N__2600));
    InMux I__264 (
            .O(N__2604),
            .I(N__2595));
    InMux I__263 (
            .O(N__2603),
            .I(N__2595));
    InMux I__262 (
            .O(N__2600),
            .I(N__2592));
    LocalMux I__261 (
            .O(N__2595),
            .I(N__2589));
    LocalMux I__260 (
            .O(N__2592),
            .I(N__2586));
    Span4Mux_v I__259 (
            .O(N__2589),
            .I(N__2583));
    Span4Mux_v I__258 (
            .O(N__2586),
            .I(N__2580));
    Sp12to4 I__257 (
            .O(N__2583),
            .I(N__2575));
    Sp12to4 I__256 (
            .O(N__2580),
            .I(N__2575));
    Odrv12 I__255 (
            .O(N__2575),
            .I(A_c_31));
    InMux I__254 (
            .O(N__2572),
            .I(N__2569));
    LocalMux I__253 (
            .O(N__2569),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ));
    CascadeMux I__252 (
            .O(N__2566),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ));
    InMux I__251 (
            .O(N__2563),
            .I(N__2560));
    LocalMux I__250 (
            .O(N__2560),
            .I(\U409_CIA.g0Z0Z_10 ));
    CascadeMux I__249 (
            .O(N__2557),
            .I(\U409_CIA.g0Z0Z_2_cascade_ ));
    InMux I__248 (
            .O(N__2554),
            .I(N__2548));
    InMux I__247 (
            .O(N__2553),
            .I(N__2548));
    LocalMux I__246 (
            .O(N__2548),
            .I(N__2545));
    Span4Mux_v I__245 (
            .O(N__2545),
            .I(N__2542));
    Sp12to4 I__244 (
            .O(N__2542),
            .I(N__2539));
    Span12Mux_s7_h I__243 (
            .O(N__2539),
            .I(N__2536));
    Span12Mux_v I__242 (
            .O(N__2536),
            .I(N__2533));
    Odrv12 I__241 (
            .O(N__2533),
            .I(A_c_18));
    CascadeMux I__240 (
            .O(N__2530),
            .I(N__2526));
    InMux I__239 (
            .O(N__2529),
            .I(N__2521));
    InMux I__238 (
            .O(N__2526),
            .I(N__2521));
    LocalMux I__237 (
            .O(N__2521),
            .I(N__2518));
    Span4Mux_v I__236 (
            .O(N__2518),
            .I(N__2515));
    Sp12to4 I__235 (
            .O(N__2515),
            .I(N__2512));
    Span12Mux_v I__234 (
            .O(N__2512),
            .I(N__2509));
    Odrv12 I__233 (
            .O(N__2509),
            .I(A_c_17));
    InMux I__232 (
            .O(N__2506),
            .I(N__2500));
    InMux I__231 (
            .O(N__2505),
            .I(N__2500));
    LocalMux I__230 (
            .O(N__2500),
            .I(N__2497));
    Span4Mux_v I__229 (
            .O(N__2497),
            .I(N__2494));
    Sp12to4 I__228 (
            .O(N__2494),
            .I(N__2491));
    Span12Mux_s3_h I__227 (
            .O(N__2491),
            .I(N__2488));
    Span12Mux_v I__226 (
            .O(N__2488),
            .I(N__2485));
    Odrv12 I__225 (
            .O(N__2485),
            .I(A_c_16));
    CascadeMux I__224 (
            .O(N__2482),
            .I(\U409_CIA.g0Z0Z_8_cascade_ ));
    InMux I__223 (
            .O(N__2479),
            .I(N__2476));
    LocalMux I__222 (
            .O(N__2476),
            .I(\U409_CIA.g0Z0Z_11 ));
    ClkMux I__221 (
            .O(N__2473),
            .I(N__2446));
    ClkMux I__220 (
            .O(N__2472),
            .I(N__2446));
    ClkMux I__219 (
            .O(N__2471),
            .I(N__2446));
    ClkMux I__218 (
            .O(N__2470),
            .I(N__2446));
    ClkMux I__217 (
            .O(N__2469),
            .I(N__2446));
    ClkMux I__216 (
            .O(N__2468),
            .I(N__2446));
    ClkMux I__215 (
            .O(N__2467),
            .I(N__2446));
    ClkMux I__214 (
            .O(N__2466),
            .I(N__2446));
    ClkMux I__213 (
            .O(N__2465),
            .I(N__2446));
    GlobalMux I__212 (
            .O(N__2446),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2468));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__2466));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__2465));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__2472));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2470));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2467));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2473));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2471));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .I(N__2469));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_12_2  (
            .in0(N__2798),
            .in1(N__2553),
            .in2(N__2530),
            .in3(N__2505),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_12_4 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_12_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_12_4  (
            .in0(N__2710),
            .in1(N__2844),
            .in2(N__3945),
            .in3(N__2554),
            .lcout(\U409_CIA.g0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_1_12_6 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_1_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_CIA.g0_8_LC_1_12_6  (
            .in0(N__2529),
            .in1(N__4028),
            .in2(_gnd_net_),
            .in3(N__5857),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_1_12_7 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_1_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_1_12_7  (
            .in0(N__2506),
            .in1(N__2799),
            .in2(N__2482),
            .in3(N__2479),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_16_2  (
            .in0(N__2648),
            .in1(N__2699),
            .in2(N__2682),
            .in3(N__2825),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_16_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_16_3  (
            .in0(N__2901),
            .in1(N__2678),
            .in2(N__2605),
            .in3(N__2650),
            .lcout(\U409_CIA.g0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_5  (
            .in0(N__2700),
            .in1(N__2900),
            .in2(N__2683),
            .in3(N__2649),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_2_16_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_2_16_0 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_2_16_0  (
            .in0(N__2604),
            .in1(_gnd_net_),
            .in2(N__2881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_2_16_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_2_16_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_2_16_1  (
            .in0(N__2949),
            .in1(N__2931),
            .in2(N__2626),
            .in3(N__2623),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_2_16_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_2_16_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_2_16_3  (
            .in0(N__5860),
            .in1(N__2617),
            .in2(_gnd_net_),
            .in3(N__2603),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_2_16_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_2_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_LC_2_16_4  (
            .in0(N__2860),
            .in1(N__2572),
            .in2(N__2566),
            .in3(N__2716),
            .lcout(AUTOVECTORm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_2_16_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_2_16_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.g0_2_LC_2_16_5  (
            .in0(N__2950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2880),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_2_16_6 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_2_16_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.g0_13_LC_2_16_6  (
            .in0(N__2563),
            .in1(N__2932),
            .in2(N__2557),
            .in3(N__4067),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_2_16_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_2_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_2_16_7  (
            .in0(N__2948),
            .in1(N__2930),
            .in2(N__2905),
            .in3(N__2876),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_3_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_3_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_0_LC_3_13_2  (
            .in0(N__3943),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2853),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_3_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_3_13_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_3_13_3  (
            .in0(N__2854),
            .in1(N__4105),
            .in2(N__2830),
            .in3(N__3944),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_3_14_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_3_14_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_3_14_6  (
            .in0(N__4104),
            .in1(N__4367),
            .in2(N__2753),
            .in3(N__2829),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_3_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_3_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_3_16_2  (
            .in0(N__4095),
            .in1(N__4030),
            .in2(N__2761),
            .in3(N__2800),
            .lcout(\U409_ADDRESS_DECODE.HIROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_16_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_16_6  (
            .in0(N__4094),
            .in1(N__4029),
            .in2(N__2760),
            .in3(N__2734),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_13_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_7_13_4  (
            .in0(N__4390),
            .in1(N__4031),
            .in2(_gnd_net_),
            .in3(N__3162),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_7_13_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3233),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3553),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_13_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__3234),
            .in2(_gnd_net_),
            .in3(N__3277),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3553),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_14_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_14_5  (
            .in0(N__5856),
            .in1(N__4001),
            .in2(N__4437),
            .in3(N__3001),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_8_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__3386),
            .in2(N__3414),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_8_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__3522),
            .in2(_gnd_net_),
            .in3(N__2971),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__5321),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_8_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__3495),
            .in2(_gnd_net_),
            .in3(N__2968),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__5321),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_8_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__3753),
            .in2(_gnd_net_),
            .in3(N__2965),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__5321),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_8_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__3366),
            .in2(_gnd_net_),
            .in3(N__2962),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_8_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__3807),
            .in2(_gnd_net_),
            .in3(N__2959),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_8_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_8_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__3768),
            .in2(_gnd_net_),
            .in3(N__2956),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__5321),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_8_8_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_8_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__3534),
            .in2(_gnd_net_),
            .in3(N__2953),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__5321),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_9_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_8_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__3717),
            .in2(_gnd_net_),
            .in3(N__3025),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_8_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__3462),
            .in2(_gnd_net_),
            .in3(N__3022),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__5323),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__3819),
            .in2(_gnd_net_),
            .in3(N__3019),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_8_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_8_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__3477),
            .in2(_gnd_net_),
            .in3(N__3016),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__5323),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_8_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__3786),
            .in2(_gnd_net_),
            .in3(N__3013),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_8_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__3585),
            .in2(_gnd_net_),
            .in3(N__3010),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_8_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__3741),
            .in2(_gnd_net_),
            .in3(N__3007),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_8_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_8_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__3510),
            .in2(_gnd_net_),
            .in3(N__3004),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5323),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_8_12_0  (
            .in0(N__3300),
            .in1(N__3340),
            .in2(N__3322),
            .in3(N__3195),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_8_12_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_8_12_2 .LUT_INIT=16'b0010001001000100;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_8_12_2  (
            .in0(N__3275),
            .in1(N__3194),
            .in2(_gnd_net_),
            .in3(N__3232),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_8_12_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_8_12_3 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \U409_CIA.VMA_LC_8_12_3  (
            .in0(N__3049),
            .in1(N__4285),
            .in2(N__3055),
            .in3(N__3196),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3551),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_12_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_12_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_12_4  (
            .in0(N__3316),
            .in1(N__3339),
            .in2(_gnd_net_),
            .in3(N__3295),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_12_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_12_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_8_12_5  (
            .in0(N__3193),
            .in1(N__3230),
            .in2(_gnd_net_),
            .in3(N__3274),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_12_6 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__4928),
            .in2(N__3052),
            .in3(N__3048),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_8_12_7 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_8_12_7 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_8_12_7  (
            .in0(N__3040),
            .in1(N__3231),
            .in2(N__3034),
            .in3(N__3276),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3551),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_13_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__3272),
            .in2(N__3235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_13_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__3337),
            .in2(_gnd_net_),
            .in3(N__3031),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__3552),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_8_13_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_8_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__3190),
            .in2(_gnd_net_),
            .in3(N__3028),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_13_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__3296),
            .in2(_gnd_net_),
            .in3(N__3349),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__3552),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_8_13_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_8_13_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__3320),
            .in2(_gnd_net_),
            .in3(N__3346),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_13_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_8_13_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_8_13_5  (
            .in0(N__3192),
            .in1(N__3250),
            .in2(N__3343),
            .in3(N__3228),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3552),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_8_13_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_8_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_8_13_6  (
            .in0(N__3338),
            .in1(N__3321),
            .in2(N__3301),
            .in3(N__3273),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_13_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_8_13_7 .LUT_INIT=16'b0010011001100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_8_13_7  (
            .in0(N__3191),
            .in1(N__3244),
            .in2(N__3238),
            .in3(N__3229),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3552),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_8_15_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_8_15_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_8_15_4  (
            .in0(N__3166),
            .in1(N__4022),
            .in2(_gnd_net_),
            .in3(N__4395),
            .lcout(U409_ADDRESS_DECODE_un1_nREGSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2  (
            .in0(N__3127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4123),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_5_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_5_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__3088),
            .in2(_gnd_net_),
            .in3(N__4119),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_8_0  (
            .in0(N__3535),
            .in1(N__3523),
            .in2(N__3511),
            .in3(N__3387),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_9_8_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_9_8_1  (
            .in0(N__3367),
            .in1(N__3496),
            .in2(_gnd_net_),
            .in3(N__3409),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_9_8_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_9_8_2  (
            .in0(N__3484),
            .in1(N__3478),
            .in2(N__3466),
            .in3(N__3463),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_9_8_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_9_8_3  (
            .in0(N__3706),
            .in1(N__3432),
            .in2(N__3451),
            .in3(N__3633),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5320),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_9_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_9_8_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_9_8_4  (
            .in0(N__3666),
            .in1(N__3705),
            .in2(N__3637),
            .in3(N__3421),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5320),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_9_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_9_8_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_9_8_5  (
            .in0(N__3703),
            .in1(N__3667),
            .in2(N__3415),
            .in3(N__3631),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5320),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_9_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_9_8_6  (
            .in0(N__3410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3388),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5320),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_9_8_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_9_8_7  (
            .in0(N__3704),
            .in1(N__3373),
            .in2(N__3676),
            .in3(N__3632),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5320),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_9_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_9_9_0  (
            .in0(N__3671),
            .in1(N__3699),
            .in2(N__3636),
            .in3(N__3355),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5322),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_9_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_9_9_1  (
            .in0(N__3820),
            .in1(N__3808),
            .in2(N__3721),
            .in3(N__3787),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_9_9_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_9_9_2  (
            .in0(N__3672),
            .in1(N__3700),
            .in2(N__3796),
            .in3(N__3793),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5322),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_9_9_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_9_9_3  (
            .in0(N__3702),
            .in1(N__3674),
            .in2(N__3635),
            .in3(N__3775),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5322),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_9_9_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_9_9_4  (
            .in0(N__3586),
            .in1(N__3769),
            .in2(N__3757),
            .in3(N__3742),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_9_9_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_9_9_5  (
            .in0(N__3624),
            .in1(N__3730),
            .in2(N__3724),
            .in3(N__3675),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5322),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_9_9_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_9_9_7  (
            .in0(N__3701),
            .in1(N__3673),
            .in2(N__3634),
            .in3(N__3592),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5322),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_9_11_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_9_11_7 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_9_11_7  (
            .in0(N__4394),
            .in1(N__4419),
            .in2(_gnd_net_),
            .in3(N__4317),
            .lcout(U409_ADDRESS_DECODE_un1_nRAMSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_9_12_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_9_12_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_9_12_0  (
            .in0(N__4235),
            .in1(N__4256),
            .in2(N__4289),
            .in3(N__4208),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3550),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_12_4 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_12_4  (
            .in0(N__4236),
            .in1(N__4257),
            .in2(N__4290),
            .in3(N__4209),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_9_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_9_13_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_LC_9_13_3  (
            .in0(N__4324),
            .in1(N__4032),
            .in2(N__3955),
            .in3(N__4102),
            .lcout(\U409_ADDRESS_DECODE.LOWROMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_9_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_9_13_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_9_13_6  (
            .in0(N__4103),
            .in1(_gnd_net_),
            .in2(N__4036),
            .in3(N__3954),
            .lcout(\U409_ADDRESS_DECODE.un5_nRAMSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_15_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_15_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_15_7  (
            .in0(N__4840),
            .in1(N__3898),
            .in2(N__3829),
            .in3(N__5100),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_16_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_9_16_4 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_9_16_4  (
            .in0(N__4386),
            .in1(N__3861),
            .in2(N__3847),
            .in3(N__5859),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_9_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_LC_9_16_5 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_LC_9_16_5  (
            .in0(N__5858),
            .in1(N__4385),
            .in2(N__3862),
            .in3(N__3843),
            .lcout(ROMENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_0  (
            .in0(N__4180),
            .in1(N__4145),
            .in2(N__4453),
            .in3(N__4627),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5668));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__4734),
            .in2(_gnd_net_),
            .in3(N__4798),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_9_2  (
            .in0(N__4662),
            .in1(N__4684),
            .in2(N__4606),
            .in3(N__4178),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_9_3  (
            .in0(N__4765),
            .in1(N__4146),
            .in2(N__4183),
            .in3(N__4161),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_9_4  (
            .in0(N__4179),
            .in1(N__4685),
            .in2(N__4778),
            .in3(N__4144),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_9_5  (
            .in0(N__4663),
            .in1(N__4603),
            .in2(N__4165),
            .in3(N__4162),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_10_9_6  (
            .in0(N__4838),
            .in1(N__5103),
            .in2(N__4153),
            .in3(N__4706),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__4449),
            .in2(N__4150),
            .in3(N__4147),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5668));
    defparam RESETn_ibuf_RNIM9SF_LC_10_10_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_10_10_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_10_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_10_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5838),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_0 .LUT_INIT=16'b1111011100000111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_0  (
            .in0(N__4965),
            .in1(N__4991),
            .in2(N__5035),
            .in3(N__5001),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_1 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_1  (
            .in0(N__5133),
            .in1(N__5840),
            .in2(N__4129),
            .in3(N__5008),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_11_2 .LUT_INIT=16'b0000010000110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_11_2  (
            .in0(N__4992),
            .in1(N__5131),
            .in2(N__4969),
            .in3(N__5002),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_11_3 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_11_3  (
            .in0(N__5132),
            .in1(N__5841),
            .in2(N__4126),
            .in3(N__5032),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_11_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_10_11_5  (
            .in0(N__4441),
            .in1(N__4420),
            .in2(N__4402),
            .in3(N__4316),
            .lcout(nBUFEN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_12_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_12_2  (
            .in0(N__4291),
            .in1(N__4261),
            .in2(N__4240),
            .in3(N__4210),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5558));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_6_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_6_0  (
            .in0(N__5236),
            .in1(N__5257),
            .in2(_gnd_net_),
            .in3(N__4858),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_6_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_11_6_1  (
            .in0(N__4189),
            .in1(N__5428),
            .in2(N__4195),
            .in3(N__5275),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_11_6_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_11_6_2  (
            .in0(N__4547),
            .in1(N__4486),
            .in2(N__4192),
            .in3(N__4859),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5317),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_6_3  (
            .in0(N__5334),
            .in1(N__4875),
            .in2(N__5293),
            .in3(N__5413),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_11_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_11_6_4 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_11_6_4  (
            .in0(N__4548),
            .in1(N__5245),
            .in2(N__4522),
            .in3(N__4487),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5317),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_11_6_5  (
            .in0(N__5380),
            .in1(N__5185),
            .in2(N__5161),
            .in3(N__5221),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_11_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_11_6_6  (
            .in0(N__4549),
            .in1(N__4521),
            .in2(N__4582),
            .in3(N__5209),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5317),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_11_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_11_6_7  (
            .in0(N__4860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4876),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5317),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_11_7_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_11_7_0  (
            .in0(N__4514),
            .in1(N__4546),
            .in2(N__5146),
            .in3(N__4484),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5319),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_11_7_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_11_7_1  (
            .in0(N__4544),
            .in1(N__4517),
            .in2(N__4489),
            .in3(N__5347),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5319),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_11_7_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_11_7_2  (
            .in0(N__4513),
            .in1(N__4545),
            .in2(N__5173),
            .in3(N__4483),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5319),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_7_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_11_7_3  (
            .in0(N__5359),
            .in1(N__5443),
            .in2(N__5398),
            .in3(N__5200),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_11_7_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_11_7_4  (
            .in0(N__4515),
            .in1(N__4560),
            .in2(N__4579),
            .in3(N__4485),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5319),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_11_7_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_11_7_7  (
            .in0(N__4543),
            .in1(N__4516),
            .in2(N__4488),
            .in3(N__5368),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5319),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_11_8_2  (
            .in0(N__4686),
            .in1(N__4799),
            .in2(N__4779),
            .in3(N__4735),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__4604),
            .in2(N__4456),
            .in3(N__4664),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_6  (
            .in0(N__4772),
            .in1(N__4800),
            .in2(_gnd_net_),
            .in3(N__4736),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_9_0 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_9_0  (
            .in0(N__4708),
            .in1(N__4839),
            .in2(N__4780),
            .in3(N__5102),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_9_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_9_1  (
            .in0(N__4737),
            .in1(N__4774),
            .in2(_gnd_net_),
            .in3(N__4801),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_9_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_9_2  (
            .in0(N__4773),
            .in1(N__4738),
            .in2(_gnd_net_),
            .in3(N__4625),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_3  (
            .in0(N__4714),
            .in1(N__5458),
            .in2(_gnd_net_),
            .in3(N__4707),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_4  (
            .in0(N__4693),
            .in1(N__4687),
            .in2(_gnd_net_),
            .in3(N__4624),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_5  (
            .in0(N__4623),
            .in1(N__4635),
            .in2(_gnd_net_),
            .in3(N__4666),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_6 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_6  (
            .in0(N__4665),
            .in1(N__4605),
            .in2(N__4639),
            .in3(N__4626),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5664));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_10_3 .LUT_INIT=16'b0100011101000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_10_3  (
            .in0(N__5034),
            .in1(N__5134),
            .in2(N__5044),
            .in3(N__5473),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5548));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_11_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_11_0  (
            .in0(N__5130),
            .in1(N__4900),
            .in2(N__5101),
            .in3(N__4914),
            .lcout(\U409_TRANSFER_ACK.N_107 ),
            .ltout(\U409_TRANSFER_ACK.N_107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_11_1 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_11_1  (
            .in0(N__5033),
            .in1(N__4959),
            .in2(N__5011),
            .in3(N__4990),
            .lcout(\U409_TRANSFER_ACK.m9_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__4899),
            .in2(_gnd_net_),
            .in3(N__4913),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4993),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5559));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_11_12_2  (
            .in0(N__4935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5559));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4915),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5559));
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__4874),
            .in2(N__4861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_12_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__5289),
            .in2(_gnd_net_),
            .in3(N__5278),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__5316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_12_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__5271),
            .in2(_gnd_net_),
            .in3(N__5260),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__5316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__5256),
            .in2(_gnd_net_),
            .in3(N__5239),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_12_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__5235),
            .in2(_gnd_net_),
            .in3(N__5224),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__5316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__5220),
            .in2(_gnd_net_),
            .in3(N__5203),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_12_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_12_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__5199),
            .in2(_gnd_net_),
            .in3(N__5188),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__5316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_12_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__5184),
            .in2(_gnd_net_),
            .in3(N__5164),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_12_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__5157),
            .in2(_gnd_net_),
            .in3(N__5137),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_12_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_12_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__5442),
            .in2(_gnd_net_),
            .in3(N__5431),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__5318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_12_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_12_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__5427),
            .in2(_gnd_net_),
            .in3(N__5416),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__5318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_12_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_12_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__5412),
            .in2(_gnd_net_),
            .in3(N__5401),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__5318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_12_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_12_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__5394),
            .in2(_gnd_net_),
            .in3(N__5383),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__5318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_12_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__5379),
            .in2(_gnd_net_),
            .in3(N__5362),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_12_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__5358),
            .in2(_gnd_net_),
            .in3(N__5341),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_12_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_12_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__5335),
            .in2(_gnd_net_),
            .in3(N__5338),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_8_7 .LUT_INIT=16'b0001000111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_8_7  (
            .in0(N__5612),
            .in1(N__5490),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_9_0 .LUT_INIT=16'b1111010010110100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_9_0  (
            .in0(N__5575),
            .in1(N__5644),
            .in2(N__5494),
            .in3(N__5637),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5560));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_9_5 .LUT_INIT=16'b0010001010001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_9_5  (
            .in0(N__5580),
            .in1(N__5614),
            .in2(N__5638),
            .in3(N__5599),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5560));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_9_6 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_9_6  (
            .in0(N__5598),
            .in1(_gnd_net_),
            .in2(N__5581),
            .in3(N__5633),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5560));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_7  (
            .in0(N__5579),
            .in1(N__5613),
            .in2(_gnd_net_),
            .in3(N__5597),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5560));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_10_0 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_10_0  (
            .in0(N__5925),
            .in1(N__5817),
            .in2(_gnd_net_),
            .in3(N__5937),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_10_1 .LUT_INIT=16'b0000101011101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_12_10_1  (
            .in0(N__5505),
            .in1(N__5926),
            .in2(N__5839),
            .in3(N__5914),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_12_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__5489),
            .in2(_gnd_net_),
            .in3(N__5472),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIURL11_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIURL11_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIURL11_LC_12_10_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIURL11_LC_12_10_4  (
            .in0(N__5924),
            .in1(N__5936),
            .in2(N__5461),
            .in3(N__5457),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5446),
            .in3(N__5792),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_10_7  (
            .in0(N__5938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5793),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_11_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_12_11_5  (
            .in0(N__5804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5913),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__5902),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_13_16_2.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_13_16_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5890),
            .lcout(N_373_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_16_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_16_11_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_16_11_1  (
            .in0(N__5788),
            .in1(N__5706),
            .in2(_gnd_net_),
            .in3(N__5689),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

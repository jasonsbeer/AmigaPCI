-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 8 2025 22:54:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \N_897_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.N_193_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_176_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_253_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_298_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.N_216\ : std_logic;
signal \U712_CHIP_RAM.N_216_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_CHIP_RAM.N_213\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_193\ : std_logic;
signal \U712_CHIP_RAM.N_177_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_223\ : std_logic;
signal \U712_CHIP_RAM.N_300\ : std_logic;
signal \U712_CHIP_RAM.N_223_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_187_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_264_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_262\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_220\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_323\ : std_logic;
signal \U712_CHIP_RAM.N_176\ : std_logic;
signal \U712_CHIP_RAM.N_242_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_319\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.N_177\ : std_logic;
signal \U712_CHIP_RAM.N_319_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_322\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_311\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_46\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_256_i\ : std_logic;
signal \U712_CYCLE_TERM.N_207_i_0_en_cascade_\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_207_i_0_en_0\ : std_logic;
signal \U712_REG_SM.N_185_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.N_197_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_42_1\ : std_logic;
signal \U712_CHIP_RAM.N_236\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_198_i\ : std_logic;
signal \U712_CHIP_RAM.N_187\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_355_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_321\ : std_logic;
signal \U712_CHIP_RAM.N_235\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_217\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_219\ : std_logic;
signal \U712_CHIP_RAM.N_117_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_197\ : std_logic;
signal \U712_REG_SM.N_215_cascade_\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_185\ : std_logic;
signal \U712_REG_SM.N_204_cascade_\ : std_logic;
signal \U712_REG_SM.N_215\ : std_logic;
signal \U712_REG_SM.N_204\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \U712_REG_SM.N_209\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_324_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_242\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0\ : std_logic;
signal \U712_CHIP_RAM.N_253\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_188\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_200\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \un1_LDSn_i_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \un1_UDSn_i_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_212\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.N_298\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_355\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_BYTE_ENABLE.N_275\ : std_logic;
signal \N_148_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_271\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_\ : std_logic;
signal \N_171_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_277\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_\ : std_logic;
signal \N_150_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_270\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_273\ : std_logic;
signal \N_172_i\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CLK40_OUT_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CLK40_OUT <= \CLK40_OUT_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3645\,
            RESETB => \N__6789\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10288\,
            DIN => \N__10287\,
            DOUT => \N__10286\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10288\,
            PADOUT => \N__10287\,
            PADIN => \N__10286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7266\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10279\,
            DIN => \N__10278\,
            DOUT => \N__10277\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10279\,
            PADOUT => \N__10278\,
            PADIN => \N__10277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10270\,
            DIN => \N__10269\,
            DOUT => \N__10268\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10270\,
            PADOUT => \N__10269\,
            PADIN => \N__10268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8742\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10261\,
            DIN => \N__10260\,
            DOUT => \N__10259\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10261\,
            PADOUT => \N__10260\,
            PADIN => \N__10259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10252\,
            DIN => \N__10251\,
            DOUT => \N__10250\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10252\,
            PADOUT => \N__10251\,
            PADIN => \N__10250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10243\,
            DIN => \N__10242\,
            DOUT => \N__10241\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10243\,
            PADOUT => \N__10242\,
            PADIN => \N__10241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10234\,
            DIN => \N__10233\,
            DOUT => \N__10232\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10234\,
            PADOUT => \N__10233\,
            PADIN => \N__10232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10225\,
            DIN => \N__10224\,
            DOUT => \N__10223\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10225\,
            PADOUT => \N__10224\,
            PADIN => \N__10223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10216\,
            DIN => \N__10215\,
            DOUT => \N__10214\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10216\,
            PADOUT => \N__10215\,
            PADIN => \N__10214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10207\,
            DIN => \N__10206\,
            DOUT => \N__10205\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10207\,
            PADOUT => \N__10206\,
            PADIN => \N__10205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10198\,
            DIN => \N__10197\,
            DOUT => \N__10196\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10198\,
            PADOUT => \N__10197\,
            PADIN => \N__10196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10189\,
            DIN => \N__10188\,
            DOUT => \N__10187\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10189\,
            PADOUT => \N__10188\,
            PADIN => \N__10187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10180\,
            DIN => \N__10179\,
            DOUT => \N__10178\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10180\,
            PADOUT => \N__10179\,
            PADIN => \N__10178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10171\,
            DIN => \N__10170\,
            DOUT => \N__10169\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10171\,
            PADOUT => \N__10170\,
            PADIN => \N__10169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10162\,
            DIN => \N__10161\,
            DOUT => \N__10160\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10162\,
            PADOUT => \N__10161\,
            PADIN => \N__10160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10153\,
            DIN => \N__10152\,
            DOUT => \N__10151\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10153\,
            PADOUT => \N__10152\,
            PADIN => \N__10151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10144\,
            DIN => \N__10143\,
            DOUT => \N__10142\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10144\,
            PADOUT => \N__10143\,
            PADIN => \N__10142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10135\,
            DIN => \N__10134\,
            DOUT => \N__10133\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10135\,
            PADOUT => \N__10134\,
            PADIN => \N__10133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10126\,
            DIN => \N__10125\,
            DOUT => \N__10124\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10126\,
            PADOUT => \N__10125\,
            PADIN => \N__10124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10117\,
            DIN => \N__10116\,
            DOUT => \N__10115\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10117\,
            PADOUT => \N__10116\,
            PADIN => \N__10115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8676\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10108\,
            DIN => \N__10107\,
            DOUT => \N__10106\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10108\,
            PADOUT => \N__10107\,
            PADIN => \N__10106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10099\,
            DIN => \N__10098\,
            DOUT => \N__10097\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10099\,
            PADOUT => \N__10098\,
            PADIN => \N__10097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10090\,
            DIN => \N__10089\,
            DOUT => \N__10088\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10090\,
            PADOUT => \N__10089\,
            PADIN => \N__10088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10081\,
            DIN => \N__10080\,
            DOUT => \N__10079\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10081\,
            PADOUT => \N__10080\,
            PADIN => \N__10079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10072\,
            DIN => \N__10071\,
            DOUT => \N__10070\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10072\,
            PADOUT => \N__10071\,
            PADIN => \N__10070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10063\,
            DIN => \N__10062\,
            DOUT => \N__10061\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10063\,
            PADOUT => \N__10062\,
            PADIN => \N__10061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10054\,
            DIN => \N__10053\,
            DOUT => \N__10052\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10054\,
            PADOUT => \N__10053\,
            PADIN => \N__10052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10045\,
            DIN => \N__10044\,
            DOUT => \N__10043\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10045\,
            PADOUT => \N__10044\,
            PADIN => \N__10043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10036\,
            DIN => \N__10035\,
            DOUT => \N__10034\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10036\,
            PADOUT => \N__10035\,
            PADIN => \N__10034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10027\,
            DIN => \N__10026\,
            DOUT => \N__10025\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10027\,
            PADOUT => \N__10026\,
            PADIN => \N__10025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10018\,
            DIN => \N__10017\,
            DOUT => \N__10016\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10018\,
            PADOUT => \N__10017\,
            PADIN => \N__10016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10009\,
            DIN => \N__10008\,
            DOUT => \N__10007\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10009\,
            PADOUT => \N__10008\,
            PADIN => \N__10007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10000\,
            DIN => \N__9999\,
            DOUT => \N__9998\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10000\,
            PADOUT => \N__9999\,
            PADIN => \N__9998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9991\,
            DIN => \N__9990\,
            DOUT => \N__9989\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9991\,
            PADOUT => \N__9990\,
            PADIN => \N__9989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9982\,
            DIN => \N__9981\,
            DOUT => \N__9980\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9982\,
            PADOUT => \N__9981\,
            PADIN => \N__9980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9973\,
            DIN => \N__9972\,
            DOUT => \N__9971\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9973\,
            PADOUT => \N__9972\,
            PADIN => \N__9971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9964\,
            DIN => \N__9963\,
            DOUT => \N__9962\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9964\,
            PADOUT => \N__9963\,
            PADIN => \N__9962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6162\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9955\,
            DIN => \N__9954\,
            DOUT => \N__9953\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9955\,
            PADOUT => \N__9954\,
            PADIN => \N__9953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9946\,
            DIN => \N__9945\,
            DOUT => \N__9944\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9946\,
            PADOUT => \N__9945\,
            PADIN => \N__9944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7641\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9937\,
            DIN => \N__9936\,
            DOUT => \N__9935\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9937\,
            PADOUT => \N__9936\,
            PADIN => \N__9935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9928\,
            DIN => \N__9927\,
            DOUT => \N__9926\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9928\,
            PADOUT => \N__9927\,
            PADIN => \N__9926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9919\,
            DIN => \N__9918\,
            DOUT => \N__9917\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9919\,
            PADOUT => \N__9918\,
            PADIN => \N__9917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3663\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9910\,
            DIN => \N__9909\,
            DOUT => \N__9908\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9910\,
            PADOUT => \N__9909\,
            PADIN => \N__9908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4998\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9901\,
            DIN => \N__9900\,
            DOUT => \N__9899\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9901\,
            PADOUT => \N__9900\,
            PADIN => \N__9899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7575\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9892\,
            DIN => \N__9891\,
            DOUT => \N__9890\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9892\,
            PADOUT => \N__9891\,
            PADIN => \N__9890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9883\,
            DIN => \N__9882\,
            DOUT => \N__9881\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9883\,
            PADOUT => \N__9882\,
            PADIN => \N__9881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9874\,
            DIN => \N__9873\,
            DOUT => \N__9872\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9874\,
            PADOUT => \N__9873\,
            PADIN => \N__9872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9865\,
            DIN => \N__9864\,
            DOUT => \N__9863\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9865\,
            PADOUT => \N__9864\,
            PADIN => \N__9863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5130\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9856\,
            DIN => \N__9855\,
            DOUT => \N__9854\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9856\,
            PADOUT => \N__9855\,
            PADIN => \N__9854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9847\,
            DIN => \N__9846\,
            DOUT => \N__9845\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9847\,
            PADOUT => \N__9846\,
            PADIN => \N__9845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8610\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9838\,
            DIN => \N__9837\,
            DOUT => \N__9836\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9838\,
            PADOUT => \N__9837\,
            PADIN => \N__9836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9829\,
            DIN => \N__9828\,
            DOUT => \N__9827\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9829\,
            PADOUT => \N__9828\,
            PADIN => \N__9827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7170\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9820\,
            DIN => \N__9819\,
            DOUT => \N__9818\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9820\,
            PADOUT => \N__9819\,
            PADIN => \N__9818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7392\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9811\,
            DIN => \N__9810\,
            DOUT => \N__9809\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9811\,
            PADOUT => \N__9810\,
            PADIN => \N__9809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9802\,
            DIN => \N__9801\,
            DOUT => \N__9800\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9802\,
            PADOUT => \N__9801\,
            PADIN => \N__9800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9793\,
            DIN => \N__9792\,
            DOUT => \N__9791\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9793\,
            PADOUT => \N__9792\,
            PADIN => \N__9791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9784\,
            DIN => \N__9783\,
            DOUT => \N__9782\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9784\,
            PADOUT => \N__9783\,
            PADIN => \N__9782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9775\,
            DIN => \N__9774\,
            DOUT => \N__9773\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9775\,
            PADOUT => \N__9774\,
            PADIN => \N__9773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9766\,
            DIN => \N__9765\,
            DOUT => \N__9764\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9766\,
            PADOUT => \N__9765\,
            PADIN => \N__9764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6681\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9757\,
            DIN => \N__9756\,
            DOUT => \N__9755\,
            PACKAGEPIN => \CLK40_OUT_wire\
        );

    \CLK40_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9757\,
            PADOUT => \N__9756\,
            PADIN => \N__9755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9748\,
            DIN => \N__9747\,
            DOUT => \N__9746\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9748\,
            PADOUT => \N__9747\,
            PADIN => \N__9746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7116\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9739\,
            DIN => \N__9738\,
            DOUT => \N__9737\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9739\,
            PADOUT => \N__9738\,
            PADIN => \N__9737\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9730\,
            DIN => \N__9729\,
            DOUT => \N__9728\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9730\,
            PADOUT => \N__9729\,
            PADIN => \N__9728\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9721\,
            DIN => \N__9720\,
            DOUT => \N__9719\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9721\,
            PADOUT => \N__9720\,
            PADIN => \N__9719\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9712\,
            DIN => \N__9711\,
            DOUT => \N__9710\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9712\,
            PADOUT => \N__9711\,
            PADIN => \N__9710\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9703\,
            DIN => \N__9702\,
            DOUT => \N__9701\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9703\,
            PADOUT => \N__9702\,
            PADIN => \N__9701\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5772\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9694\,
            DIN => \N__9693\,
            DOUT => \N__9692\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9694\,
            PADOUT => \N__9693\,
            PADIN => \N__9692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9685\,
            DIN => \N__9684\,
            DOUT => \N__9683\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9685\,
            PADOUT => \N__9684\,
            PADIN => \N__9683\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9676\,
            DIN => \N__9675\,
            DOUT => \N__9674\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9676\,
            PADOUT => \N__9675\,
            PADIN => \N__9674\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3678\,
            DIN0 => OPEN,
            DOUT0 => \N__6357\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9667\,
            DIN => \N__9666\,
            DOUT => \N__9665\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9667\,
            PADOUT => \N__9666\,
            PADIN => \N__9665\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9658\,
            DIN => \N__9657\,
            DOUT => \N__9656\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9658\,
            PADOUT => \N__9657\,
            PADIN => \N__9656\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9649\,
            DIN => \N__9648\,
            DOUT => \N__9647\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9649\,
            PADOUT => \N__9648\,
            PADIN => \N__9647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9640\,
            DIN => \N__9639\,
            DOUT => \N__9638\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9640\,
            PADOUT => \N__9639\,
            PADIN => \N__9638\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9631\,
            DIN => \N__9630\,
            DOUT => \N__9629\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9631\,
            PADOUT => \N__9630\,
            PADIN => \N__9629\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9622\,
            DIN => \N__9621\,
            DOUT => \N__9620\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9622\,
            PADOUT => \N__9621\,
            PADIN => \N__9620\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9613\,
            DIN => \N__9612\,
            DOUT => \N__9611\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9613\,
            PADOUT => \N__9612\,
            PADIN => \N__9611\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9604\,
            DIN => \N__9603\,
            DOUT => \N__9602\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9604\,
            PADOUT => \N__9603\,
            PADIN => \N__9602\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9595\,
            DIN => \N__9594\,
            DOUT => \N__9593\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9595\,
            PADOUT => \N__9594\,
            PADIN => \N__9593\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5742\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9586\,
            DIN => \N__9585\,
            DOUT => \N__9584\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9586\,
            PADOUT => \N__9585\,
            PADIN => \N__9584\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2291\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__9558\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9552\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9552\,
            I => \N__9548\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9545\
        );

    \I__2284\ : Span4Mux_v
    port map (
            O => \N__9548\,
            I => \N__9542\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9539\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__9542\,
            I => \N__9536\
        );

    \I__2281\ : Sp12to4
    port map (
            O => \N__9539\,
            I => \N__9533\
        );

    \I__2280\ : Sp12to4
    port map (
            O => \N__9536\,
            I => \N__9528\
        );

    \I__2279\ : Span12Mux_v
    port map (
            O => \N__9533\,
            I => \N__9528\
        );

    \I__2278\ : Span12Mux_h
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2277\ : Odrv12
    port map (
            O => \N__9525\,
            I => \DRA_c_7\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9516\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__9513\,
            I => \N__9510\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__9510\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2271\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__9504\,
            I => \N__9495\
        );

    \I__2269\ : ClkMux
    port map (
            O => \N__9503\,
            I => \N__9480\
        );

    \I__2268\ : ClkMux
    port map (
            O => \N__9502\,
            I => \N__9480\
        );

    \I__2267\ : ClkMux
    port map (
            O => \N__9501\,
            I => \N__9480\
        );

    \I__2266\ : ClkMux
    port map (
            O => \N__9500\,
            I => \N__9480\
        );

    \I__2265\ : ClkMux
    port map (
            O => \N__9499\,
            I => \N__9480\
        );

    \I__2264\ : ClkMux
    port map (
            O => \N__9498\,
            I => \N__9480\
        );

    \I__2263\ : Glb2LocalMux
    port map (
            O => \N__9495\,
            I => \N__9480\
        );

    \I__2262\ : GlobalMux
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2261\ : gio2CtrlBuf
    port map (
            O => \N__9477\,
            I => \C3_c_g\
        );

    \I__2260\ : CEMux
    port map (
            O => \N__9474\,
            I => \N__9471\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9471\,
            I => \N__9464\
        );

    \I__2258\ : CEMux
    port map (
            O => \N__9470\,
            I => \N__9461\
        );

    \I__2257\ : CEMux
    port map (
            O => \N__9469\,
            I => \N__9458\
        );

    \I__2256\ : CEMux
    port map (
            O => \N__9468\,
            I => \N__9455\
        );

    \I__2255\ : CEMux
    port map (
            O => \N__9467\,
            I => \N__9452\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__9464\,
            I => \N__9446\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9446\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9443\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9438\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__9452\,
            I => \N__9438\
        );

    \I__2249\ : CEMux
    port map (
            O => \N__9451\,
            I => \N__9435\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__9446\,
            I => \N__9430\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__9443\,
            I => \N__9430\
        );

    \I__2246\ : Span4Mux_v
    port map (
            O => \N__9438\,
            I => \N__9427\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9435\,
            I => \N__9424\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9430\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__9427\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2242\ : Odrv12
    port map (
            O => \N__9424\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9409\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9406\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9403\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9400\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9397\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9394\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9409\,
            I => \N__9388\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9382\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9372\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9360\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9397\,
            I => \N__9351\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N__9342\
        );

    \I__2229\ : SRMux
    port map (
            O => \N__9393\,
            I => \N__9246\
        );

    \I__2228\ : SRMux
    port map (
            O => \N__9392\,
            I => \N__9246\
        );

    \I__2227\ : SRMux
    port map (
            O => \N__9391\,
            I => \N__9246\
        );

    \I__2226\ : Glb2LocalMux
    port map (
            O => \N__9388\,
            I => \N__9246\
        );

    \I__2225\ : SRMux
    port map (
            O => \N__9387\,
            I => \N__9246\
        );

    \I__2224\ : SRMux
    port map (
            O => \N__9386\,
            I => \N__9246\
        );

    \I__2223\ : SRMux
    port map (
            O => \N__9385\,
            I => \N__9246\
        );

    \I__2222\ : Glb2LocalMux
    port map (
            O => \N__9382\,
            I => \N__9246\
        );

    \I__2221\ : SRMux
    port map (
            O => \N__9381\,
            I => \N__9246\
        );

    \I__2220\ : SRMux
    port map (
            O => \N__9380\,
            I => \N__9246\
        );

    \I__2219\ : SRMux
    port map (
            O => \N__9379\,
            I => \N__9246\
        );

    \I__2218\ : SRMux
    port map (
            O => \N__9378\,
            I => \N__9246\
        );

    \I__2217\ : SRMux
    port map (
            O => \N__9377\,
            I => \N__9246\
        );

    \I__2216\ : SRMux
    port map (
            O => \N__9376\,
            I => \N__9246\
        );

    \I__2215\ : SRMux
    port map (
            O => \N__9375\,
            I => \N__9246\
        );

    \I__2214\ : Glb2LocalMux
    port map (
            O => \N__9372\,
            I => \N__9246\
        );

    \I__2213\ : SRMux
    port map (
            O => \N__9371\,
            I => \N__9246\
        );

    \I__2212\ : SRMux
    port map (
            O => \N__9370\,
            I => \N__9246\
        );

    \I__2211\ : SRMux
    port map (
            O => \N__9369\,
            I => \N__9246\
        );

    \I__2210\ : SRMux
    port map (
            O => \N__9368\,
            I => \N__9246\
        );

    \I__2209\ : SRMux
    port map (
            O => \N__9367\,
            I => \N__9246\
        );

    \I__2208\ : SRMux
    port map (
            O => \N__9366\,
            I => \N__9246\
        );

    \I__2207\ : SRMux
    port map (
            O => \N__9365\,
            I => \N__9246\
        );

    \I__2206\ : SRMux
    port map (
            O => \N__9364\,
            I => \N__9246\
        );

    \I__2205\ : SRMux
    port map (
            O => \N__9363\,
            I => \N__9246\
        );

    \I__2204\ : Glb2LocalMux
    port map (
            O => \N__9360\,
            I => \N__9246\
        );

    \I__2203\ : SRMux
    port map (
            O => \N__9359\,
            I => \N__9246\
        );

    \I__2202\ : SRMux
    port map (
            O => \N__9358\,
            I => \N__9246\
        );

    \I__2201\ : SRMux
    port map (
            O => \N__9357\,
            I => \N__9246\
        );

    \I__2200\ : SRMux
    port map (
            O => \N__9356\,
            I => \N__9246\
        );

    \I__2199\ : SRMux
    port map (
            O => \N__9355\,
            I => \N__9246\
        );

    \I__2198\ : SRMux
    port map (
            O => \N__9354\,
            I => \N__9246\
        );

    \I__2197\ : Glb2LocalMux
    port map (
            O => \N__9351\,
            I => \N__9246\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9350\,
            I => \N__9246\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9349\,
            I => \N__9246\
        );

    \I__2194\ : SRMux
    port map (
            O => \N__9348\,
            I => \N__9246\
        );

    \I__2193\ : SRMux
    port map (
            O => \N__9347\,
            I => \N__9246\
        );

    \I__2192\ : SRMux
    port map (
            O => \N__9346\,
            I => \N__9246\
        );

    \I__2191\ : SRMux
    port map (
            O => \N__9345\,
            I => \N__9246\
        );

    \I__2190\ : Glb2LocalMux
    port map (
            O => \N__9342\,
            I => \N__9246\
        );

    \I__2189\ : SRMux
    port map (
            O => \N__9341\,
            I => \N__9246\
        );

    \I__2188\ : SRMux
    port map (
            O => \N__9340\,
            I => \N__9246\
        );

    \I__2187\ : SRMux
    port map (
            O => \N__9339\,
            I => \N__9246\
        );

    \I__2186\ : SRMux
    port map (
            O => \N__9338\,
            I => \N__9246\
        );

    \I__2185\ : SRMux
    port map (
            O => \N__9337\,
            I => \N__9246\
        );

    \I__2184\ : GlobalMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__2183\ : gio2CtrlBuf
    port map (
            O => \N__9243\,
            I => \RESETn_c_i_g\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__9234\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__9216\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9209\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9206\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9209\,
            I => \N__9203\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9206\,
            I => \N__9200\
        );

    \I__2169\ : Span4Mux_h
    port map (
            O => \N__9203\,
            I => \N__9197\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__9200\,
            I => \N__9194\
        );

    \I__2167\ : Sp12to4
    port map (
            O => \N__9197\,
            I => \N__9191\
        );

    \I__2166\ : Sp12to4
    port map (
            O => \N__9194\,
            I => \N__9188\
        );

    \I__2165\ : Span12Mux_v
    port map (
            O => \N__9191\,
            I => \N__9185\
        );

    \I__2164\ : Span12Mux_h
    port map (
            O => \N__9188\,
            I => \N__9182\
        );

    \I__2163\ : Span12Mux_h
    port map (
            O => \N__9185\,
            I => \N__9177\
        );

    \I__2162\ : Span12Mux_v
    port map (
            O => \N__9182\,
            I => \N__9177\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__9177\,
            I => \DRA_c_4\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__9165\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__2154\ : Span4Mux_h
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__9153\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9146\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9146\,
            I => \N__9138\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9143\,
            I => \N__9138\
        );

    \I__2148\ : Span12Mux_v
    port map (
            O => \N__9138\,
            I => \N__9135\
        );

    \I__2147\ : Span12Mux_h
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__2146\ : Span12Mux_v
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__9129\,
            I => \DRA_c_9\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__9120\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9113\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9110\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9105\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9105\
        );

    \I__2137\ : Span12Mux_v
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__2136\ : Span12Mux_h
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__2135\ : Span12Mux_v
    port map (
            O => \N__9099\,
            I => \N__9096\
        );

    \I__2134\ : Odrv12
    port map (
            O => \N__9096\,
            I => \DRA_c_1\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__2131\ : Odrv12
    port map (
            O => \N__9087\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2130\ : CEMux
    port map (
            O => \N__9084\,
            I => \N__9078\
        );

    \I__2129\ : CEMux
    port map (
            O => \N__9083\,
            I => \N__9075\
        );

    \I__2128\ : CEMux
    port map (
            O => \N__9082\,
            I => \N__9072\
        );

    \I__2127\ : CEMux
    port map (
            O => \N__9081\,
            I => \N__9069\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9066\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9075\,
            I => \N__9062\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9072\,
            I => \N__9059\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9056\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__9066\,
            I => \N__9053\
        );

    \I__2121\ : CEMux
    port map (
            O => \N__9065\,
            I => \N__9050\
        );

    \I__2120\ : Span4Mux_h
    port map (
            O => \N__9062\,
            I => \N__9047\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__9059\,
            I => \N__9038\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9056\,
            I => \N__9038\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__9053\,
            I => \N__9038\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__9038\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__9047\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__9038\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9033\,
            I => \N__9029\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9026\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__9021\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9021\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__9021\,
            I => \N__9018\
        );

    \I__2108\ : Sp12to4
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__2107\ : Span12Mux_v
    port map (
            O => \N__9015\,
            I => \N__9012\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__9012\,
            I => \DRA_c_5\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__9003\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8993\
        );

    \I__2100\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8990\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__8993\,
            I => \N__8985\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8985\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__2096\ : Span4Mux_v
    port map (
            O => \N__8982\,
            I => \N__8979\
        );

    \I__2095\ : Sp12to4
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__8976\,
            I => \DRA_c_8\
        );

    \I__2093\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8970\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__8967\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2090\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__8961\,
            I => \N__8958\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__8955\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2086\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8945\
        );

    \I__2084\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8942\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8939\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8936\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__8939\,
            I => \N__8933\
        );

    \I__2080\ : Span12Mux_h
    port map (
            O => \N__8936\,
            I => \N__8930\
        );

    \I__2079\ : Span12Mux_h
    port map (
            O => \N__8933\,
            I => \N__8927\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__8930\,
            I => \RAS0n_c\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__8927\,
            I => \RAS0n_c\
        );

    \I__2076\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__8919\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8913\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__8913\,
            I => \N__8909\
        );

    \I__2072\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8906\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__8909\,
            I => \N__8901\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8906\,
            I => \N__8901\
        );

    \I__2069\ : Sp12to4
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__2068\ : Span12Mux_v
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__2067\ : Span12Mux_h
    port map (
            O => \N__8895\,
            I => \N__8892\
        );

    \I__2066\ : Odrv12
    port map (
            O => \N__8892\,
            I => \DRA_c_6\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8883\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8883\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8880\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__8877\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2060\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__2058\ : ClkMux
    port map (
            O => \N__8870\,
            I => \N__8847\
        );

    \I__2057\ : ClkMux
    port map (
            O => \N__8869\,
            I => \N__8847\
        );

    \I__2056\ : ClkMux
    port map (
            O => \N__8868\,
            I => \N__8847\
        );

    \I__2055\ : ClkMux
    port map (
            O => \N__8867\,
            I => \N__8847\
        );

    \I__2054\ : ClkMux
    port map (
            O => \N__8866\,
            I => \N__8847\
        );

    \I__2053\ : ClkMux
    port map (
            O => \N__8865\,
            I => \N__8847\
        );

    \I__2052\ : Glb2LocalMux
    port map (
            O => \N__8862\,
            I => \N__8847\
        );

    \I__2051\ : GlobalMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__2050\ : gio2CtrlBuf
    port map (
            O => \N__8844\,
            I => \C1_c_g\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8837\
        );

    \I__2048\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8833\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8830\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8827\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8824\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__8830\,
            I => \N__8819\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8827\,
            I => \N__8819\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__8824\,
            I => \N__8816\
        );

    \I__2041\ : Sp12to4
    port map (
            O => \N__8819\,
            I => \N__8813\
        );

    \I__2040\ : Sp12to4
    port map (
            O => \N__8816\,
            I => \N__8810\
        );

    \I__2039\ : Span12Mux_v
    port map (
            O => \N__8813\,
            I => \N__8807\
        );

    \I__2038\ : Span12Mux_h
    port map (
            O => \N__8810\,
            I => \N__8804\
        );

    \I__2037\ : Span12Mux_h
    port map (
            O => \N__8807\,
            I => \N__8801\
        );

    \I__2036\ : Span12Mux_v
    port map (
            O => \N__8804\,
            I => \N__8798\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__8801\,
            I => \DBRn_c\
        );

    \I__2034\ : Odrv12
    port map (
            O => \N__8798\,
            I => \DBRn_c\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8790\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2031\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__8781\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8774\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8771\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8768\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8765\
        );

    \I__2024\ : Span12Mux_h
    port map (
            O => \N__8768\,
            I => \N__8762\
        );

    \I__2023\ : Span12Mux_v
    port map (
            O => \N__8765\,
            I => \N__8759\
        );

    \I__2022\ : Span12Mux_v
    port map (
            O => \N__8762\,
            I => \N__8754\
        );

    \I__2021\ : Span12Mux_h
    port map (
            O => \N__8759\,
            I => \N__8754\
        );

    \I__2020\ : Odrv12
    port map (
            O => \N__8754\,
            I => \DRA_c_3\
        );

    \I__2019\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__2017\ : Odrv12
    port map (
            O => \N__8745\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2016\ : IoInMux
    port map (
            O => \N__8742\,
            I => \N__8739\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__2014\ : Span4Mux_s2_v
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__8724\,
            I => \CASn_c\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8715\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__8720\,
            I => \N__8712\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__8719\,
            I => \N__8709\
        );

    \I__2006\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8706\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8703\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8699\
        );

    \I__2003\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8696\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__8706\,
            I => \N__8691\
        );

    \I__2001\ : Span4Mux_h
    port map (
            O => \N__8703\,
            I => \N__8691\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8688\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8685\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8696\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__8691\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8688\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__8685\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1994\ : IoInMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1992\ : Span4Mux_s2_v
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__8661\,
            I => \CRCSn_c\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8655\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1984\ : Span4Mux_s3_v
    port map (
            O => \N__8646\,
            I => \N__8643\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__8640\,
            I => \CMA_c_0\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8631\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8631\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__8625\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8619\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__8613\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1972\ : IoInMux
    port map (
            O => \N__8610\,
            I => \N__8607\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1970\ : IoSpan4Mux
    port map (
            O => \N__8604\,
            I => \N__8601\
        );

    \I__1969\ : Sp12to4
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__1968\ : Span12Mux_s7_v
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__1967\ : Span12Mux_h
    port map (
            O => \N__8595\,
            I => \N__8592\
        );

    \I__1966\ : Odrv12
    port map (
            O => \N__8592\,
            I => \CMA_c_4\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__8589\,
            I => \N__8585\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__8588\,
            I => \N__8580\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8573\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__8584\,
            I => \N__8566\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__8583\,
            I => \N__8563\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8559\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8556\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__8578\,
            I => \N__8553\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__8577\,
            I => \N__8549\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__8576\,
            I => \N__8545\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8540\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8535\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8532\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8521\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8521\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8521\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8521\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8518\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8512\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8512\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8509\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8506\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8497\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8497\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8497\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8497\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8493\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8490\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8487\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8484\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8481\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8478\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8473\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8473\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8468\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8468\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8465\
        );

    \I__1928\ : Span4Mux_h
    port map (
            O => \N__8512\,
            I => \N__8456\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8456\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8456\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8456\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8453\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8444\
        );

    \I__1922\ : Sp12to4
    port map (
            O => \N__8490\,
            I => \N__8444\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8444\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8444\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__8481\,
            I => \N__8437\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__8478\,
            I => \N__8437\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8473\,
            I => \N__8437\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__8468\,
            I => \N__8432\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8432\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__8456\,
            I => \N__8429\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8424\
        );

    \I__1912\ : Span12Mux_h
    port map (
            O => \N__8444\,
            I => \N__8424\
        );

    \I__1911\ : Span4Mux_h
    port map (
            O => \N__8437\,
            I => \N__8421\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__8432\,
            I => \CPU_CYCLEm\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__8429\,
            I => \CPU_CYCLEm\
        );

    \I__1908\ : Odrv12
    port map (
            O => \N__8424\,
            I => \CPU_CYCLEm\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__8421\,
            I => \CPU_CYCLEm\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__8406\,
            I => \N__8403\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__8403\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__8400\,
            I => \N__8395\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8390\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__8398\,
            I => \N__8387\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8382\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8379\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__8393\,
            I => \N__8376\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8373\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8370\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8365\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8365\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8361\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8353\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8350\
        );

    \I__1889\ : Span4Mux_h
    port map (
            O => \N__8373\,
            I => \N__8343\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8343\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8343\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__8364\,
            I => \N__8331\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__8361\,
            I => \N__8327\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8318\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8318\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8318\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8318\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8315\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__8353\,
            I => \N__8312\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8307\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__8343\,
            I => \N__8307\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8302\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8302\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8291\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8291\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8291\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8291\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8291\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8282\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8282\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8282\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8282\
        );

    \I__1865\ : Sp12to4
    port map (
            O => \N__8327\,
            I => \N__8275\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8318\,
            I => \N__8275\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8275\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__8312\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__8307\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8302\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8291\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8282\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__8275\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__8262\,
            I => \N__8259\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8253\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__8258\,
            I => \N__8249\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__8257\,
            I => \N__8246\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__8256\,
            I => \N__8242\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8253\,
            I => \N__8239\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8234\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8234\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8231\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8226\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8226\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__8239\,
            I => \N__8219\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8219\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8214\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8214\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__8225\,
            I => \N__8211\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8207\
        );

    \I__1839\ : Span4Mux_h
    port map (
            O => \N__8219\,
            I => \N__8204\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__8214\,
            I => \N__8201\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8196\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8196\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8207\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__8204\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__8201\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8196\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8179\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8176\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8173\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8170\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8167\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8164\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8179\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8176\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8173\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8170\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8167\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8164\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__8151\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\
        );

    \I__1818\ : IoInMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8142\
        );

    \I__1816\ : IoSpan4Mux
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1815\ : Span4Mux_s2_h
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1813\ : Span12Mux_h
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__8130\,
            I => \CMA_c_7\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8124\,
            I => \N__8096\
        );

    \I__1809\ : ClkMux
    port map (
            O => \N__8123\,
            I => \N__8019\
        );

    \I__1808\ : ClkMux
    port map (
            O => \N__8122\,
            I => \N__8019\
        );

    \I__1807\ : ClkMux
    port map (
            O => \N__8121\,
            I => \N__8019\
        );

    \I__1806\ : ClkMux
    port map (
            O => \N__8120\,
            I => \N__8019\
        );

    \I__1805\ : ClkMux
    port map (
            O => \N__8119\,
            I => \N__8019\
        );

    \I__1804\ : ClkMux
    port map (
            O => \N__8118\,
            I => \N__8019\
        );

    \I__1803\ : ClkMux
    port map (
            O => \N__8117\,
            I => \N__8019\
        );

    \I__1802\ : ClkMux
    port map (
            O => \N__8116\,
            I => \N__8019\
        );

    \I__1801\ : ClkMux
    port map (
            O => \N__8115\,
            I => \N__8019\
        );

    \I__1800\ : ClkMux
    port map (
            O => \N__8114\,
            I => \N__8019\
        );

    \I__1799\ : ClkMux
    port map (
            O => \N__8113\,
            I => \N__8019\
        );

    \I__1798\ : ClkMux
    port map (
            O => \N__8112\,
            I => \N__8019\
        );

    \I__1797\ : ClkMux
    port map (
            O => \N__8111\,
            I => \N__8019\
        );

    \I__1796\ : ClkMux
    port map (
            O => \N__8110\,
            I => \N__8019\
        );

    \I__1795\ : ClkMux
    port map (
            O => \N__8109\,
            I => \N__8019\
        );

    \I__1794\ : ClkMux
    port map (
            O => \N__8108\,
            I => \N__8019\
        );

    \I__1793\ : ClkMux
    port map (
            O => \N__8107\,
            I => \N__8019\
        );

    \I__1792\ : ClkMux
    port map (
            O => \N__8106\,
            I => \N__8019\
        );

    \I__1791\ : ClkMux
    port map (
            O => \N__8105\,
            I => \N__8019\
        );

    \I__1790\ : ClkMux
    port map (
            O => \N__8104\,
            I => \N__8019\
        );

    \I__1789\ : ClkMux
    port map (
            O => \N__8103\,
            I => \N__8019\
        );

    \I__1788\ : ClkMux
    port map (
            O => \N__8102\,
            I => \N__8019\
        );

    \I__1787\ : ClkMux
    port map (
            O => \N__8101\,
            I => \N__8019\
        );

    \I__1786\ : ClkMux
    port map (
            O => \N__8100\,
            I => \N__8019\
        );

    \I__1785\ : ClkMux
    port map (
            O => \N__8099\,
            I => \N__8019\
        );

    \I__1784\ : Glb2LocalMux
    port map (
            O => \N__8096\,
            I => \N__8019\
        );

    \I__1783\ : ClkMux
    port map (
            O => \N__8095\,
            I => \N__8019\
        );

    \I__1782\ : ClkMux
    port map (
            O => \N__8094\,
            I => \N__8019\
        );

    \I__1781\ : ClkMux
    port map (
            O => \N__8093\,
            I => \N__8019\
        );

    \I__1780\ : ClkMux
    port map (
            O => \N__8092\,
            I => \N__8019\
        );

    \I__1779\ : ClkMux
    port map (
            O => \N__8091\,
            I => \N__8019\
        );

    \I__1778\ : ClkMux
    port map (
            O => \N__8090\,
            I => \N__8019\
        );

    \I__1777\ : ClkMux
    port map (
            O => \N__8089\,
            I => \N__8019\
        );

    \I__1776\ : ClkMux
    port map (
            O => \N__8088\,
            I => \N__8019\
        );

    \I__1775\ : GlobalMux
    port map (
            O => \N__8019\,
            I => \CLK80_PLL\
        );

    \I__1774\ : CEMux
    port map (
            O => \N__8016\,
            I => \N__8012\
        );

    \I__1773\ : CEMux
    port map (
            O => \N__8015\,
            I => \N__8009\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8012\,
            I => \N__8004\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__8001\
        );

    \I__1770\ : CEMux
    port map (
            O => \N__8008\,
            I => \N__7997\
        );

    \I__1769\ : CEMux
    port map (
            O => \N__8007\,
            I => \N__7994\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__8004\,
            I => \N__7989\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__8001\,
            I => \N__7989\
        );

    \I__1766\ : CEMux
    port map (
            O => \N__8000\,
            I => \N__7986\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7997\,
            I => \N__7981\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7994\,
            I => \N__7978\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__7989\,
            I => \N__7973\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7973\
        );

    \I__1761\ : CEMux
    port map (
            O => \N__7985\,
            I => \N__7970\
        );

    \I__1760\ : CEMux
    port map (
            O => \N__7984\,
            I => \N__7967\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__7981\,
            I => \N__7964\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__7978\,
            I => \N__7959\
        );

    \I__1757\ : Span4Mux_h
    port map (
            O => \N__7973\,
            I => \N__7959\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7954\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7967\,
            I => \N__7954\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__7964\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__7959\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__7954\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__7941\,
            I => \N__7937\
        );

    \I__1748\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7934\
        );

    \I__1747\ : Sp12to4
    port map (
            O => \N__7937\,
            I => \N__7931\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7934\,
            I => \N__7928\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__7931\,
            I => \N__7925\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__7928\,
            I => \N__7922\
        );

    \I__1743\ : Span12Mux_v
    port map (
            O => \N__7925\,
            I => \N__7919\
        );

    \I__1742\ : Span12Mux_v
    port map (
            O => \N__7922\,
            I => \N__7916\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__7919\,
            I => \DRA_c_2\
        );

    \I__1740\ : Odrv12
    port map (
            O => \N__7916\,
            I => \DRA_c_2\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7908\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__7905\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7898\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7895\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7898\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7895\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7890\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7883\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7880\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7877\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7880\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__7877\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7872\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__7869\,
            I => \N__7865\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7862\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7859\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7862\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7859\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1720\ : InMux
    port map (
            O => \N__7854\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7847\
        );

    \I__1718\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7844\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7847\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7844\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1715\ : InMux
    port map (
            O => \N__7839\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1714\ : InMux
    port map (
            O => \N__7836\,
            I => \N__7832\
        );

    \I__1713\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7829\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7832\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__7829\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1710\ : InMux
    port map (
            O => \N__7824\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7821\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__7818\,
            I => \N__7815\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7811\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7808\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7805\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7808\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1703\ : Odrv12
    port map (
            O => \N__7805\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1702\ : SRMux
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__7791\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__7788\,
            I => \N__7785\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7774\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7774\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7766\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7766\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7766\
        );

    \I__1692\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7761\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7761\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7774\,
            I => \N__7756\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7753\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7750\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7747\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7742\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7742\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__7756\,
            I => \N__7737\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7737\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__7750\,
            I => \N__7734\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__7747\,
            I => \N__7729\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7729\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7725\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__7734\,
            I => \N__7720\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__7729\,
            I => \N__7720\
        );

    \I__1676\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7717\
        );

    \I__1675\ : Sp12to4
    port map (
            O => \N__7725\,
            I => \N__7712\
        );

    \I__1674\ : Sp12to4
    port map (
            O => \N__7720\,
            I => \N__7712\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7717\,
            I => \N__7709\
        );

    \I__1672\ : Span12Mux_h
    port map (
            O => \N__7712\,
            I => \N__7706\
        );

    \I__1671\ : Span12Mux_h
    port map (
            O => \N__7709\,
            I => \N__7703\
        );

    \I__1670\ : Odrv12
    port map (
            O => \N__7706\,
            I => \RESETn_c\
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__7703\,
            I => \RESETn_c\
        );

    \I__1668\ : IoInMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__1666\ : Span12Mux_s7_v
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__7689\,
            I => \RESETn_c_i\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7683\,
            I => \N__7678\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7675\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7668\
        );

    \I__1660\ : Span4Mux_h
    port map (
            O => \N__7678\,
            I => \N__7663\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7675\,
            I => \N__7663\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7660\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7653\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7653\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7671\,
            I => \N__7653\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7668\,
            I => \N__7650\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__7663\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7660\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7653\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7650\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__7641\,
            I => \N__7638\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__1647\ : Span12Mux_s6_v
    port map (
            O => \N__7635\,
            I => \N__7632\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__7632\,
            I => \RASn_c\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1642\ : Span4Mux_h
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__7617\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7611\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7611\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1638\ : IoInMux
    port map (
            O => \N__7608\,
            I => \N__7605\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1636\ : Span4Mux_s3_h
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1634\ : Span4Mux_h
    port map (
            O => \N__7596\,
            I => \N__7593\
        );

    \I__1633\ : Span4Mux_h
    port map (
            O => \N__7593\,
            I => \N__7590\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__7587\,
            I => \CMA_c_6\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1628\ : Odrv12
    port map (
            O => \N__7578\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1627\ : IoInMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1625\ : IoSpan4Mux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1624\ : IoSpan4Mux
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1623\ : Span4Mux_s2_h
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1622\ : Sp12to4
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1621\ : Span12Mux_h
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__7554\,
            I => \CMA_c_3\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7548\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1617\ : Span12Mux_v
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1616\ : Span12Mux_h
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1615\ : Odrv12
    port map (
            O => \N__7539\,
            I => \A_c_17\
        );

    \I__1614\ : IoInMux
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1612\ : Span4Mux_s3_h
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1609\ : Span4Mux_h
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__7515\,
            I => \CMA_c_8\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7505\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7501\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7496\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__7504\,
            I => \N__7492\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7501\,
            I => \N__7489\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7500\,
            I => \N__7486\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__7499\,
            I => \N__7483\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__7496\,
            I => \N__7480\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__7495\,
            I => \N__7477\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7473\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7489\,
            I => \N__7468\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7486\,
            I => \N__7468\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7465\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__7480\,
            I => \N__7462\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7457\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7457\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7473\,
            I => \N__7454\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__7468\,
            I => \N__7451\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7465\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__7462\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7457\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__7454\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__7451\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7436\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7433\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7430\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7433\,
            I => \N__7427\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__7430\,
            I => \N__7422\
        );

    \I__1577\ : Span4Mux_h
    port map (
            O => \N__7427\,
            I => \N__7419\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7414\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7414\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__7422\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__7419\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7414\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7404\,
            I => \N__7401\
        );

    \I__1569\ : Span12Mux_v
    port map (
            O => \N__7401\,
            I => \N__7398\
        );

    \I__1568\ : Span12Mux_h
    port map (
            O => \N__7398\,
            I => \N__7395\
        );

    \I__1567\ : Odrv12
    port map (
            O => \N__7395\,
            I => \A_c_19\
        );

    \I__1566\ : IoInMux
    port map (
            O => \N__7392\,
            I => \N__7389\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7389\,
            I => \N__7386\
        );

    \I__1564\ : Span4Mux_s3_h
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__1562\ : Span4Mux_h
    port map (
            O => \N__7380\,
            I => \N__7377\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__7377\,
            I => \N__7374\
        );

    \I__1560\ : Span4Mux_h
    port map (
            O => \N__7374\,
            I => \N__7371\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__7371\,
            I => \CMA_c_9\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7364\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7361\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7364\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7361\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7356\,
            I => \bfn_12_8_0_\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7349\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7346\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7349\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7346\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7341\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__7338\,
            I => \N__7335\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7330\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7327\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7324\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7330\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7324\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7313\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7310\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7313\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7310\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7302\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__7293\,
            I => \U712_BYTE_ENABLE.N_271\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__7290\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_\
        );

    \I__1531\ : IoInMux
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7284\,
            I => \N__7281\
        );

    \I__1529\ : IoSpan4Mux
    port map (
            O => \N__7281\,
            I => \N__7278\
        );

    \I__1528\ : Span4Mux_s3_h
    port map (
            O => \N__7278\,
            I => \N__7275\
        );

    \I__1527\ : Sp12to4
    port map (
            O => \N__7275\,
            I => \N__7272\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__7272\,
            I => \N__7269\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7269\,
            I => \N_171_i\
        );

    \I__1524\ : IoInMux
    port map (
            O => \N__7266\,
            I => \N__7263\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1522\ : Span4Mux_s1_v
    port map (
            O => \N__7260\,
            I => \N__7255\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7250\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7250\
        );

    \I__1519\ : Sp12to4
    port map (
            O => \N__7255\,
            I => \N__7247\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7250\,
            I => \N__7244\
        );

    \I__1517\ : Span12Mux_h
    port map (
            O => \N__7247\,
            I => \N__7240\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__7244\,
            I => \N__7237\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7234\
        );

    \I__1514\ : Odrv12
    port map (
            O => \N__7240\,
            I => \DBENn_c\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__7237\,
            I => \DBENn_c\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7234\,
            I => \DBENn_c\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7223\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7220\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7213\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7220\,
            I => \N__7213\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7208\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7208\
        );

    \I__1505\ : Span12Mux_v
    port map (
            O => \N__7213\,
            I => \N__7203\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7200\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7197\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7194\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__7203\,
            I => \DMA_CYCLEm\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__7200\,
            I => \DMA_CYCLEm\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7197\,
            I => \DMA_CYCLEm\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7194\,
            I => \DMA_CYCLEm\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7182\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7182\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7176\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7176\,
            I => \U712_BYTE_ENABLE.N_277\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__7173\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_\
        );

    \I__1492\ : IoInMux
    port map (
            O => \N__7170\,
            I => \N__7167\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__1490\ : Span4Mux_s3_v
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__7161\,
            I => \N__7158\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__7158\,
            I => \N__7155\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__7152\,
            I => \N_150_i\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7143\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7136\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7136\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7136\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7143\,
            I => \U712_BYTE_ENABLE.N_270\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7136\,
            I => \U712_BYTE_ENABLE.N_270\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7128\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7128\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__7125\,
            I => \N__7122\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7119\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7119\,
            I => \U712_BYTE_ENABLE.N_273\
        );

    \I__1474\ : IoInMux
    port map (
            O => \N__7116\,
            I => \N__7113\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7113\,
            I => \N__7110\
        );

    \I__1472\ : IoSpan4Mux
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1471\ : Span4Mux_s2_h
    port map (
            O => \N__7107\,
            I => \N__7104\
        );

    \I__1470\ : Sp12to4
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__1469\ : Span12Mux_h
    port map (
            O => \N__7101\,
            I => \N__7098\
        );

    \I__1468\ : Span12Mux_v
    port map (
            O => \N__7098\,
            I => \N__7095\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__7095\,
            I => \N_172_i\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7086\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7086\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7082\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7079\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__7082\,
            I => \N__7074\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7074\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1459\ : Span12Mux_v
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1458\ : Span12Mux_h
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__7065\,
            I => \CASLn_c\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7062\,
            I => \N__7058\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7053\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7053\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__7050\,
            I => \N__7046\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7043\
        );

    \I__1450\ : Sp12to4
    port map (
            O => \N__7046\,
            I => \N__7038\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7043\,
            I => \N__7038\
        );

    \I__1448\ : Span12Mux_h
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1447\ : Span12Mux_v
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__7032\,
            I => \CASUn_c\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7025\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7022\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7025\,
            I => \N__7017\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__7017\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__7017\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1440\ : IoInMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1438\ : Span12Mux_s4_h
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1437\ : Span12Mux_h
    port map (
            O => \N__7005\,
            I => \N__7002\
        );

    \I__1436\ : Odrv12
    port map (
            O => \N__7002\,
            I => \WEn_c\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6996\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6996\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6990\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6990\,
            I => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6984\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6973\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6973\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6970\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6967\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6973\,
            I => \N__6962\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6970\,
            I => \N__6962\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6967\,
            I => \N__6959\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__1421\ : Span12Mux_v
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1420\ : Sp12to4
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1419\ : Span12Mux_h
    port map (
            O => \N__6953\,
            I => \N__6945\
        );

    \I__1418\ : Span12Mux_v
    port map (
            O => \N__6950\,
            I => \N__6945\
        );

    \I__1417\ : Odrv12
    port map (
            O => \N__6945\,
            I => \CLK40_PLL_i\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6936\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6929\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6929\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6929\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6936\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6929\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6920\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6917\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6920\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6917\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__6903\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__6900\,
            I => \N__6896\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__6899\,
            I => \N__6893\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6890\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6887\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6890\,
            I => \N__6884\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6887\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1396\ : Odrv12
    port map (
            O => \N__6884\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__6873\,
            I => \U712_BYTE_ENABLE.N_275\
        );

    \I__1392\ : IoInMux
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1390\ : Span4Mux_s1_h
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__1389\ : Span4Mux_h
    port map (
            O => \N__6861\,
            I => \N__6858\
        );

    \I__1388\ : Sp12to4
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1387\ : Span12Mux_s11_v
    port map (
            O => \N__6855\,
            I => \N__6852\
        );

    \I__1386\ : Span12Mux_h
    port map (
            O => \N__6852\,
            I => \N__6849\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__6849\,
            I => \N_148_i\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6839\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6836\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__6839\,
            I => \N__6833\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6830\
        );

    \I__1379\ : Sp12to4
    port map (
            O => \N__6833\,
            I => \N__6827\
        );

    \I__1378\ : Sp12to4
    port map (
            O => \N__6830\,
            I => \N__6824\
        );

    \I__1377\ : Span12Mux_h
    port map (
            O => \N__6827\,
            I => \N__6821\
        );

    \I__1376\ : Span12Mux_v
    port map (
            O => \N__6824\,
            I => \N__6818\
        );

    \I__1375\ : Span12Mux_v
    port map (
            O => \N__6821\,
            I => \N__6813\
        );

    \I__1374\ : Span12Mux_h
    port map (
            O => \N__6818\,
            I => \N__6813\
        );

    \I__1373\ : Odrv12
    port map (
            O => \N__6813\,
            I => \RnW_c\
        );

    \I__1372\ : IoInMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1370\ : Span4Mux_s1_h
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1368\ : Span12Mux_s8_v
    port map (
            O => \N__6798\,
            I => \N__6795\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__6792\,
            I => \N_212\
        );

    \I__1365\ : IoInMux
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6786\,
            I => \N__6782\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6779\
        );

    \I__1362\ : Span4Mux_s3_v
    port map (
            O => \N__6782\,
            I => \N__6776\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6773\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__6776\,
            I => \N__6770\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__6773\,
            I => \N__6767\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__6770\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__6767\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1356\ : IoInMux
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1354\ : Span12Mux_s2_v
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1353\ : Odrv12
    port map (
            O => \N__6753\,
            I => \CMA_c_2\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6747\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6732\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6723\,
            I => \N__6718\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6715\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6712\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__6718\,
            I => \N__6707\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6715\,
            I => \N__6707\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6712\,
            I => \N__6704\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__6707\,
            I => \N__6701\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__6704\,
            I => \N__6698\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__6701\,
            I => \N__6695\
        );

    \I__1334\ : Sp12to4
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1333\ : Sp12to4
    port map (
            O => \N__6695\,
            I => \N__6689\
        );

    \I__1332\ : Span12Mux_h
    port map (
            O => \N__6692\,
            I => \N__6686\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6689\,
            I => \AWEn_c\
        );

    \I__1330\ : Odrv12
    port map (
            O => \N__6686\,
            I => \AWEn_c\
        );

    \I__1329\ : IoInMux
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1327\ : Span4Mux_s3_v
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__6669\,
            I => \N__6665\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6662\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6665\,
            I => \DBDIR_c\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6662\,
            I => \DBDIR_c\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__6651\,
            I => \N__6647\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6644\
        );

    \I__1317\ : Odrv4
    port map (
            O => \N__6647\,
            I => \U712_CHIP_RAM.N_298\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6644\,
            I => \U712_CHIP_RAM.N_298\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__6639\,
            I => \N__6632\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__6638\,
            I => \N__6628\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6625\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6622\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6619\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6616\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6609\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6609\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6625\,
            I => \N__6601\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6622\,
            I => \N__6601\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6619\,
            I => \N__6601\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6616\,
            I => \N__6598\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6595\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6589\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6609\,
            I => \N__6586\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6583\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__6601\,
            I => \N__6580\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__6598\,
            I => \N__6575\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6595\,
            I => \N__6575\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6568\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6568\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6568\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6589\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__6586\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6583\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__6580\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__6575\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6552\,
            I => \N__6546\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6543\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6539\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6536\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__6546\,
            I => \N__6529\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6543\,
            I => \N__6529\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6526\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6523\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6520\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6515\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6515\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__6529\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6526\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__6523\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__6520\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6515\,
            I => \U712_CHIP_RAM.N_355\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__6504\,
            I => \N__6499\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6496\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6491\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6491\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6496\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6491\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6481\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6478\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6475\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6472\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6478\,
            I => \N__6469\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6465\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__6472\,
            I => \N__6462\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__6469\,
            I => \N__6459\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6456\
        );

    \I__1255\ : Odrv12
    port map (
            O => \N__6465\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__6462\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__6459\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6456\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6440\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6435\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6440\,
            I => \N__6432\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6429\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6426\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6435\,
            I => \N__6423\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__6432\,
            I => \N__6418\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6418\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6415\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__6423\,
            I => \N__6409\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__6418\,
            I => \N__6404\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__6415\,
            I => \N__6404\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6397\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6397\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6397\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__6409\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6404\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6397\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6381\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6378\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6373\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6373\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__6381\,
            I => \N__6368\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6368\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6373\,
            I => \N__6365\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__6368\,
            I => \N__6362\
        );

    \I__1223\ : Odrv12
    port map (
            O => \N__6365\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6362\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1221\ : IoInMux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__1219\ : Span12Mux_s1_h
    port map (
            O => \N__6351\,
            I => \N__6348\
        );

    \I__1218\ : Span12Mux_v
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1217\ : Span12Mux_h
    port map (
            O => \N__6345\,
            I => \N__6341\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6338\
        );

    \I__1215\ : Odrv12
    port map (
            O => \N__6341\,
            I => \TACK_OUTn\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6338\,
            I => \TACK_OUTn\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6327\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6327\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6327\,
            I => \N__6322\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6317\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6317\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__6322\,
            I => \N__6314\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__6314\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__6311\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__6306\,
            I => \N__6301\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6296\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6296\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6293\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6290\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6293\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__6290\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6276\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6276\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6276\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6273\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__6270\,
            I => \N__6266\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6263\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__6266\,
            I => \N__6260\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6263\,
            I => \N__6257\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__6257\,
            I => \N__6251\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__6254\,
            I => \N__6246\
        );

    \I__1185\ : Span12Mux_v
    port map (
            O => \N__6251\,
            I => \N__6246\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__6246\,
            I => \A_c_1\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6234\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6234\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6234\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6231\
        );

    \I__1179\ : Span4Mux_v
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__1178\ : Sp12to4
    port map (
            O => \N__6228\,
            I => \N__6225\
        );

    \I__1177\ : Span12Mux_v
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__1176\ : Span12Mux_h
    port map (
            O => \N__6222\,
            I => \N__6219\
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__6219\,
            I => \SIZ_c_1\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6213\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6209\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6206\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__6209\,
            I => \N__6203\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6206\,
            I => \N__6200\
        );

    \I__1169\ : Span4Mux_v
    port map (
            O => \N__6203\,
            I => \N__6194\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6191\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__6194\,
            I => \REG_CYCLEm\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6191\,
            I => \REG_CYCLEm\
        );

    \I__1164\ : IoInMux
    port map (
            O => \N__6186\,
            I => \N__6183\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6180\
        );

    \I__1162\ : Span4Mux_s2_v
    port map (
            O => \N__6180\,
            I => \N__6177\
        );

    \I__1161\ : Span4Mux_h
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__6174\,
            I => \N__6171\
        );

    \I__1159\ : Sp12to4
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__1158\ : Span12Mux_s11_v
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__6165\,
            I => \DRDENn_c\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__6162\,
            I => \N__6159\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6159\,
            I => \N__6156\
        );

    \I__1154\ : IoSpan4Mux
    port map (
            O => \N__6156\,
            I => \N__6153\
        );

    \I__1153\ : IoSpan4Mux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__1152\ : Span4Mux_s1_v
    port map (
            O => \N__6150\,
            I => \N__6147\
        );

    \I__1151\ : Sp12to4
    port map (
            O => \N__6147\,
            I => \N__6144\
        );

    \I__1150\ : Span12Mux_s9_v
    port map (
            O => \N__6144\,
            I => \N__6141\
        );

    \I__1149\ : Odrv12
    port map (
            O => \N__6141\,
            I => \un1_LDSn_i_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6129\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6129\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6129\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6129\,
            I => \N__6126\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__6126\,
            I => \N__6120\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6115\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6115\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6112\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__6120\,
            I => \N__6107\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6107\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6104\
        );

    \I__1137\ : Span4Mux_v
    port map (
            O => \N__6107\,
            I => \N__6101\
        );

    \I__1136\ : Sp12to4
    port map (
            O => \N__6104\,
            I => \N__6098\
        );

    \I__1135\ : Sp12to4
    port map (
            O => \N__6101\,
            I => \N__6095\
        );

    \I__1134\ : Span12Mux_v
    port map (
            O => \N__6098\,
            I => \N__6092\
        );

    \I__1133\ : Span12Mux_h
    port map (
            O => \N__6095\,
            I => \N__6089\
        );

    \I__1132\ : Odrv12
    port map (
            O => \N__6092\,
            I => \A_c_0\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__6089\,
            I => \A_c_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6081\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6081\,
            I => \N__6077\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__6077\,
            I => \N__6070\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6065\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6065\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6070\,
            I => \N__6060\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6060\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6060\,
            I => \N__6057\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__6057\,
            I => \N__6054\
        );

    \I__1120\ : Sp12to4
    port map (
            O => \N__6054\,
            I => \N__6051\
        );

    \I__1119\ : Span12Mux_h
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1118\ : Odrv12
    port map (
            O => \N__6048\,
            I => \SIZ_c_0\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6039\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6039\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6039\,
            I => \N__6036\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__6036\,
            I => \N__6033\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6033\,
            I => \N__6029\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6026\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__6029\,
            I => \DS_ENm\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6026\,
            I => \DS_ENm\
        );

    \I__1109\ : IoInMux
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__1107\ : Span12Mux_s9_v
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__1106\ : Span12Mux_h
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__6009\,
            I => \un1_UDSn_i_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__6000\,
            I => \U712_CHIP_RAM.N_242\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__5988\,
            I => \U712_CHIP_RAM.DBENn_7_0\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__5979\,
            I => \U712_CHIP_RAM.N_253\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__5976\,
            I => \N__5973\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5969\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5966\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5969\,
            I => \REG_TACK\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5966\,
            I => \REG_TACK\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5958\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5951\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5948\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5951\,
            I => \N__5945\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5948\,
            I => \N__5942\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__5945\,
            I => \N__5937\
        );

    \I__1082\ : Span4Mux_h
    port map (
            O => \N__5942\,
            I => \N__5934\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5931\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5928\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__5937\,
            I => \U712_REG_SM.N_188\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__5934\,
            I => \U712_REG_SM.N_188\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5931\,
            I => \U712_REG_SM.N_188\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5928\,
            I => \U712_REG_SM.N_188\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5919\,
            I => \N__5914\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5911\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5908\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5905\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5902\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5908\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5905\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__5902\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__1064\ : Sp12to4
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__1063\ : Span12Mux_h
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1062\ : Odrv12
    port map (
            O => \N__5880\,
            I => \RAS1n_c\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5873\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5873\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5870\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5860\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5855\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5855\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5860\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5855\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5843\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5839\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5836\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5833\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5839\,
            I => \N__5830\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__5836\,
            I => \U712_REG_SM.N_200\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5833\,
            I => \U712_REG_SM.N_200\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__5830\,
            I => \U712_REG_SM.N_200\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__5823\,
            I => \N__5818\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5814\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5821\,
            I => \N__5811\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5808\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5805\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5800\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5800\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5808\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5805\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__5800\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5790\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5790\,
            I => \N__5787\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__5787\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5781\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1026\ : IoInMux
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5766\
        );

    \I__1024\ : IoSpan4Mux
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__1023\ : Sp12to4
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__1022\ : Span12Mux_s9_v
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__5757\,
            I => \CMA_c_1\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5751\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5751\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5745\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5745\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__5742\,
            I => \N__5739\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__1014\ : IoSpan4Mux
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__1013\ : IoSpan4Mux
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__1012\ : Sp12to4
    port map (
            O => \N__5730\,
            I => \N__5727\
        );

    \I__1011\ : Span12Mux_s9_h
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__5724\,
            I => \CMA_c_5\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__1007\ : Span12Mux_v
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__1006\ : Span12Mux_h
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__1005\ : Odrv12
    port map (
            O => \N__5709\,
            I => \A_c_6\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1002\ : Span12Mux_h
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__1001\ : Odrv12
    port map (
            O => \N__5697\,
            I => \A_c_13\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__5694\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__999\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__997\ : Span12Mux_v
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__996\ : Span12Mux_h
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__995\ : Odrv12
    port map (
            O => \N__5679\,
            I => \A_c_4\
        );

    \I__994\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5673\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5670\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__991\ : Sp12to4
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__990\ : Span12Mux_h
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__989\ : Odrv12
    port map (
            O => \N__5661\,
            I => \A_c_11\
        );

    \I__988\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5655\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__985\ : Span4Mux_v
    port map (
            O => \N__5649\,
            I => \N__5646\
        );

    \I__984\ : Sp12to4
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__983\ : Span12Mux_h
    port map (
            O => \N__5643\,
            I => \N__5640\
        );

    \I__982\ : Odrv12
    port map (
            O => \N__5640\,
            I => \A_c_7\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.N_324_cascade_\
        );

    \I__980\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5631\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__978\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5620\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__5627\,
            I => \N__5617\
        );

    \I__976\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5610\
        );

    \I__975\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5610\
        );

    \I__974\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5597\
        );

    \I__973\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5597\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5620\,
            I => \N__5593\
        );

    \I__971\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5590\
        );

    \I__970\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5587\
        );

    \I__969\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5579\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5610\,
            I => \N__5576\
        );

    \I__967\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5573\
        );

    \I__966\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5570\
        );

    \I__965\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5563\
        );

    \I__964\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5563\
        );

    \I__963\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5563\
        );

    \I__962\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5556\
        );

    \I__961\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5556\
        );

    \I__960\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5556\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5597\,
            I => \N__5553\
        );

    \I__958\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5550\
        );

    \I__957\ : Span4Mux_h
    port map (
            O => \N__5593\,
            I => \N__5543\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5590\,
            I => \N__5543\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5587\,
            I => \N__5543\
        );

    \I__954\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5538\
        );

    \I__953\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5538\
        );

    \I__952\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5531\
        );

    \I__951\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5531\
        );

    \I__950\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5531\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5579\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__5576\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5573\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5556\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__5553\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5550\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__5543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5538\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5531\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__5508\,
            I => \N__5504\
        );

    \I__937\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5500\
        );

    \I__936\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5497\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__5503\,
            I => \N__5487\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5482\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5474\
        );

    \I__932\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5469\
        );

    \I__931\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5469\
        );

    \I__930\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5466\
        );

    \I__929\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5459\
        );

    \I__928\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5459\
        );

    \I__927\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5459\
        );

    \I__926\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5456\
        );

    \I__925\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5449\
        );

    \I__924\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5449\
        );

    \I__923\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5449\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__5482\,
            I => \N__5446\
        );

    \I__921\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5443\
        );

    \I__920\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5440\
        );

    \I__919\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5437\
        );

    \I__918\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5432\
        );

    \I__917\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5432\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__5474\,
            I => \N__5423\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5469\,
            I => \N__5423\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5423\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5423\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5418\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5418\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__5446\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5443\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5440\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5437\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5432\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__5418\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__903\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5400\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5400\,
            I => \N__5394\
        );

    \I__901\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5391\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5398\,
            I => \N__5387\
        );

    \I__899\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5382\
        );

    \I__898\ : Span4Mux_h
    port map (
            O => \N__5394\,
            I => \N__5379\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5391\,
            I => \N__5376\
        );

    \I__896\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5373\
        );

    \I__895\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5368\
        );

    \I__894\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5368\
        );

    \I__893\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5365\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5382\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__5379\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5368\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__886\ : IoInMux
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__884\ : IoSpan4Mux
    port map (
            O => \N__5346\,
            I => \N__5343\
        );

    \I__883\ : Span4Mux_s1_h
    port map (
            O => \N__5343\,
            I => \N__5340\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__880\ : Span12Mux_s10_h
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__5331\,
            I => \CLK_EN_c\
        );

    \I__878\ : CEMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5325\,
            I => \N__5322\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__5322\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5319\,
            I => \U712_REG_SM.N_204_cascade_\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__873\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5308\
        );

    \I__872\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5305\
        );

    \I__871\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5302\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5308\,
            I => \U712_REG_SM.N_215\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5305\,
            I => \U712_REG_SM.N_215\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5302\,
            I => \U712_REG_SM.N_215\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__5295\,
            I => \N__5291\
        );

    \I__866\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5288\
        );

    \I__865\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5288\,
            I => \U712_REG_SM.N_204\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U712_REG_SM.N_204\
        );

    \I__862\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5275\
        );

    \I__861\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5270\
        );

    \I__860\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5270\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5275\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__857\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5262\,
            I => \N__5258\
        );

    \I__855\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5255\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__5258\,
            I => \N__5250\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5250\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__850\ : Sp12to4
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__849\ : Span12Mux_h
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__5238\,
            I => \TSn_c\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__846\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__842\ : Sp12to4
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__841\ : Span12Mux_h
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__840\ : Odrv12
    port map (
            O => \N__5214\,
            I => \REGSPACEn_c\
        );

    \I__839\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5205\
        );

    \I__838\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5205\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5205\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__836\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5198\
        );

    \I__835\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5195\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U712_REG_SM.N_209\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5195\,
            I => \U712_REG_SM.N_209\
        );

    \I__832\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5180\
        );

    \I__831\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5180\
        );

    \I__830\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5180\
        );

    \I__829\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5177\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5177\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__826\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5165\
        );

    \I__825\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5165\
        );

    \I__824\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5162\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5165\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa\
        );

    \I__821\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5152\
        );

    \I__820\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5147\
        );

    \I__819\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5147\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5147\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__816\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5136\
        );

    \I__815\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5136\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5136\,
            I => \N__5133\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__5133\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__812\ : IoInMux
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5127\,
            I => \N__5124\
        );

    \I__810\ : Span4Mux_s0_v
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__809\ : Sp12to4
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__808\ : Span12Mux_h
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__807\ : Odrv12
    port map (
            O => \N__5115\,
            I => \CMA_c_10\
        );

    \I__806\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5106\
        );

    \I__805\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5106\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5106\,
            I => \CPU_TACKm\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \N__5096\
        );

    \I__802\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5091\
        );

    \I__801\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5091\
        );

    \I__800\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5088\
        );

    \I__799\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5083\
        );

    \I__798\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5083\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5080\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5077\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5072\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5080\,
            I => \N__5072\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__5077\,
            I => \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__5072\,
            I => \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__790\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__787\ : Sp12to4
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__786\ : Span12Mux_h
    port map (
            O => \N__5052\,
            I => \N__5049\
        );

    \I__785\ : Span12Mux_v
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__5046\,
            I => \RAMSPACEn_c\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__5043\,
            I => \N__5039\
        );

    \I__782\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5036\
        );

    \I__781\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5033\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5036\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5033\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__778\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5022\
        );

    \I__777\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5022\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5022\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__774\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5010\
        );

    \I__773\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5010\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__771\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U712_REG_SM.N_197\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__5001\,
            I => \U712_REG_SM.N_215_cascade_\
        );

    \I__768\ : IoInMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__766\ : IoInMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__765\ : Span4Mux_s2_v
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4982\
        );

    \I__763\ : Span4Mux_h
    port map (
            O => \N__4985\,
            I => \N__4979\
        );

    \I__762\ : IoSpan4Mux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__4979\,
            I => \N__4973\
        );

    \I__760\ : IoSpan4Mux
    port map (
            O => \N__4976\,
            I => \N__4970\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__4973\,
            I => \N__4967\
        );

    \I__758\ : Sp12to4
    port map (
            O => \N__4970\,
            I => \N__4964\
        );

    \I__757\ : Span12Mux_h
    port map (
            O => \N__4967\,
            I => \N__4958\
        );

    \I__756\ : Span12Mux_s6_v
    port map (
            O => \N__4964\,
            I => \N__4958\
        );

    \I__755\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4955\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__4958\,
            I => \ASn_c\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4955\,
            I => \ASn_c\
        );

    \I__752\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4943\
        );

    \I__751\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4943\
        );

    \I__750\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4938\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4943\,
            I => \N__4935\
        );

    \I__748\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4932\
        );

    \I__747\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4929\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4938\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__4935\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4932\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4929\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__741\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4907\
        );

    \I__739\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4904\
        );

    \I__738\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4900\
        );

    \I__737\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4895\
        );

    \I__736\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4895\
        );

    \I__735\ : Span4Mux_v
    port map (
            O => \N__4907\,
            I => \N__4890\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4890\
        );

    \I__733\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4887\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4900\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4895\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4890\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__728\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4875\,
            I => \U712_REG_SM.N_185\
        );

    \I__726\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4865\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__4871\,
            I => \N__4861\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__4870\,
            I => \N__4857\
        );

    \I__723\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4846\
        );

    \I__722\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4846\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4843\
        );

    \I__720\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4840\
        );

    \I__719\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4837\
        );

    \I__718\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4834\
        );

    \I__717\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4831\
        );

    \I__716\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4826\
        );

    \I__715\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4826\
        );

    \I__714\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4821\
        );

    \I__713\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4821\
        );

    \I__712\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4816\
        );

    \I__711\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4816\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4813\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4840\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4837\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4834\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4831\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4826\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4821\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4816\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__4813\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__700\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4791\,
            I => \U712_CHIP_RAM.N_198_i\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__4788\,
            I => \N__4784\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__4787\,
            I => \N__4781\
        );

    \I__696\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4778\
        );

    \I__695\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4772\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4778\,
            I => \N__4769\
        );

    \I__693\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4766\
        );

    \I__692\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4763\
        );

    \I__691\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4760\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4772\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4766\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4763\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U712_CHIP_RAM.N_187\
        );

    \I__685\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4745\
        );

    \I__684\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4742\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4745\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4742\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__681\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4733\
        );

    \I__680\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4730\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4733\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4730\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \N__4721\
        );

    \I__676\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4718\
        );

    \I__675\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__672\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4706\
        );

    \I__671\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4703\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4706\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__4698\,
            I => \U712_CHIP_RAM.N_355_cascade_\
        );

    \I__667\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__4689\,
            I => \N__4685\
        );

    \I__664\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4682\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4685\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__661\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4674\,
            I => \U712_CHIP_RAM.N_235\
        );

    \I__659\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4666\
        );

    \I__658\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4663\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4669\,
            I => \N__4655\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4666\,
            I => \N__4651\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4648\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4644\
        );

    \I__653\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4639\
        );

    \I__652\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4636\
        );

    \I__651\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4633\
        );

    \I__650\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4630\
        );

    \I__649\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4625\
        );

    \I__648\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4625\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__4651\,
            I => \N__4622\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__4648\,
            I => \N__4619\
        );

    \I__645\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4614\
        );

    \I__644\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4614\
        );

    \I__643\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4609\
        );

    \I__642\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4609\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4604\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4604\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4633\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4625\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4622\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4619\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4614\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4609\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__4604\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__631\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4580\
        );

    \I__629\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__628\ : Span4Mux_h
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4577\,
            I => \U712_CHIP_RAM.N_217\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__4574\,
            I => \U712_CHIP_RAM.N_217\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_\
        );

    \I__624\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__622\ : Span4Mux_h
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__4557\,
            I => \U712_CHIP_RAM.N_219\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__4554\,
            I => \U712_CHIP_RAM.N_117_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4548\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1\
        );

    \I__617\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4538\
        );

    \I__616\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4538\
        );

    \I__615\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4535\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4535\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__612\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4524\
        );

    \I__611\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4524\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4524\,
            I => \U712_CHIP_RAM.N_42_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__607\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4512\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__605\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4506\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0\
        );

    \I__603\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4500\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4497\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__4494\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4491\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4482\
        );

    \I__597\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4482\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__594\ : Span4Mux_h
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__593\ : Sp12to4
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__4470\,
            I => \A_c_14\
        );

    \I__591\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4464\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__589\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4446\,
            I => \A_c_15\
        );

    \I__583\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__581\ : Sp12to4
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__580\ : Span12Mux_v
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__579\ : Span12Mux_h
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__578\ : Odrv12
    port map (
            O => \N__4428\,
            I => \A_c_8\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__4425\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4422\,
            I => \U712_REG_SM.N_185_cascade_\
        );

    \I__575\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4412\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__4412\,
            I => \N__4406\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4403\
        );

    \I__570\ : Sp12to4
    port map (
            O => \N__4406\,
            I => \N__4400\
        );

    \I__569\ : Span4Mux_s3_h
    port map (
            O => \N__4403\,
            I => \N__4397\
        );

    \I__568\ : Span12Mux_h
    port map (
            O => \N__4400\,
            I => \N__4392\
        );

    \I__567\ : Sp12to4
    port map (
            O => \N__4397\,
            I => \N__4392\
        );

    \I__566\ : Span12Mux_v
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__565\ : Odrv12
    port map (
            O => \N__4389\,
            I => \C1_c\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__4386\,
            I => \U712_REG_SM.N_197_cascade_\
        );

    \I__563\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4376\
        );

    \I__562\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__561\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4373\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4376\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4373\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__557\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4361\
        );

    \I__556\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4356\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N__4353\
        );

    \I__554\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4350\
        );

    \I__553\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4347\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__4353\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4350\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4347\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__548\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4330\
        );

    \I__547\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4330\
        );

    \I__546\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4327\
        );

    \I__545\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4324\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4330\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4327\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4324\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__4317\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__4314\,
            I => \N__4308\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__4313\,
            I => \N__4305\
        );

    \I__538\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4298\
        );

    \I__537\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4298\
        );

    \I__536\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4298\
        );

    \I__535\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4295\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4295\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__4290\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_cascade_\
        );

    \I__531\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__530\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4281\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__528\ : InMux
    port map (
            O => \N__4278\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__527\ : InMux
    port map (
            O => \N__4275\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__526\ : InMux
    port map (
            O => \N__4272\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__525\ : InMux
    port map (
            O => \N__4269\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__523\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4260\,
            I => \N__4250\
        );

    \I__521\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4243\
        );

    \I__520\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4243\
        );

    \I__519\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4243\
        );

    \I__518\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4236\
        );

    \I__517\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4236\
        );

    \I__516\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4236\
        );

    \I__515\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4233\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__4250\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4243\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4236\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4233\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__510\ : InMux
    port map (
            O => \N__4224\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__509\ : CEMux
    port map (
            O => \N__4221\,
            I => \N__4217\
        );

    \I__508\ : CEMux
    port map (
            O => \N__4220\,
            I => \N__4214\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4217\,
            I => \U712_CHIP_RAM.N_256_i\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4214\,
            I => \U712_CHIP_RAM.N_256_i\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__4209\,
            I => \U712_CYCLE_TERM.N_207_i_0_en_cascade_\
        );

    \I__504\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__502\ : Span12Mux_v
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__501\ : Odrv12
    port map (
            O => \N__4197\,
            I => \TACK_EN_i_ess\
        );

    \I__500\ : CEMux
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__4188\,
            I => \U712_CYCLE_TERM.N_207_i_0_en_0\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4185\,
            I => \U712_CHIP_RAM.N_242_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__4176\,
            I => \U712_CHIP_RAM.N_319\
        );

    \I__493\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4168\
        );

    \I__492\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4163\
        );

    \I__491\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4163\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4168\,
            I => \N__4160\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__4160\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__487\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4151\
        );

    \I__486\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4148\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4143\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4148\,
            I => \N__4140\
        );

    \I__483\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4137\
        );

    \I__482\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4134\
        );

    \I__481\ : Span4Mux_v
    port map (
            O => \N__4143\,
            I => \N__4129\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4140\,
            I => \N__4129\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4137\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4134\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__4129\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4122\,
            I => \U712_CHIP_RAM.N_319_cascade_\
        );

    \I__475\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4115\
        );

    \I__474\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4112\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4115\,
            I => \U712_CHIP_RAM.N_322\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4112\,
            I => \U712_CHIP_RAM.N_322\
        );

    \I__471\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4102\
        );

    \I__470\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4095\
        );

    \I__469\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4095\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4102\,
            I => \N__4092\
        );

    \I__467\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4089\
        );

    \I__466\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4086\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4095\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__464\ : Odrv4
    port map (
            O => \N__4092\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4089\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4086\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__461\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4072\
        );

    \I__460\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4067\
        );

    \I__459\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4067\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4072\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4067\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__456\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4059\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\
        );

    \I__454\ : InMux
    port map (
            O => \N__4056\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__453\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4050\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__451\ : InMux
    port map (
            O => \N__4047\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__4044\,
            I => \U712_CHIP_RAM.N_187_cascade_\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4041\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__4038\,
            I => \U712_CHIP_RAM.N_264_cascade_\
        );

    \I__447\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4032\,
            I => \U712_CHIP_RAM.N_262\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__4029\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__444\ : CEMux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__4017\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\
        );

    \I__440\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4008\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4008\,
            I => \U712_CHIP_RAM.N_220\
        );

    \I__437\ : InMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4002\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__434\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__3990\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__431\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3984\,
            I => \U712_CHIP_RAM.N_176\
        );

    \I__429\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__426\ : Span4Mux_h
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__425\ : Span4Mux_h
    port map (
            O => \N__3969\,
            I => \N__3966\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__3966\,
            I => \A_c_10\
        );

    \I__423\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3960\,
            I => \N__3957\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__419\ : Span12Mux_h
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__418\ : Span12Mux_v
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__3945\,
            I => \A_c_3\
        );

    \I__416\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__414\ : Span12Mux_v
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__413\ : Odrv12
    port map (
            O => \N__3933\,
            I => \A_c_9\
        );

    \I__412\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__410\ : Span12Mux_v
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__409\ : Span12Mux_v
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__3918\,
            I => \A_c_2\
        );

    \I__407\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__3909\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3906\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_\
        );

    \I__403\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3900\,
            I => \U712_CHIP_RAM.N_193\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__3897\,
            I => \U712_CHIP_RAM.N_177_cascade_\
        );

    \I__400\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3891\,
            I => \U712_CHIP_RAM.N_223\
        );

    \I__398\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3885\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3882\,
            I => \U712_CHIP_RAM.N_223_cascade_\
        );

    \I__395\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3876\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3876\,
            I => \N__3872\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__3875\,
            I => \N__3869\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__3872\,
            I => \N__3866\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3869\,
            I => \N__3863\
        );

    \I__390\ : Sp12to4
    port map (
            O => \N__3866\,
            I => \N__3860\
        );

    \I__389\ : IoSpan4Mux
    port map (
            O => \N__3863\,
            I => \N__3857\
        );

    \I__388\ : Span12Mux_h
    port map (
            O => \N__3860\,
            I => \N__3854\
        );

    \I__387\ : IoSpan4Mux
    port map (
            O => \N__3857\,
            I => \N__3851\
        );

    \I__386\ : Span12Mux_v
    port map (
            O => \N__3854\,
            I => \N__3848\
        );

    \I__385\ : IoSpan4Mux
    port map (
            O => \N__3851\,
            I => \N__3845\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__3848\,
            I => \C3_c\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__3845\,
            I => \C3_c\
        );

    \I__382\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__380\ : Odrv4
    port map (
            O => \N__3834\,
            I => \U712_CHIP_RAM.N_213\
        );

    \I__379\ : IoInMux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__377\ : Span12Mux_s3_v
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__376\ : Odrv12
    port map (
            O => \N__3822\,
            I => \VBENn_c\
        );

    \I__375\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__373\ : Span4Mux_v
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__372\ : Sp12to4
    port map (
            O => \N__3810\,
            I => \N__3807\
        );

    \I__371\ : Span12Mux_h
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__3804\,
            I => \A_c_12\
        );

    \I__369\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__367\ : Span12Mux_v
    port map (
            O => \N__3795\,
            I => \N__3792\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__3792\,
            I => \A_c_5\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__3789\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__364\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__362\ : Span4Mux_h
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__361\ : Sp12to4
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__360\ : Span12Mux_v
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__359\ : Odrv12
    port map (
            O => \N__3771\,
            I => \A_c_18\
        );

    \I__358\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__355\ : Span4Mux_v
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__354\ : Span4Mux_h
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__353\ : Sp12to4
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__3750\,
            I => \A_c_16\
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__3747\,
            I => \U712_CHIP_RAM.N_253_cascade_\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__3744\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_\
        );

    \I__349\ : CEMux
    port map (
            O => \N__3741\,
            I => \N__3738\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__347\ : Sp12to4
    port map (
            O => \N__3735\,
            I => \N__3732\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3732\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__3729\,
            I => \U712_CHIP_RAM.N_298_cascade_\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__3726\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__343\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3716\
        );

    \I__342\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__341\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3713\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3716\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3713\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__338\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3705\,
            I => \U712_CHIP_RAM.N_216\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__3702\,
            I => \U712_CHIP_RAM.N_216_cascade_\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__3699\,
            I => \U712_CHIP_RAM.N_193_cascade_\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3696\,
            I => \U712_CHIP_RAM.N_176_cascade_\
        );

    \I__333\ : IoInMux
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__331\ : IoSpan4Mux
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__330\ : Span4Mux_s1_h
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__329\ : Odrv4
    port map (
            O => \N__3681\,
            I => \CLK40_PLL_i_i\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3675\,
            I => \N__3672\
        );

    \I__326\ : Span4Mux_s3_h
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__325\ : Span4Mux_v
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__3666\,
            I => \N_897_i\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__3663\,
            I => \N__3660\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__321\ : Span4Mux_s2_v
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__320\ : Span4Mux_v
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__319\ : Span4Mux_h
    port map (
            O => \N__3651\,
            I => \N__3648\
        );

    \I__318\ : Odrv4
    port map (
            O => \N__3648\,
            I => \CLK80_PLL_i_i\
        );

    \I__317\ : IoInMux
    port map (
            O => \N__3645\,
            I => \N__3642\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__315\ : IoSpan4Mux
    port map (
            O => \N__3639\,
            I => \N__3636\
        );

    \I__314\ : Span4Mux_s2_v
    port map (
            O => \N__3636\,
            I => \N__3633\
        );

    \I__313\ : Sp12to4
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__312\ : Span12Mux_v
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__311\ : Odrv12
    port map (
            O => \N__3627\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__8866\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__8867\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__8869\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__8870\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__8868\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7698\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4415\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3875\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLK40_OUT_obuf_RNO_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4206\,
            lcout => \N_897_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8127\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4182\,
            in1 => \N__6614\,
            in2 => \_gnd_net_\,
            in3 => \N__4695\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8106\,
            ce => 'H',
            sr => \N__9391\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100010011"
        )
    port map (
            in0 => \N__4107\,
            in1 => \N__4661\,
            in2 => \N__4871\,
            in3 => \N__5603\,
            lcout => \U712_CHIP_RAM.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6592\,
            in2 => \_gnd_net_\,
            in3 => \N__5485\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__5486\,
            in1 => \N__7784\,
            in2 => \_gnd_net_\,
            in3 => \N__5602\,
            lcout => \U712_CHIP_RAM.N_193\,
            ltout => \U712_CHIP_RAM.N_193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__6555\,
            in1 => \N__4583\,
            in2 => \N__3699\,
            in3 => \N__5615\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__6593\,
            in1 => \N__5604\,
            in2 => \N__5503\,
            in3 => \N__4147\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110000"
        )
    port map (
            in0 => \N__6486\,
            in1 => \N__6439\,
            in2 => \N__7788\,
            in3 => \N__6594\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_i_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__4077\,
            in2 => \_gnd_net_\,
            in3 => \N__6385\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8114\,
            ce => \N__3741\,
            sr => \N__9376\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001000100"
        )
    port map (
            in0 => \N__5478\,
            in1 => \N__4100\,
            in2 => \_gnd_net_\,
            in3 => \N__4856\,
            lcout => \U712_CHIP_RAM.N_176\,
            ltout => \U712_CHIP_RAM.N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4647\,
            in1 => \N__4775\,
            in2 => \N__3696\,
            in3 => \N__5586\,
            lcout => \U712_CHIP_RAM.N_253\,
            ltout => \U712_CHIP_RAM.N_253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__6384\,
            in1 => \N__3721\,
            in2 => \N__3747\,
            in3 => \N__5101\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9416\,
            in1 => \_gnd_net_\,
            in2 => \N__3744\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__5477\,
            in2 => \N__4662\,
            in3 => \N__5585\,
            lcout => \U712_CHIP_RAM.N_298\,
            ltout => \U712_CHIP_RAM.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__6636\,
            in1 => \_gnd_net_\,
            in2 => \N__3729\,
            in3 => \N__6549\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIV2P76_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__6484\,
            in2 => \N__6447\,
            in3 => \N__5099\,
            lcout => \U712_CHIP_RAM.N_323\,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__3840\,
            in1 => \_gnd_net_\,
            in2 => \N__3726\,
            in3 => \N__4106\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8118\,
            ce => 'H',
            sr => \N__9369\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILCLN6_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7773\,
            in1 => \N__3723\,
            in2 => \N__5103\,
            in3 => \N__6390\,
            lcout => \U712_CHIP_RAM.N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6637\,
            in1 => \N__3708\,
            in2 => \_gnd_net_\,
            in3 => \N__4155\,
            lcout => \U712_CHIP_RAM.N_220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__5616\,
            in1 => \N__5480\,
            in2 => \_gnd_net_\,
            in3 => \N__4860\,
            lcout => \U712_CHIP_RAM.N_216\,
            ltout => \U712_CHIP_RAM.N_216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4105\,
            in2 => \N__3702\,
            in3 => \N__4658\,
            lcout => \U712_CHIP_RAM.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3879\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8121\,
            ce => 'H',
            sr => \N__9364\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4364\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8121\,
            ce => 'H',
            sr => \N__9364\
        );

    \U712_REG_SM.C3_SYNC_2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4912\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8121\,
            ce => 'H',
            sr => \N__9364\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6123\,
            in1 => \N__6269\,
            in2 => \_gnd_net_\,
            in3 => \N__8496\,
            lcout => \U712_BYTE_ENABLE.N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__6722\,
            in2 => \_gnd_net_\,
            in3 => \N__6438\,
            lcout => \U712_CHIP_RAM.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__8543\,
            in1 => \N__6216\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3819\,
            in1 => \N__3801\,
            in2 => \_gnd_net_\,
            in3 => \N__8339\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8340\,
            in1 => \N__8552\,
            in2 => \N__3789\,
            in3 => \N__9240\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__3786\,
            in2 => \_gnd_net_\,
            in3 => \N__3768\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3981\,
            in1 => \N__3963\,
            in2 => \_gnd_net_\,
            in3 => \N__8338\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3942\,
            in1 => \N__3930\,
            in2 => \_gnd_net_\,
            in3 => \N__8336\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4172\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5399\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4521\,
            in1 => \N__3915\,
            in2 => \N__3906\,
            in3 => \N__3894\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8104\,
            ce => \N__4026\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5623\,
            in1 => \N__6608\,
            in2 => \_gnd_net_\,
            in3 => \N__4146\,
            lcout => \U712_CHIP_RAM.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4660\,
            in2 => \_gnd_net_\,
            in3 => \N__4868\,
            lcout => \U712_CHIP_RAM.N_177\,
            ltout => \U712_CHIP_RAM.N_177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNINB8M4_0_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__3903\,
            in2 => \N__3897\,
            in3 => \N__6550\,
            lcout => \U712_CHIP_RAM.N_223\,
            ltout => \U712_CHIP_RAM.N_223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI63MN7_2_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__4171\,
            in1 => \N__3888\,
            in2 => \N__3882\,
            in3 => \N__4869\,
            lcout => \U712_CHIP_RAM.N_42_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6650\,
            lcout => \U712_CHIP_RAM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6635\,
            in2 => \_gnd_net_\,
            in3 => \N__6534\,
            lcout => \U712_CHIP_RAM.N_187\,
            ltout => \U712_CHIP_RAM.N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__4794\,
            in2 => \N__4044\,
            in3 => \N__4670\,
            lcout => \U712_CHIP_RAM.N_262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5596\,
            in1 => \N__7781\,
            in2 => \N__4870\,
            in3 => \N__5494\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILJN86_2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6386\,
            in1 => \N__5100\,
            in2 => \N__4041\,
            in3 => \N__4776\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ3ENG_3_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4118\,
            in1 => \N__7783\,
            in2 => \N__4038\,
            in3 => \N__4035\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4029\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__4014\,
            in1 => \N__4543\,
            in2 => \N__7499\,
            in3 => \N__4005\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__4253\,
            in1 => \N__7779\,
            in2 => \N__3999\,
            in3 => \N__4053\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8111\,
            ce => \N__4221\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5609\,
            in1 => \N__3987\,
            in2 => \N__4788\,
            in3 => \N__4643\,
            lcout => \U712_CHIP_RAM.N_242\,
            ltout => \U712_CHIP_RAM.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9NL8E_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__4075\,
            in2 => \N__4185\,
            in3 => \N__7780\,
            lcout => \U712_CHIP_RAM.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6615\,
            in1 => \N__5490\,
            in2 => \_gnd_net_\,
            in3 => \N__5385\,
            lcout => \U712_CHIP_RAM.N_319\,
            ltout => \U712_CHIP_RAM.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINL0R5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__4173\,
            in1 => \N__4154\,
            in2 => \N__4122\,
            in3 => \N__4688\,
            lcout => \U712_CHIP_RAM.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4642\,
            in2 => \_gnd_net_\,
            in3 => \N__4851\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4852\,
            in1 => \N__5479\,
            in2 => \N__5627\,
            in3 => \N__4101\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4076\,
            in1 => \N__4515\,
            in2 => \N__4266\,
            in3 => \N__4062\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8111\,
            ce => \N__4221\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5608\,
            in2 => \_gnd_net_\,
            in3 => \N__9093\,
            lcout => \U712_CHIP_RAM.DBENn_7_0\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4257\,
            in1 => \N__5481\,
            in2 => \_gnd_net_\,
            in3 => \N__4056\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4864\,
            in2 => \_gnd_net_\,
            in3 => \N__4047\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4258\,
            in1 => \N__4659\,
            in2 => \_gnd_net_\,
            in3 => \N__4278\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4254\,
            in1 => \N__4724\,
            in2 => \_gnd_net_\,
            in3 => \N__4275\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4259\,
            in1 => \N__4737\,
            in2 => \_gnd_net_\,
            in3 => \N__4272\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4255\,
            in1 => \N__4749\,
            in2 => \_gnd_net_\,
            in3 => \N__4269\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4710\,
            in1 => \N__4256\,
            in2 => \_gnd_net_\,
            in3 => \N__4224\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8115\,
            ce => \N__4220\,
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__7760\,
            in1 => \N__6304\,
            in2 => \N__6900\,
            in3 => \N__6325\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_207_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9414\,
            in1 => \_gnd_net_\,
            in2 => \N__4209\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_207_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__7759\,
            in1 => \N__6305\,
            in2 => \_gnd_net_\,
            in3 => \N__6326\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8119\,
            ce => \N__4194\,
            sr => \N__9354\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_0_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4381\,
            in1 => \N__4335\,
            in2 => \N__4313\,
            in3 => \N__4359\,
            lcout => \U712_REG_SM.N_185\,
            ltout => \U712_REG_SM.N_185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4941\,
            in2 => \N__4422\,
            in3 => \N__4903\,
            lcout => \U712_REG_SM.N_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8122\,
            ce => 'H',
            sr => \N__9346\
        );

    \U712_REG_SM.C1_SYNC_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8122\,
            ce => 'H',
            sr => \N__9346\
        );

    \U712_REG_SM.C1_SYNC_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4338\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8122\,
            ce => 'H',
            sr => \N__9346\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4382\,
            in1 => \N__4336\,
            in2 => \N__4314\,
            in3 => \N__4360\,
            lcout => \U712_REG_SM.N_197\,
            ltout => \U712_REG_SM.N_197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4911\,
            in1 => \_gnd_net_\,
            in2 => \N__4386\,
            in3 => \N__4948\,
            lcout => \U712_REG_SM.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIFFTG1_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4383\,
            in1 => \N__4910\,
            in2 => \N__4368\,
            in3 => \N__4942\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_0_sqmuxa_0_a2_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4286\,
            in1 => \N__4337\,
            in2 => \N__4317\,
            in3 => \N__4311\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa\,
            ltout => \U712_REG_SM.DS_EN_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__5817\,
            in1 => \N__4287\,
            in2 => \N__4290\,
            in3 => \N__5201\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8122\,
            ce => 'H',
            sr => \N__9346\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__7674\,
            in1 => \N__8330\,
            in2 => \N__7504\,
            in3 => \N__8702\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9417\,
            in1 => \_gnd_net_\,
            in2 => \N__4491\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__4488\,
            in1 => \N__7426\,
            in2 => \N__8576\,
            in3 => \N__8889\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__4487\,
            in1 => \N__7425\,
            in2 => \N__8577\,
            in3 => \N__8888\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8334\,
            in1 => \N__4467\,
            in2 => \N__8578\,
            in3 => \N__8751\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__8548\,
            in1 => \N__8636\,
            in2 => \N__8225\,
            in3 => \N__8335\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101111"
        )
    port map (
            in0 => \N__8637\,
            in1 => \N__8544\,
            in2 => \N__8364\,
            in3 => \N__8210\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8341\,
            in1 => \N__4461\,
            in2 => \_gnd_net_\,
            in3 => \N__4443\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001100"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__4872\,
            in2 => \N__5508\,
            in3 => \N__5626\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__4529\,
            in1 => \N__4544\,
            in2 => \N__4425\,
            in3 => \N__7673\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111100100"
        )
    port map (
            in0 => \N__4545\,
            in1 => \N__4530\,
            in2 => \N__8719\,
            in3 => \N__4509\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__7672\,
            in1 => \_gnd_net_\,
            in2 => \N__7495\,
            in3 => \N__8342\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7671\,
            in2 => \_gnd_net_\,
            in3 => \N__7476\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__6485\,
            in1 => \N__6443\,
            in2 => \N__6638\,
            in3 => \N__5625\,
            lcout => \U712_CHIP_RAM.N_236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5607\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__5606\,
            in1 => \N__5493\,
            in2 => \N__5398\,
            in3 => \N__4854\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5492\,
            in1 => \N__5605\,
            in2 => \_gnd_net_\,
            in3 => \N__5386\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__4503\,
            in1 => \N__4671\,
            in2 => \N__4497\,
            in3 => \N__4777\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9415\,
            in1 => \_gnd_net_\,
            in2 => \N__4494\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5491\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \U712_CHIP_RAM.N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5390\,
            in2 => \N__4787\,
            in3 => \N__4677\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4748\,
            in1 => \N__4736\,
            in2 => \N__4725\,
            in3 => \N__4709\,
            lcout => \U712_CHIP_RAM.N_355\,
            ltout => \U712_CHIP_RAM.N_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4698\,
            in3 => \N__5582\,
            lcout => \U712_CHIP_RAM.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__5495\,
            in2 => \_gnd_net_\,
            in3 => \N__4654\,
            lcout => \U712_CHIP_RAM.N_235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__5496\,
            in1 => \N__5584\,
            in2 => \N__4669\,
            in3 => \N__6542\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4587\,
            in1 => \N__8517\,
            in2 => \N__4569\,
            in3 => \N__5397\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__5112\,
            in1 => \N__4566\,
            in2 => \N__4554\,
            in3 => \N__4551\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8108\,
            ce => 'H',
            sr => \N__9365\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5111\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111111"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5961\,
            in2 => \N__5043\,
            in3 => \N__5027\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101011"
        )
    port map (
            in0 => \N__5042\,
            in1 => \N__5265\,
            in2 => \N__5067\,
            in3 => \N__8562\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8112\,
            ce => 'H',
            sr => \N__9355\
        );

    \DBR_SYNC_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5142\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8112\,
            ce => 'H',
            sr => \N__9355\
        );

    \U712_REG_SM.C3_SYNC_RNIBM0G2_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__5028\,
            in1 => \N__5141\,
            in2 => \_gnd_net_\,
            in3 => \N__5940\,
            lcout => \U712_REG_SM.N_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__5187\,
            in1 => \N__5157\,
            in2 => \N__5019\,
            in3 => \N__5312\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8116\,
            ce => 'H',
            sr => \N__9347\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__4950\,
            in1 => \N__5015\,
            in2 => \N__4920\,
            in3 => \N__5007\,
            lcout => \U712_REG_SM.N_215\,
            ltout => \U712_REG_SM.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4963\,
            in2 => \N__5001\,
            in3 => \N__5172\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8116\,
            ce => 'H',
            sr => \N__9347\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4949\,
            in1 => \N__4913\,
            in2 => \_gnd_net_\,
            in3 => \N__4878\,
            lcout => \U712_REG_SM.N_204\,
            ltout => \U712_REG_SM.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__6032\,
            in1 => \N__5279\,
            in2 => \N__5319\,
            in3 => \N__5171\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8116\,
            ce => 'H',
            sr => \N__9347\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__5865\,
            in1 => \N__5278\,
            in2 => \N__5295\,
            in3 => \N__5846\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8116\,
            ce => 'H',
            sr => \N__9347\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__5155\,
            in1 => \N__5210\,
            in2 => \N__5316\,
            in3 => \N__5189\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8120\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__5311\,
            in1 => \N__5280\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8120\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__5261\,
            in1 => \N__5190\,
            in2 => \N__5235\,
            in3 => \N__5211\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8120\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__5202\,
            in1 => \N__5918\,
            in2 => \N__5823\,
            in3 => \N__5941\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8120\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__5156\,
            in1 => \N__5188\,
            in2 => \_gnd_net_\,
            in3 => \N__5170\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8120\,
            ce => 'H',
            sr => \N__9340\
        );

    \DBR_SYNC_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8840\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8123\,
            ce => 'H',
            sr => \N__9338\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7682\,
            in1 => \N__8394\,
            in2 => \N__7512\,
            in3 => \N__8718\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8092\,
            ce => \N__7985\,
            sr => \N__9392\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__5784\,
            in2 => \_gnd_net_\,
            in3 => \N__5778\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8099\,
            ce => \N__7984\,
            sr => \N__9377\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5754\,
            in1 => \N__5748\,
            in2 => \_gnd_net_\,
            in3 => \N__5634\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8099\,
            ce => \N__7984\,
            sr => \N__9377\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5721\,
            in1 => \N__8358\,
            in2 => \_gnd_net_\,
            in3 => \N__5706\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8359\,
            in1 => \N__8530\,
            in2 => \N__5694\,
            in3 => \N__8973\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5691\,
            in1 => \N__8357\,
            in2 => \_gnd_net_\,
            in3 => \N__5676\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5658\,
            in1 => \N__8531\,
            in2 => \_gnd_net_\,
            in3 => \N__9231\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8360\,
            in2 => \N__5637\,
            in3 => \N__8224\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5628\,
            in1 => \N__5507\,
            in2 => \_gnd_net_\,
            in3 => \N__5403\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8102\,
            ce => \N__5328\,
            sr => \N__9366\
        );

    \U712_CHIP_RAM.DBENn_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001011111110"
        )
    port map (
            in0 => \N__7243\,
            in1 => \N__6006\,
            in2 => \N__6504\,
            in3 => \N__5997\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8105\,
            ce => 'H',
            sr => \N__9356\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__7207\,
            in1 => \N__6502\,
            in2 => \_gnd_net_\,
            in3 => \N__5985\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8105\,
            ce => 'H',
            sr => \N__9356\
        );

    \U712_REG_SM.REG_TACK_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011100"
        )
    port map (
            in0 => \N__5821\,
            in1 => \N__5917\,
            in2 => \N__5976\,
            in3 => \N__5955\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8105\,
            ce => 'H',
            sr => \N__9356\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5877\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8109\,
            ce => 'H',
            sr => \N__9348\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__5864\,
            in1 => \N__5842\,
            in2 => \N__5919\,
            in3 => \N__5954\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8109\,
            ce => 'H',
            sr => \N__9348\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__5895\,
            in1 => \N__8948\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8109\,
            ce => 'H',
            sr => \N__9348\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001110"
        )
    port map (
            in0 => \N__5863\,
            in1 => \N__6199\,
            in2 => \N__5850\,
            in3 => \N__5822\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8109\,
            ce => 'H',
            sr => \N__9348\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__7887\,
            in1 => \N__6999\,
            in2 => \N__7818\,
            in3 => \N__6987\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8109\,
            ce => 'H',
            sr => \N__9348\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__6980\,
            in1 => \N__6941\,
            in2 => \N__6306\,
            in3 => \N__6333\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8113\,
            ce => 'H',
            sr => \N__9341\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__6940\,
            in1 => \N__6344\,
            in2 => \N__7338\,
            in3 => \N__6981\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8113\,
            ce => 'H',
            sr => \N__9341\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__7305\,
            in1 => \N__6939\,
            in2 => \N__6899\,
            in3 => \N__6332\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8113\,
            ce => 'H',
            sr => \N__9341\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6138\,
            in1 => \N__6285\,
            in2 => \_gnd_net_\,
            in3 => \N__8569\,
            lcout => \U712_BYTE_ENABLE.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__6283\,
            in1 => \N__6136\,
            in2 => \N__8583\,
            in3 => \N__6241\,
            lcout => \U712_BYTE_ENABLE.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__6284\,
            in1 => \N__6137\,
            in2 => \N__8584\,
            in3 => \N__6242\,
            lcout => \U712_BYTE_ENABLE.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__8570\,
            in1 => \N__6243\,
            in2 => \_gnd_net_\,
            in3 => \N__6084\,
            lcout => \U712_BYTE_ENABLE.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7226\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6212\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__6044\,
            in1 => \N__6124\,
            in2 => \_gnd_net_\,
            in3 => \N__6073\,
            lcout => \un1_LDSn_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111111"
        )
    port map (
            in0 => \N__6125\,
            in1 => \_gnd_net_\,
            in2 => \N__6080\,
            in3 => \N__6045\,
            lcout => \un1_UDSn_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__6721\,
            in1 => \N__6842\,
            in2 => \_gnd_net_\,
            in3 => \N__7227\,
            lcout => \N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8182\,
            in1 => \N__8787\,
            in2 => \N__8257\,
            in3 => \N__6744\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8093\,
            ce => \N__8015\,
            sr => \N__9378\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__6750\,
            in1 => \N__8572\,
            in2 => \N__8398\,
            in3 => \N__8964\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__8571\,
            in1 => \N__9222\,
            in2 => \N__8393\,
            in3 => \N__6738\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__6729\,
            in1 => \N__6503\,
            in2 => \_gnd_net_\,
            in3 => \N__6668\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8100\,
            ce => 'H',
            sr => \N__9357\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6413\,
            in1 => \N__6657\,
            in2 => \N__6639\,
            in3 => \N__6551\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__6414\,
            in1 => \N__7206\,
            in2 => \N__6912\,
            in3 => \N__6993\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8103\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6468\,
            in2 => \_gnd_net_\,
            in3 => \N__6412\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7835\,
            in2 => \_gnd_net_\,
            in3 => \N__7850\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6923\,
            lcout => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__7901\,
            in1 => \N__7352\,
            in2 => \N__7869\,
            in3 => \N__7367\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7317\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8110\,
            ce => 'H',
            sr => \N__9339\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6979\,
            in2 => \_gnd_net_\,
            in3 => \N__6942\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8110\,
            ce => 'H',
            sr => \N__9339\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7029\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8110\,
            ce => 'H',
            sr => \N__9339\
        );

    \U712_CHIP_RAM.CAS_SYNC_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6924\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8110\,
            ce => 'H',
            sr => \N__9339\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7334\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8110\,
            ce => 'H',
            sr => \N__9339\
        );

    \U712_BYTE_ENABLE.N_148_i_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__7185\,
            in1 => \N__6879\,
            in2 => \N__7062\,
            in3 => \N__7146\,
            lcout => \N_148_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7333\,
            in2 => \_gnd_net_\,
            in3 => \N__7316\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7219\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_171_i_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__7299\,
            in1 => \N__7149\,
            in2 => \N__7290\,
            in3 => \N__7061\,
            lcout => \N_171_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7258\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7218\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_150_i_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__7147\,
            in1 => \N__7179\,
            in2 => \N__7173\,
            in3 => \N__7091\,
            lcout => \N_150_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_172_i_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__7148\,
            in1 => \N__7131\,
            in2 => \N__7125\,
            in3 => \N__7092\,
            lcout => \N_172_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7049\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8117\,
            ce => 'H',
            sr => \N__9337\
        );

    \U712_CHIP_RAM.WEn_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7508\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8088\,
            ce => 'H',
            sr => \N__9375\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8386\,
            in1 => \N__8539\,
            in2 => \N__7629\,
            in3 => \N__7911\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496_1_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8538\,
            in2 => \_gnd_net_\,
            in3 => \N__8385\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI4496Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__8184\,
            in1 => \N__8245\,
            in2 => \N__9522\,
            in3 => \N__7614\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8091\,
            ce => \N__8000\,
            sr => \N__9363\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8183\,
            in1 => \N__9174\,
            in2 => \N__8256\,
            in3 => \N__7584\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8091\,
            ce => \N__8000\,
            sr => \N__9363\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__7551\,
            in1 => \N__7439\,
            in2 => \N__8588\,
            in3 => \N__9162\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8091\,
            ce => \N__8000\,
            sr => \N__9363\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7681\,
            in1 => \N__8356\,
            in2 => \N__8720\,
            in3 => \N__7500\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__7440\,
            in1 => \N__7407\,
            in2 => \N__8589\,
            in3 => \N__8922\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8095\,
            ce => \N__8016\,
            sr => \N__9345\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7368\,
            in2 => \_gnd_net_\,
            in3 => \N__7356\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7353\,
            in2 => \_gnd_net_\,
            in3 => \N__7341\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7902\,
            in2 => \_gnd_net_\,
            in3 => \N__7890\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7886\,
            in2 => \_gnd_net_\,
            in3 => \N__7872\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7868\,
            in2 => \_gnd_net_\,
            in3 => \N__7854\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7851\,
            in2 => \_gnd_net_\,
            in3 => \N__7839\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7836\,
            in2 => \_gnd_net_\,
            in3 => \N__7824\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7814\,
            in2 => \_gnd_net_\,
            in3 => \N__7821\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8865\,
            ce => 'H',
            sr => \N__7800\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7728\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_13_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7686\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8089\,
            ce => 'H',
            sr => \N__9393\
        );

    \U712_CHIP_RAM.CASn_LC_13_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8399\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8089\,
            ce => 'H',
            sr => \N__9393\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8721\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8089\,
            ce => 'H',
            sr => \N__9393\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8185\,
            in1 => \N__8793\,
            in2 => \N__8262\,
            in3 => \N__8658\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8090\,
            ce => \N__8008\,
            sr => \N__9385\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7947\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9500\,
            ce => \N__9469\,
            sr => \N__9379\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8186\,
            in1 => \N__9009\,
            in2 => \N__8258\,
            in3 => \N__8622\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8094\,
            ce => \N__8007\,
            sr => \N__9370\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8579\,
            in1 => \N__8412\,
            in2 => \N__8400\,
            in3 => \N__9126\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__8252\,
            in1 => \N__8187\,
            in2 => \N__8151\,
            in3 => \N__9567\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8094\,
            ce => \N__8007\,
            sr => \N__9370\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7940\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9083\,
            sr => \N__9367\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8916\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9083\,
            sr => \N__9367\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9213\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9083\,
            sr => \N__9367\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9498\,
            ce => \N__9451\,
            sr => \N__9358\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8912\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9498\,
            ce => \N__9451\,
            sr => \N__9358\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9413\,
            in1 => \N__8841\,
            in2 => \_gnd_net_\,
            in3 => \N__8874\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__8836\,
            in2 => \_gnd_net_\,
            in3 => \N__9507\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9117\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9502\,
            ce => \N__9474\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9502\,
            ce => \N__9474\,
            sr => \N__9386\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8777\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9082\,
            sr => \N__9380\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9033\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9082\,
            sr => \N__9380\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9555\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9081\,
            sr => \N__9371\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9000\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9081\,
            sr => \N__9371\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9212\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9499\,
            ce => \N__9467\,
            sr => \N__9368\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9499\,
            ce => \N__9467\,
            sr => \N__9368\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9149\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9084\,
            sr => \N__9359\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9116\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__9065\,
            sr => \N__9350\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9503\,
            ce => \N__9468\,
            sr => \N__9387\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8996\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9501\,
            ce => \N__9470\,
            sr => \N__9381\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9551\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9501\,
            ce => \N__9470\,
            sr => \N__9381\
        );
end \INTERFACE\;

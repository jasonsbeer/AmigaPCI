-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 14 2025 20:14:53

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    PRnW : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    BLSn : out std_logic;
    TCIn : out std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \A_c_8\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m104_ns_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_105_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_106_0\ : std_logic;
signal \U712_CHIP_RAM.N_106_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0\ : std_logic;
signal \U712_CHIP_RAM.N_233\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_206_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_214_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.N_216_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_217_0\ : std_logic;
signal \U712_CHIP_RAM.N_216_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_195_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_213_0\ : std_logic;
signal \U712_CHIP_RAM.N_189_0\ : std_logic;
signal \U712_CHIP_RAM.N_195_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_111_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_50\ : std_logic;
signal \U712_CHIP_RAM.m138_0\ : std_logic;
signal \U712_CHIP_RAM.N_352_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_183_0\ : std_logic;
signal \U712_CHIP_RAM.N_137_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_178_0\ : std_logic;
signal \U712_CHIP_RAM.N_94_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_96_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.m92_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_190_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_222_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_358_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m219_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_137_0\ : std_logic;
signal \U712_CHIP_RAM.N_142_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER43\ : std_logic;
signal \U712_CHIP_RAM.m207_ns_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_206_0\ : std_logic;
signal \U712_CHIP_RAM.N_208_0\ : std_logic;
signal \U712_CHIP_RAM.m141_ns_1\ : std_logic;
signal \U712_CHIP_RAM.N_140_0\ : std_logic;
signal \U712_CHIP_RAM.N_140_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_103_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_358\ : std_logic;
signal \U712_CHIP_RAM.N_188_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_344\ : std_logic;
signal \U712_CHIP_RAM.N_96_0\ : std_logic;
signal \U712_CHIP_RAM.m123_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_117_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.m92_0\ : std_logic;
signal \U712_CHIP_RAM.N_130_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.m203_ns_1\ : std_logic;
signal \U712_CHIP_RAM.N_363_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m186_0\ : std_logic;
signal \U712_CHIP_RAM.N_363\ : std_logic;
signal \U712_CHIP_RAM.m225_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_110_0\ : std_logic;
signal \U712_CHIP_RAM.N_112_0\ : std_logic;
signal \U712_CHIP_RAM.N_112_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_94_0\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM_START_RST\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_111_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_359_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_130_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_135_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_125_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_204_0\ : std_logic;
signal \U712_CHIP_RAM.N_120_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_28_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_16_0\ : std_logic;
signal \U712_CHIP_RAM.N_16_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_66_0_cascade_\ : std_logic;
signal \A_c_0\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_168_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_RST_0_i\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \N_10_0_cascade_\ : std_logic;
signal \U712_REG_SM_REG_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.N_84_0_cascade_\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_0\ : std_logic;
signal \i66_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m40_nsZ0Z_1\ : std_logic;
signal \N_10_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_7\ : std_logic;
signal \U712_CHIP_RAM.N_21_0\ : std_logic;
signal \U712_CHIP_RAM.N_21_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_31_0\ : std_logic;
signal \U712_CHIP_RAM.N_329\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_1\ : std_logic;
signal \N_20_0_cascade_\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_2\ : std_logic;
signal \U712_CHIP_RAM.N_37_0\ : std_logic;
signal \N_174_0\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_CHIP_RAM.N_326_mux\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.m154_0_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.m154_0_0\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.m157_xx_mm_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m157_xx_mm_0_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\ : std_logic;
signal \U712_CHIP_RAM.m162_xx_mm_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m162_xx_mm_0_2_cascade_\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM_m45_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM_REG_TACK_7_0\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_8\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_3\ : std_logic;
signal \N_44_0\ : std_logic;
signal \N_175_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM_WRITE_CYCLE\ : std_logic;
signal \N_20_0\ : std_logic;
signal \PRnW_c\ : std_logic;
signal \U712_REG_SM_C3_SYNC_1\ : std_logic;
signal \BLSn_c\ : std_logic;
signal \U712_REG_SM.N_20_0_0\ : std_logic;
signal \N_172_0\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.m161_xx_mm_0_0_cascade_\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.m159_xx_mm_0_0_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.m156_xx_mm_0_2\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m156_xx_mm_0_0\ : std_logic;
signal \N_144_0\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_325\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \N_33_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.m160_xx_mm_0_0\ : std_logic;
signal \U712_CHIP_RAM.m164_0\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.m159_xx_mm_0_2\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.m161_xx_mm_0_2\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.m155_0_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m155_0_2\ : std_logic;
signal \N_68_0\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \N_145_0\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \N_71_0\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.N_36_0_cascade_\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_OUTC_net\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STARTZ0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_ENC_net\ : std_logic;
signal \U712_REG_SM_C1_SYNC_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_33_0_0\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \U712_CHIP_RAM.m160_xx_mm_0_2\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.m228_0\ : std_logic;
signal \U712_CHIP_RAM.N_343\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.N_342\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.N_3_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.m158_xx_mm_0_0\ : std_logic;
signal \U712_CHIP_RAM.m154_a2_0\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.m158_xx_mm_0_2\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_168_0_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\ : std_logic;
signal \N_323_mux\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLEm\ : std_logic;
signal \N_333_mux\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \PRnW_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \BLSn_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    PRnW <= \PRnW_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    BLSn <= \BLSn_wire\;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4517\,
            RESETB => \N__4634\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => \GNDG0\
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13239\,
            DIN => \N__13238\,
            DOUT => \N__13237\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13239\,
            PADOUT => \N__13238\,
            PADIN => \N__13237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13230\,
            DIN => \N__13229\,
            DOUT => \N__13228\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13230\,
            PADOUT => \N__13229\,
            PADIN => \N__13228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13221\,
            DIN => \N__13220\,
            DOUT => \N__13219\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13221\,
            PADOUT => \N__13220\,
            PADIN => \N__13219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10595\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13212\,
            DIN => \N__13211\,
            DOUT => \N__13210\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13212\,
            PADOUT => \N__13211\,
            PADIN => \N__13210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11315\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13203\,
            DIN => \N__13202\,
            DOUT => \N__13201\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13203\,
            PADOUT => \N__13202\,
            PADIN => \N__13201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13194\,
            DIN => \N__13193\,
            DOUT => \N__13192\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13194\,
            PADOUT => \N__13193\,
            PADIN => \N__13192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13185\,
            DIN => \N__13184\,
            DOUT => \N__13183\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13185\,
            PADOUT => \N__13184\,
            PADIN => \N__13183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13176\,
            DIN => \N__13175\,
            DOUT => \N__13174\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13176\,
            PADOUT => \N__13175\,
            PADIN => \N__13174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13167\,
            DIN => \N__13166\,
            DOUT => \N__13165\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13167\,
            PADOUT => \N__13166\,
            PADIN => \N__13165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13158\,
            DIN => \N__13157\,
            DOUT => \N__13156\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13158\,
            PADOUT => \N__13157\,
            PADIN => \N__13156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13149\,
            DIN => \N__13148\,
            DOUT => \N__13147\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13149\,
            PADOUT => \N__13148\,
            PADIN => \N__13147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13140\,
            DIN => \N__13139\,
            DOUT => \N__13138\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13140\,
            PADOUT => \N__13139\,
            PADIN => \N__13138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8543\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13131\,
            DIN => \N__13130\,
            DOUT => \N__13129\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13131\,
            PADOUT => \N__13130\,
            PADIN => \N__13129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13122\,
            DIN => \N__13121\,
            DOUT => \N__13120\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13122\,
            PADOUT => \N__13121\,
            PADIN => \N__13120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13113\,
            DIN => \N__13112\,
            DOUT => \N__13111\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13113\,
            PADOUT => \N__13112\,
            PADIN => \N__13111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5752\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13104\,
            DIN => \N__13103\,
            DOUT => \N__13102\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13104\,
            PADOUT => \N__13103\,
            PADIN => \N__13102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13095\,
            DIN => \N__13094\,
            DOUT => \N__13093\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13095\,
            PADOUT => \N__13094\,
            PADIN => \N__13093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13086\,
            DIN => \N__13085\,
            DOUT => \N__13084\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13086\,
            PADOUT => \N__13085\,
            PADIN => \N__13084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5042\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13077\,
            DIN => \N__13076\,
            DOUT => \N__13075\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13077\,
            PADOUT => \N__13076\,
            PADIN => \N__13075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13068\,
            DIN => \N__13067\,
            DOUT => \N__13066\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13068\,
            PADOUT => \N__13067\,
            PADIN => \N__13066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13059\,
            DIN => \N__13058\,
            DOUT => \N__13057\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13059\,
            PADOUT => \N__13058\,
            PADIN => \N__13057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8384\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13050\,
            DIN => \N__13049\,
            DOUT => \N__13048\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13050\,
            PADOUT => \N__13049\,
            PADIN => \N__13048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13041\,
            DIN => \N__13040\,
            DOUT => \N__13039\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13041\,
            PADOUT => \N__13040\,
            PADIN => \N__13039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13032\,
            DIN => \N__13031\,
            DOUT => \N__13030\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13032\,
            PADOUT => \N__13031\,
            PADIN => \N__13030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13023\,
            DIN => \N__13022\,
            DOUT => \N__13021\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13023\,
            PADOUT => \N__13022\,
            PADIN => \N__13021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13014\,
            DIN => \N__13013\,
            DOUT => \N__13012\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13014\,
            PADOUT => \N__13013\,
            PADIN => \N__13012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9441\,
            DIN0 => OPEN,
            DOUT0 => \N__8898\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13005\,
            DIN => \N__13004\,
            DOUT => \N__13003\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13005\,
            PADOUT => \N__13004\,
            PADIN => \N__13003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12996\,
            DIN => \N__12995\,
            DOUT => \N__12994\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12996\,
            PADOUT => \N__12995\,
            PADIN => \N__12994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12987\,
            DIN => \N__12986\,
            DOUT => \N__12985\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12987\,
            PADOUT => \N__12986\,
            PADIN => \N__12985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12978\,
            DIN => \N__12977\,
            DOUT => \N__12976\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12978\,
            PADOUT => \N__12977\,
            PADIN => \N__12976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12969\,
            DIN => \N__12968\,
            DOUT => \N__12967\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12969\,
            PADOUT => \N__12968\,
            PADIN => \N__12967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12960\,
            DIN => \N__12959\,
            DOUT => \N__12958\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12960\,
            PADOUT => \N__12959\,
            PADIN => \N__12958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9260\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12951\,
            DIN => \N__12950\,
            DOUT => \N__12949\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12951\,
            PADOUT => \N__12950\,
            PADIN => \N__12949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12942\,
            DIN => \N__12941\,
            DOUT => \N__12940\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12942\,
            PADOUT => \N__12941\,
            PADIN => \N__12940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12933\,
            DIN => \N__12932\,
            DOUT => \N__12931\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12933\,
            PADOUT => \N__12932\,
            PADIN => \N__12931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12924\,
            DIN => \N__12923\,
            DOUT => \N__12922\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12924\,
            PADOUT => \N__12923\,
            PADIN => \N__12922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12915\,
            DIN => \N__12914\,
            DOUT => \N__12913\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12915\,
            PADOUT => \N__12914\,
            PADIN => \N__12913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12906\,
            DIN => \N__12905\,
            DOUT => \N__12904\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12906\,
            PADOUT => \N__12905\,
            PADIN => \N__12904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12897\,
            DIN => \N__12896\,
            DOUT => \N__12895\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12897\,
            PADOUT => \N__12896\,
            PADIN => \N__12895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12888\,
            DIN => \N__12887\,
            DOUT => \N__12886\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12888\,
            PADOUT => \N__12887\,
            PADIN => \N__12886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12879\,
            DIN => \N__12878\,
            DOUT => \N__12877\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12879\,
            PADOUT => \N__12878\,
            PADIN => \N__12877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12870\,
            DIN => \N__12869\,
            DOUT => \N__12868\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12870\,
            PADOUT => \N__12869\,
            PADIN => \N__12868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8321\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12861\,
            DIN => \N__12860\,
            DOUT => \N__12859\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12861\,
            PADOUT => \N__12860\,
            PADIN => \N__12859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12852\,
            DIN => \N__12851\,
            DOUT => \N__12850\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12852\,
            PADOUT => \N__12851\,
            PADIN => \N__12850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10175\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12843\,
            DIN => \N__12842\,
            DOUT => \N__12841\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12843\,
            PADOUT => \N__12842\,
            PADIN => \N__12841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8570\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12834\,
            DIN => \N__12833\,
            DOUT => \N__12832\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12834\,
            PADOUT => \N__12833\,
            PADIN => \N__12832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8048\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12825\,
            DIN => \N__12824\,
            DOUT => \N__12823\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12825\,
            PADOUT => \N__12824\,
            PADIN => \N__12823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12816\,
            DIN => \N__12815\,
            DOUT => \N__12814\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12816\,
            PADOUT => \N__12815\,
            PADIN => \N__12814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12807\,
            DIN => \N__12806\,
            DOUT => \N__12805\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12807\,
            PADOUT => \N__12806\,
            PADIN => \N__12805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9445\,
            DIN0 => OPEN,
            DOUT0 => \N__8912\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12798\,
            DIN => \N__12797\,
            DOUT => \N__12796\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12798\,
            PADOUT => \N__12797\,
            PADIN => \N__12796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7961\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12789\,
            DIN => \N__12788\,
            DOUT => \N__12787\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12789\,
            PADOUT => \N__12788\,
            PADIN => \N__12787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4748\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12780\,
            DIN => \N__12779\,
            DOUT => \N__12778\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12780\,
            PADOUT => \N__12779\,
            PADIN => \N__12778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8990\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12771\,
            DIN => \N__12770\,
            DOUT => \N__12769\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12771\,
            PADOUT => \N__12770\,
            PADIN => \N__12769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12762\,
            DIN => \N__12761\,
            DOUT => \N__12760\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12762\,
            PADOUT => \N__12761\,
            PADIN => \N__12760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12753\,
            DIN => \N__12752\,
            DOUT => \N__12751\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12753\,
            PADOUT => \N__12752\,
            PADIN => \N__12751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7604\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12744\,
            DIN => \N__12743\,
            DOUT => \N__12742\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12744\,
            PADOUT => \N__12743\,
            PADIN => \N__12742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12735\,
            DIN => \N__12734\,
            DOUT => \N__12733\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12735\,
            PADOUT => \N__12734\,
            PADIN => \N__12733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12726\,
            DIN => \N__12725\,
            DOUT => \N__12724\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12726\,
            PADOUT => \N__12725\,
            PADIN => \N__12724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7694\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12717\,
            DIN => \N__12716\,
            DOUT => \N__12715\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12717\,
            PADOUT => \N__12716\,
            PADIN => \N__12715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8273\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12708\,
            DIN => \N__12707\,
            DOUT => \N__12706\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12708\,
            PADOUT => \N__12707\,
            PADIN => \N__12706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12699\,
            DIN => \N__12698\,
            DOUT => \N__12697\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12699\,
            PADOUT => \N__12698\,
            PADIN => \N__12697\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12690\,
            DIN => \N__12689\,
            DOUT => \N__12688\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12690\,
            PADOUT => \N__12689\,
            PADIN => \N__12688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9446\,
            DIN0 => OPEN,
            DOUT0 => \N__8911\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12681\,
            DIN => \N__12680\,
            DOUT => \N__12679\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12681\,
            PADOUT => \N__12680\,
            PADIN => \N__12679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6686\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12672\,
            DIN => \N__12671\,
            DOUT => \N__12670\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12672\,
            PADOUT => \N__12671\,
            PADIN => \N__12670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12663\,
            DIN => \N__12662\,
            DOUT => \N__12661\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12663\,
            PADOUT => \N__12662\,
            PADIN => \N__12661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12654\,
            DIN => \N__12653\,
            DOUT => \N__12652\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12654\,
            PADOUT => \N__12653\,
            PADIN => \N__12652\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7859\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12645\,
            DIN => \N__12644\,
            DOUT => \N__12643\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12645\,
            PADOUT => \N__12644\,
            PADIN => \N__12643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12636\,
            DIN => \N__12635\,
            DOUT => \N__12634\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12636\,
            PADOUT => \N__12635\,
            PADIN => \N__12634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12627\,
            DIN => \N__12626\,
            DOUT => \N__12625\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12627\,
            PADOUT => \N__12626\,
            PADIN => \N__12625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12618\,
            DIN => \N__12617\,
            DOUT => \N__12616\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12618\,
            PADOUT => \N__12617\,
            PADIN => \N__12616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12609\,
            DIN => \N__12608\,
            DOUT => \N__12607\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12609\,
            PADOUT => \N__12608\,
            PADIN => \N__12607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12600\,
            DIN => \N__12599\,
            DOUT => \N__12598\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12600\,
            PADOUT => \N__12599\,
            PADIN => \N__12598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12591\,
            DIN => \N__12590\,
            DOUT => \N__12589\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12591\,
            PADOUT => \N__12590\,
            PADIN => \N__12589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7475\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12582\,
            DIN => \N__12581\,
            DOUT => \N__12580\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12582\,
            PADOUT => \N__12581\,
            PADIN => \N__12580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9016\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12573\,
            DIN => \N__12572\,
            DOUT => \N__12571\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12573\,
            PADOUT => \N__12572\,
            PADIN => \N__12571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12564\,
            DIN => \N__12563\,
            DOUT => \N__12562\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12564\,
            PADOUT => \N__12563\,
            PADIN => \N__12562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12555\,
            DIN => \N__12554\,
            DOUT => \N__12553\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12555\,
            PADOUT => \N__12554\,
            PADIN => \N__12553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12546\,
            DIN => \N__12545\,
            DOUT => \N__12544\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12546\,
            PADOUT => \N__12545\,
            PADIN => \N__12544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12537\,
            DIN => \N__12536\,
            DOUT => \N__12535\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12537\,
            PADOUT => \N__12536\,
            PADIN => \N__12535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12528\,
            DIN => \N__12527\,
            DOUT => \N__12526\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12528\,
            PADOUT => \N__12527\,
            PADIN => \N__12526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12519\,
            DIN => \N__12518\,
            DOUT => \N__12517\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12519\,
            PADOUT => \N__12518\,
            PADIN => \N__12517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4544\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12510\,
            DIN => \N__12509\,
            DOUT => \N__12508\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12510\,
            PADOUT => \N__12509\,
            PADIN => \N__12508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12501\,
            DIN => \N__12500\,
            DOUT => \N__12499\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12501\,
            PADOUT => \N__12500\,
            PADIN => \N__12499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRnW_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12492\,
            DIN => \N__12491\,
            DOUT => \N__12490\,
            PACKAGEPIN => \PRnW_wire\
        );

    \PRnW_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12492\,
            PADOUT => \N__12491\,
            PADIN => \N__12490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8150\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12483\,
            DIN => \N__12482\,
            DOUT => \N__12481\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12483\,
            PADOUT => \N__12482\,
            PADIN => \N__12481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12474\,
            DIN => \N__12473\,
            DOUT => \N__12472\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12474\,
            PADOUT => \N__12473\,
            PADIN => \N__12472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12465\,
            DIN => \N__12464\,
            DOUT => \N__12463\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12465\,
            PADOUT => \N__12464\,
            PADIN => \N__12463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12456\,
            DIN => \N__12455\,
            DOUT => \N__12454\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12456\,
            PADOUT => \N__12455\,
            PADIN => \N__12454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10346\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12447\,
            DIN => \N__12446\,
            DOUT => \N__12445\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12447\,
            PADOUT => \N__12446\,
            PADIN => \N__12445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12438\,
            DIN => \N__12437\,
            DOUT => \N__12436\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12438\,
            PADOUT => \N__12437\,
            PADIN => \N__12436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12429\,
            DIN => \N__12428\,
            DOUT => \N__12427\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12429\,
            PADOUT => \N__12428\,
            PADIN => \N__12427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BLSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12420\,
            DIN => \N__12419\,
            DOUT => \N__12418\,
            PACKAGEPIN => \BLSn_wire\
        );

    \BLSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12420\,
            PADOUT => \N__12419\,
            PADIN => \N__12418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12411\,
            DIN => \N__12410\,
            DOUT => \N__12409\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12411\,
            PADOUT => \N__12410\,
            PADIN => \N__12409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12402\,
            DIN => \N__12401\,
            DOUT => \N__12400\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12402\,
            PADOUT => \N__12401\,
            PADIN => \N__12400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12393\,
            DIN => \N__12392\,
            DOUT => \N__12391\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12393\,
            PADOUT => \N__12392\,
            PADIN => \N__12391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10853\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12384\,
            DIN => \N__12383\,
            DOUT => \N__12382\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12384\,
            PADOUT => \N__12383\,
            PADIN => \N__12382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9095\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12375\,
            DIN => \N__12374\,
            DOUT => \N__12373\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12375\,
            PADOUT => \N__12374\,
            PADIN => \N__12373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12366\,
            DIN => \N__12365\,
            DOUT => \N__12364\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12366\,
            PADOUT => \N__12365\,
            PADIN => \N__12364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3007\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12344\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__3005\ : Odrv12
    port map (
            O => \N__12341\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__3004\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__12335\,
            I => \N__12329\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12326\
        );

    \I__3001\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12323\
        );

    \I__3000\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12320\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__12329\,
            I => \N__12313\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__12326\,
            I => \N__12313\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__12323\,
            I => \N__12313\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12308\
        );

    \I__2995\ : Sp12to4
    port map (
            O => \N__12313\,
            I => \N__12308\
        );

    \I__2994\ : Span12Mux_v
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__2993\ : Odrv12
    port map (
            O => \N__12305\,
            I => \DRA_c_3\
        );

    \I__2992\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12296\
        );

    \I__2991\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12293\
        );

    \I__2990\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12290\
        );

    \I__2989\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12287\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__12296\,
            I => \N__12280\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__12293\,
            I => \N__12280\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__12290\,
            I => \N__12280\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__12287\,
            I => \N__12277\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__12277\,
            I => \N__12271\
        );

    \I__2982\ : Span4Mux_v
    port map (
            O => \N__12274\,
            I => \N__12268\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__12271\,
            I => \N__12265\
        );

    \I__2980\ : Sp12to4
    port map (
            O => \N__12268\,
            I => \N__12262\
        );

    \I__2979\ : Sp12to4
    port map (
            O => \N__12265\,
            I => \N__12259\
        );

    \I__2978\ : Span12Mux_h
    port map (
            O => \N__12262\,
            I => \N__12256\
        );

    \I__2977\ : Odrv12
    port map (
            O => \N__12259\,
            I => \DRA_c_4\
        );

    \I__2976\ : Odrv12
    port map (
            O => \N__12256\,
            I => \DRA_c_4\
        );

    \I__2975\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__12245\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__12239\,
            I => \N__12235\
        );

    \I__2970\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12230\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__12235\,
            I => \N__12227\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12224\
        );

    \I__2967\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12221\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12218\
        );

    \I__2965\ : Sp12to4
    port map (
            O => \N__12227\,
            I => \N__12209\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__12224\,
            I => \N__12209\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__12221\,
            I => \N__12209\
        );

    \I__2962\ : Sp12to4
    port map (
            O => \N__12218\,
            I => \N__12209\
        );

    \I__2961\ : Span12Mux_v
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__2960\ : Odrv12
    port map (
            O => \N__12206\,
            I => \DRA_c_2\
        );

    \I__2959\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12200\,
            I => \N__12197\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__12197\,
            I => \N__12194\
        );

    \I__2956\ : Span4Mux_h
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__12191\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2954\ : InMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__2952\ : Span12Mux_h
    port map (
            O => \N__12182\,
            I => \N__12179\
        );

    \I__2951\ : Odrv12
    port map (
            O => \N__12179\,
            I => \RAS1n_c\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12172\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__12172\,
            I => \N__12166\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12163\
        );

    \I__2946\ : Span12Mux_v
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__2945\ : Span12Mux_h
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__2944\ : Odrv12
    port map (
            O => \N__12160\,
            I => \RAS0n_c\
        );

    \I__2943\ : Odrv12
    port map (
            O => \N__12157\,
            I => \RAS0n_c\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12149\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__12149\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__12137\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2936\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12089\
        );

    \I__2934\ : ClkMux
    port map (
            O => \N__12130\,
            I => \N__11975\
        );

    \I__2933\ : ClkMux
    port map (
            O => \N__12129\,
            I => \N__11975\
        );

    \I__2932\ : ClkMux
    port map (
            O => \N__12128\,
            I => \N__11975\
        );

    \I__2931\ : ClkMux
    port map (
            O => \N__12127\,
            I => \N__11975\
        );

    \I__2930\ : ClkMux
    port map (
            O => \N__12126\,
            I => \N__11975\
        );

    \I__2929\ : ClkMux
    port map (
            O => \N__12125\,
            I => \N__11975\
        );

    \I__2928\ : ClkMux
    port map (
            O => \N__12124\,
            I => \N__11975\
        );

    \I__2927\ : ClkMux
    port map (
            O => \N__12123\,
            I => \N__11975\
        );

    \I__2926\ : ClkMux
    port map (
            O => \N__12122\,
            I => \N__11975\
        );

    \I__2925\ : ClkMux
    port map (
            O => \N__12121\,
            I => \N__11975\
        );

    \I__2924\ : ClkMux
    port map (
            O => \N__12120\,
            I => \N__11975\
        );

    \I__2923\ : ClkMux
    port map (
            O => \N__12119\,
            I => \N__11975\
        );

    \I__2922\ : ClkMux
    port map (
            O => \N__12118\,
            I => \N__11975\
        );

    \I__2921\ : ClkMux
    port map (
            O => \N__12117\,
            I => \N__11975\
        );

    \I__2920\ : ClkMux
    port map (
            O => \N__12116\,
            I => \N__11975\
        );

    \I__2919\ : ClkMux
    port map (
            O => \N__12115\,
            I => \N__11975\
        );

    \I__2918\ : ClkMux
    port map (
            O => \N__12114\,
            I => \N__11975\
        );

    \I__2917\ : ClkMux
    port map (
            O => \N__12113\,
            I => \N__11975\
        );

    \I__2916\ : ClkMux
    port map (
            O => \N__12112\,
            I => \N__11975\
        );

    \I__2915\ : ClkMux
    port map (
            O => \N__12111\,
            I => \N__11975\
        );

    \I__2914\ : ClkMux
    port map (
            O => \N__12110\,
            I => \N__11975\
        );

    \I__2913\ : ClkMux
    port map (
            O => \N__12109\,
            I => \N__11975\
        );

    \I__2912\ : ClkMux
    port map (
            O => \N__12108\,
            I => \N__11975\
        );

    \I__2911\ : ClkMux
    port map (
            O => \N__12107\,
            I => \N__11975\
        );

    \I__2910\ : ClkMux
    port map (
            O => \N__12106\,
            I => \N__11975\
        );

    \I__2909\ : ClkMux
    port map (
            O => \N__12105\,
            I => \N__11975\
        );

    \I__2908\ : ClkMux
    port map (
            O => \N__12104\,
            I => \N__11975\
        );

    \I__2907\ : ClkMux
    port map (
            O => \N__12103\,
            I => \N__11975\
        );

    \I__2906\ : ClkMux
    port map (
            O => \N__12102\,
            I => \N__11975\
        );

    \I__2905\ : ClkMux
    port map (
            O => \N__12101\,
            I => \N__11975\
        );

    \I__2904\ : ClkMux
    port map (
            O => \N__12100\,
            I => \N__11975\
        );

    \I__2903\ : ClkMux
    port map (
            O => \N__12099\,
            I => \N__11975\
        );

    \I__2902\ : ClkMux
    port map (
            O => \N__12098\,
            I => \N__11975\
        );

    \I__2901\ : ClkMux
    port map (
            O => \N__12097\,
            I => \N__11975\
        );

    \I__2900\ : ClkMux
    port map (
            O => \N__12096\,
            I => \N__11975\
        );

    \I__2899\ : ClkMux
    port map (
            O => \N__12095\,
            I => \N__11975\
        );

    \I__2898\ : ClkMux
    port map (
            O => \N__12094\,
            I => \N__11975\
        );

    \I__2897\ : ClkMux
    port map (
            O => \N__12093\,
            I => \N__11975\
        );

    \I__2896\ : ClkMux
    port map (
            O => \N__12092\,
            I => \N__11975\
        );

    \I__2895\ : Glb2LocalMux
    port map (
            O => \N__12089\,
            I => \N__11975\
        );

    \I__2894\ : ClkMux
    port map (
            O => \N__12088\,
            I => \N__11975\
        );

    \I__2893\ : ClkMux
    port map (
            O => \N__12087\,
            I => \N__11975\
        );

    \I__2892\ : ClkMux
    port map (
            O => \N__12086\,
            I => \N__11975\
        );

    \I__2891\ : ClkMux
    port map (
            O => \N__12085\,
            I => \N__11975\
        );

    \I__2890\ : ClkMux
    port map (
            O => \N__12084\,
            I => \N__11975\
        );

    \I__2889\ : ClkMux
    port map (
            O => \N__12083\,
            I => \N__11975\
        );

    \I__2888\ : ClkMux
    port map (
            O => \N__12082\,
            I => \N__11975\
        );

    \I__2887\ : ClkMux
    port map (
            O => \N__12081\,
            I => \N__11975\
        );

    \I__2886\ : ClkMux
    port map (
            O => \N__12080\,
            I => \N__11975\
        );

    \I__2885\ : ClkMux
    port map (
            O => \N__12079\,
            I => \N__11975\
        );

    \I__2884\ : ClkMux
    port map (
            O => \N__12078\,
            I => \N__11975\
        );

    \I__2883\ : GlobalMux
    port map (
            O => \N__11975\,
            I => \CLK80_PLL\
        );

    \I__2882\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11968\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__11968\,
            I => \N__11962\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11959\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__11962\,
            I => \N__11956\
        );

    \I__2877\ : Span4Mux_v
    port map (
            O => \N__11959\,
            I => \N__11953\
        );

    \I__2876\ : Sp12to4
    port map (
            O => \N__11956\,
            I => \N__11948\
        );

    \I__2875\ : Sp12to4
    port map (
            O => \N__11953\,
            I => \N__11948\
        );

    \I__2874\ : Span12Mux_h
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__2873\ : Span12Mux_v
    port map (
            O => \N__11945\,
            I => \N__11942\
        );

    \I__2872\ : Odrv12
    port map (
            O => \N__11942\,
            I => \DRA_c_0\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2870\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__11930\,
            I => \N__11920\
        );

    \I__2867\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11913\
        );

    \I__2866\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11913\
        );

    \I__2865\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11910\
        );

    \I__2864\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11907\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \N__11904\
        );

    \I__2862\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11899\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__11923\,
            I => \N__11896\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__11920\,
            I => \N__11889\
        );

    \I__2859\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11886\
        );

    \I__2858\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11883\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__11913\,
            I => \N__11876\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__11910\,
            I => \N__11876\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__11907\,
            I => \N__11876\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11871\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11871\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11866\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11863\
        );

    \I__2850\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11858\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11858\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11894\,
            I => \N__11855\
        );

    \I__2847\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11852\
        );

    \I__2846\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11849\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__11889\,
            I => \N__11840\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11840\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11840\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__11876\,
            I => \N__11840\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__11871\,
            I => \N__11837\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11834\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11831\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__11866\,
            I => \N__11818\
        );

    \I__2837\ : Span4Mux_h
    port map (
            O => \N__11863\,
            I => \N__11818\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11858\,
            I => \N__11818\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11855\,
            I => \N__11818\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11852\,
            I => \N__11818\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__11849\,
            I => \N__11818\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__11840\,
            I => \N__11810\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__11837\,
            I => \N__11810\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11803\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11831\,
            I => \N__11803\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__11818\,
            I => \N__11803\
        );

    \I__2827\ : InMux
    port map (
            O => \N__11817\,
            I => \N__11798\
        );

    \I__2826\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11798\
        );

    \I__2825\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11795\
        );

    \I__2824\ : Sp12to4
    port map (
            O => \N__11810\,
            I => \N__11790\
        );

    \I__2823\ : Sp12to4
    port map (
            O => \N__11803\,
            I => \N__11790\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11798\,
            I => \N__11785\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11785\
        );

    \I__2820\ : Span12Mux_h
    port map (
            O => \N__11790\,
            I => \N__11782\
        );

    \I__2819\ : Span12Mux_h
    port map (
            O => \N__11785\,
            I => \N__11779\
        );

    \I__2818\ : Span12Mux_v
    port map (
            O => \N__11782\,
            I => \N__11776\
        );

    \I__2817\ : Span12Mux_v
    port map (
            O => \N__11779\,
            I => \N__11773\
        );

    \I__2816\ : Odrv12
    port map (
            O => \N__11776\,
            I => \AGNUS_REV_c\
        );

    \I__2815\ : Odrv12
    port map (
            O => \N__11773\,
            I => \AGNUS_REV_c\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11760\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11755\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11755\
        );

    \I__2810\ : Span4Mux_v
    port map (
            O => \N__11760\,
            I => \N__11749\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__2808\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11746\
        );

    \I__2807\ : Sp12to4
    port map (
            O => \N__11749\,
            I => \N__11741\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11741\
        );

    \I__2805\ : Span12Mux_v
    port map (
            O => \N__11741\,
            I => \N__11738\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__11738\,
            I => \DRA_c_1\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__2801\ : Span12Mux_v
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__11726\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2799\ : ClkMux
    port map (
            O => \N__11723\,
            I => \N__11702\
        );

    \I__2798\ : ClkMux
    port map (
            O => \N__11722\,
            I => \N__11702\
        );

    \I__2797\ : ClkMux
    port map (
            O => \N__11721\,
            I => \N__11702\
        );

    \I__2796\ : ClkMux
    port map (
            O => \N__11720\,
            I => \N__11702\
        );

    \I__2795\ : ClkMux
    port map (
            O => \N__11719\,
            I => \N__11702\
        );

    \I__2794\ : ClkMux
    port map (
            O => \N__11718\,
            I => \N__11702\
        );

    \I__2793\ : ClkMux
    port map (
            O => \N__11717\,
            I => \N__11702\
        );

    \I__2792\ : GlobalMux
    port map (
            O => \N__11702\,
            I => \N__11699\
        );

    \I__2791\ : gio2CtrlBuf
    port map (
            O => \N__11699\,
            I => \C3_c_g\
        );

    \I__2790\ : CEMux
    port map (
            O => \N__11696\,
            I => \N__11651\
        );

    \I__2789\ : CEMux
    port map (
            O => \N__11695\,
            I => \N__11651\
        );

    \I__2788\ : CEMux
    port map (
            O => \N__11694\,
            I => \N__11651\
        );

    \I__2787\ : CEMux
    port map (
            O => \N__11693\,
            I => \N__11651\
        );

    \I__2786\ : CEMux
    port map (
            O => \N__11692\,
            I => \N__11651\
        );

    \I__2785\ : CEMux
    port map (
            O => \N__11691\,
            I => \N__11651\
        );

    \I__2784\ : CEMux
    port map (
            O => \N__11690\,
            I => \N__11651\
        );

    \I__2783\ : CEMux
    port map (
            O => \N__11689\,
            I => \N__11651\
        );

    \I__2782\ : CEMux
    port map (
            O => \N__11688\,
            I => \N__11651\
        );

    \I__2781\ : CEMux
    port map (
            O => \N__11687\,
            I => \N__11651\
        );

    \I__2780\ : CEMux
    port map (
            O => \N__11686\,
            I => \N__11651\
        );

    \I__2779\ : CEMux
    port map (
            O => \N__11685\,
            I => \N__11651\
        );

    \I__2778\ : CEMux
    port map (
            O => \N__11684\,
            I => \N__11651\
        );

    \I__2777\ : CEMux
    port map (
            O => \N__11683\,
            I => \N__11651\
        );

    \I__2776\ : CEMux
    port map (
            O => \N__11682\,
            I => \N__11651\
        );

    \I__2775\ : GlobalMux
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__2774\ : gio2CtrlBuf
    port map (
            O => \N__11648\,
            I => \DBRn_c_i_0_g\
        );

    \I__2773\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11638\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11635\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11643\,
            I => \N__11632\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11629\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11626\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11612\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11635\,
            I => \N__11587\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__11632\,
            I => \N__11581\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11629\,
            I => \N__11565\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__11626\,
            I => \N__11559\
        );

    \I__2763\ : SRMux
    port map (
            O => \N__11625\,
            I => \N__11435\
        );

    \I__2762\ : SRMux
    port map (
            O => \N__11624\,
            I => \N__11435\
        );

    \I__2761\ : SRMux
    port map (
            O => \N__11623\,
            I => \N__11435\
        );

    \I__2760\ : SRMux
    port map (
            O => \N__11622\,
            I => \N__11435\
        );

    \I__2759\ : SRMux
    port map (
            O => \N__11621\,
            I => \N__11435\
        );

    \I__2758\ : SRMux
    port map (
            O => \N__11620\,
            I => \N__11435\
        );

    \I__2757\ : SRMux
    port map (
            O => \N__11619\,
            I => \N__11435\
        );

    \I__2756\ : SRMux
    port map (
            O => \N__11618\,
            I => \N__11435\
        );

    \I__2755\ : SRMux
    port map (
            O => \N__11617\,
            I => \N__11435\
        );

    \I__2754\ : SRMux
    port map (
            O => \N__11616\,
            I => \N__11435\
        );

    \I__2753\ : SRMux
    port map (
            O => \N__11615\,
            I => \N__11435\
        );

    \I__2752\ : Glb2LocalMux
    port map (
            O => \N__11612\,
            I => \N__11435\
        );

    \I__2751\ : SRMux
    port map (
            O => \N__11611\,
            I => \N__11435\
        );

    \I__2750\ : SRMux
    port map (
            O => \N__11610\,
            I => \N__11435\
        );

    \I__2749\ : SRMux
    port map (
            O => \N__11609\,
            I => \N__11435\
        );

    \I__2748\ : SRMux
    port map (
            O => \N__11608\,
            I => \N__11435\
        );

    \I__2747\ : SRMux
    port map (
            O => \N__11607\,
            I => \N__11435\
        );

    \I__2746\ : SRMux
    port map (
            O => \N__11606\,
            I => \N__11435\
        );

    \I__2745\ : SRMux
    port map (
            O => \N__11605\,
            I => \N__11435\
        );

    \I__2744\ : SRMux
    port map (
            O => \N__11604\,
            I => \N__11435\
        );

    \I__2743\ : SRMux
    port map (
            O => \N__11603\,
            I => \N__11435\
        );

    \I__2742\ : SRMux
    port map (
            O => \N__11602\,
            I => \N__11435\
        );

    \I__2741\ : SRMux
    port map (
            O => \N__11601\,
            I => \N__11435\
        );

    \I__2740\ : SRMux
    port map (
            O => \N__11600\,
            I => \N__11435\
        );

    \I__2739\ : SRMux
    port map (
            O => \N__11599\,
            I => \N__11435\
        );

    \I__2738\ : SRMux
    port map (
            O => \N__11598\,
            I => \N__11435\
        );

    \I__2737\ : SRMux
    port map (
            O => \N__11597\,
            I => \N__11435\
        );

    \I__2736\ : SRMux
    port map (
            O => \N__11596\,
            I => \N__11435\
        );

    \I__2735\ : SRMux
    port map (
            O => \N__11595\,
            I => \N__11435\
        );

    \I__2734\ : SRMux
    port map (
            O => \N__11594\,
            I => \N__11435\
        );

    \I__2733\ : SRMux
    port map (
            O => \N__11593\,
            I => \N__11435\
        );

    \I__2732\ : SRMux
    port map (
            O => \N__11592\,
            I => \N__11435\
        );

    \I__2731\ : SRMux
    port map (
            O => \N__11591\,
            I => \N__11435\
        );

    \I__2730\ : SRMux
    port map (
            O => \N__11590\,
            I => \N__11435\
        );

    \I__2729\ : Glb2LocalMux
    port map (
            O => \N__11587\,
            I => \N__11435\
        );

    \I__2728\ : SRMux
    port map (
            O => \N__11586\,
            I => \N__11435\
        );

    \I__2727\ : SRMux
    port map (
            O => \N__11585\,
            I => \N__11435\
        );

    \I__2726\ : SRMux
    port map (
            O => \N__11584\,
            I => \N__11435\
        );

    \I__2725\ : Glb2LocalMux
    port map (
            O => \N__11581\,
            I => \N__11435\
        );

    \I__2724\ : SRMux
    port map (
            O => \N__11580\,
            I => \N__11435\
        );

    \I__2723\ : SRMux
    port map (
            O => \N__11579\,
            I => \N__11435\
        );

    \I__2722\ : SRMux
    port map (
            O => \N__11578\,
            I => \N__11435\
        );

    \I__2721\ : SRMux
    port map (
            O => \N__11577\,
            I => \N__11435\
        );

    \I__2720\ : SRMux
    port map (
            O => \N__11576\,
            I => \N__11435\
        );

    \I__2719\ : SRMux
    port map (
            O => \N__11575\,
            I => \N__11435\
        );

    \I__2718\ : SRMux
    port map (
            O => \N__11574\,
            I => \N__11435\
        );

    \I__2717\ : SRMux
    port map (
            O => \N__11573\,
            I => \N__11435\
        );

    \I__2716\ : SRMux
    port map (
            O => \N__11572\,
            I => \N__11435\
        );

    \I__2715\ : SRMux
    port map (
            O => \N__11571\,
            I => \N__11435\
        );

    \I__2714\ : SRMux
    port map (
            O => \N__11570\,
            I => \N__11435\
        );

    \I__2713\ : SRMux
    port map (
            O => \N__11569\,
            I => \N__11435\
        );

    \I__2712\ : SRMux
    port map (
            O => \N__11568\,
            I => \N__11435\
        );

    \I__2711\ : Glb2LocalMux
    port map (
            O => \N__11565\,
            I => \N__11435\
        );

    \I__2710\ : SRMux
    port map (
            O => \N__11564\,
            I => \N__11435\
        );

    \I__2709\ : SRMux
    port map (
            O => \N__11563\,
            I => \N__11435\
        );

    \I__2708\ : SRMux
    port map (
            O => \N__11562\,
            I => \N__11435\
        );

    \I__2707\ : Glb2LocalMux
    port map (
            O => \N__11559\,
            I => \N__11435\
        );

    \I__2706\ : SRMux
    port map (
            O => \N__11558\,
            I => \N__11435\
        );

    \I__2705\ : SRMux
    port map (
            O => \N__11557\,
            I => \N__11435\
        );

    \I__2704\ : SRMux
    port map (
            O => \N__11556\,
            I => \N__11435\
        );

    \I__2703\ : GlobalMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__2702\ : gio2CtrlBuf
    port map (
            O => \N__11432\,
            I => \RESETn_c_i_g\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__11429\,
            I => \N__11426\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11421\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11418\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11415\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11421\,
            I => \N__11412\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11418\,
            I => \N__11408\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11415\,
            I => \N__11405\
        );

    \I__2694\ : Span4Mux_v
    port map (
            O => \N__11412\,
            I => \N__11402\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11399\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__11408\,
            I => \N__11395\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__11405\,
            I => \N__11392\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__11402\,
            I => \N__11389\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11386\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11383\
        );

    \I__2687\ : Sp12to4
    port map (
            O => \N__11395\,
            I => \N__11378\
        );

    \I__2686\ : Sp12to4
    port map (
            O => \N__11392\,
            I => \N__11378\
        );

    \I__2685\ : Sp12to4
    port map (
            O => \N__11389\,
            I => \N__11375\
        );

    \I__2684\ : Sp12to4
    port map (
            O => \N__11386\,
            I => \N__11370\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11370\
        );

    \I__2682\ : Span12Mux_h
    port map (
            O => \N__11378\,
            I => \N__11367\
        );

    \I__2681\ : Span12Mux_h
    port map (
            O => \N__11375\,
            I => \N__11362\
        );

    \I__2680\ : Span12Mux_v
    port map (
            O => \N__11370\,
            I => \N__11362\
        );

    \I__2679\ : Span12Mux_v
    port map (
            O => \N__11367\,
            I => \N__11357\
        );

    \I__2678\ : Span12Mux_h
    port map (
            O => \N__11362\,
            I => \N__11357\
        );

    \I__2677\ : Odrv12
    port map (
            O => \N__11357\,
            I => \RnW_c\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11350\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11347\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11344\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__2671\ : Span12Mux_v
    port map (
            O => \N__11341\,
            I => \N__11335\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__11338\,
            I => \N__11332\
        );

    \I__2669\ : Span12Mux_h
    port map (
            O => \N__11335\,
            I => \N__11328\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__11332\,
            I => \N__11325\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11322\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__11328\,
            I => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__11325\,
            I => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11322\,
            I => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\
        );

    \I__2663\ : IoInMux
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__2661\ : IoSpan4Mux
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__2660\ : Span4Mux_s3_h
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__11303\,
            I => \N_323_mux\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__11294\,
            I => \N__11290\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__11290\,
            I => \N__11281\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11287\,
            I => \N__11281\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11276\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__11281\,
            I => \N__11273\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11268\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11268\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11265\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__11273\,
            I => \N__11262\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11259\
        );

    \I__2645\ : Span12Mux_h
    port map (
            O => \N__11265\,
            I => \N__11256\
        );

    \I__2644\ : Sp12to4
    port map (
            O => \N__11262\,
            I => \N__11253\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__11259\,
            I => \N__11250\
        );

    \I__2642\ : Span12Mux_v
    port map (
            O => \N__11256\,
            I => \N__11247\
        );

    \I__2641\ : Span12Mux_h
    port map (
            O => \N__11253\,
            I => \N__11244\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__11250\,
            I => \N__11241\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__11247\,
            I => \CASLn_c\
        );

    \I__2638\ : Odrv12
    port map (
            O => \N__11244\,
            I => \CASLn_c\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__11241\,
            I => \CASLn_c\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11220\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11215\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11223\,
            I => \N__11212\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__11220\,
            I => \N__11209\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11204\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11204\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__11215\,
            I => \N__11199\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11199\
        );

    \I__2625\ : Span4Mux_h
    port map (
            O => \N__11209\,
            I => \N__11194\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__11204\,
            I => \N__11194\
        );

    \I__2623\ : Span12Mux_v
    port map (
            O => \N__11199\,
            I => \N__11191\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__2621\ : Span12Mux_h
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__2619\ : Odrv12
    port map (
            O => \N__11185\,
            I => \CASUn_c\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__11182\,
            I => \CASUn_c\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11171\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__11171\,
            I => \N__11167\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__2609\ : Sp12to4
    port map (
            O => \N__11155\,
            I => \N__11147\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__11152\,
            I => \N__11144\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11139\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11139\
        );

    \I__2605\ : Odrv12
    port map (
            O => \N__11147\,
            I => \REG_CYCLEm\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__11144\,
            I => \REG_CYCLEm\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__11139\,
            I => \REG_CYCLEm\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11126\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__11131\,
            I => \N__11120\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__11130\,
            I => \N__11116\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__11129\,
            I => \N__11109\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11105\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__11125\,
            I => \N__11097\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11090\
        );

    \I__2595\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11085\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11085\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__11119\,
            I => \N__11082\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11077\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11077\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11072\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11072\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11067\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11067\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11062\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__11105\,
            I => \N__11059\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__11104\,
            I => \N__11055\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11052\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__11102\,
            I => \N__11049\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__11101\,
            I => \N__11045\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11041\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11097\,
            I => \N__11038\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11033\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11033\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11028\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11028\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11025\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11022\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11019\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__11077\,
            I => \N__11012\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11012\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11067\,
            I => \N__11012\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11005\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11005\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11005\
        );

    \I__2565\ : Sp12to4
    port map (
            O => \N__11059\,
            I => \N__11002\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \N__10998\
        );

    \I__2563\ : InMux
    port map (
            O => \N__11055\,
            I => \N__10989\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11052\,
            I => \N__10986\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11049\,
            I => \N__10983\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11048\,
            I => \N__10980\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11045\,
            I => \N__10977\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11044\,
            I => \N__10974\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11041\,
            I => \N__10970\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11038\,
            I => \N__10963\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__11033\,
            I => \N__10963\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__11028\,
            I => \N__10963\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__11025\,
            I => \N__10948\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__11022\,
            I => \N__10948\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__10948\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__11012\,
            I => \N__10948\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__11005\,
            I => \N__10948\
        );

    \I__2548\ : Span12Mux_s11_h
    port map (
            O => \N__11002\,
            I => \N__10945\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10942\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10939\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10934\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10934\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10931\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10928\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10925\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10922\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10911\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10986\,
            I => \N__10911\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10911\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10980\,
            I => \N__10911\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10911\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10908\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10905\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__10970\,
            I => \N__10900\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10963\,
            I => \N__10900\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10891\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10891\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10891\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10891\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__10948\,
            I => \N__10888\
        );

    \I__2525\ : Span12Mux_v
    port map (
            O => \N__10945\,
            I => \N__10873\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__10942\,
            I => \N__10873\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10873\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10873\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10873\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10873\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10873\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10922\,
            I => \N__10868\
        );

    \I__2517\ : Span12Mux_h
    port map (
            O => \N__10911\,
            I => \N__10868\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__10908\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10905\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__10900\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10891\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__10888\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2511\ : Odrv12
    port map (
            O => \N__10873\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2510\ : Odrv12
    port map (
            O => \N__10868\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2509\ : IoInMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__2507\ : Span4Mux_s3_v
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__10841\,
            I => \N_333_mux\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10834\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10830\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10834\,
            I => \N__10826\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10823\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10820\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10817\
        );

    \I__2498\ : Span4Mux_h
    port map (
            O => \N__10826\,
            I => \N__10814\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10811\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__10820\,
            I => \N__10806\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10806\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__10814\,
            I => \N__10803\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10798\
        );

    \I__2492\ : Span4Mux_h
    port map (
            O => \N__10806\,
            I => \N__10798\
        );

    \I__2491\ : Sp12to4
    port map (
            O => \N__10803\,
            I => \N__10793\
        );

    \I__2490\ : Sp12to4
    port map (
            O => \N__10798\,
            I => \N__10793\
        );

    \I__2489\ : Span12Mux_v
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__10790\,
            I => \DRA_c_9\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__2485\ : Span4Mux_h
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__10778\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__10769\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__2477\ : Span4Mux_h
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__10754\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10746\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10743\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10749\,
            I => \N__10740\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10736\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10743\,
            I => \N__10731\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10740\,
            I => \N__10731\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10728\
        );

    \I__2468\ : Span4Mux_h
    port map (
            O => \N__10736\,
            I => \N__10725\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__10731\,
            I => \N__10720\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10728\,
            I => \N__10720\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__10725\,
            I => \N__10717\
        );

    \I__2464\ : Sp12to4
    port map (
            O => \N__10720\,
            I => \N__10714\
        );

    \I__2463\ : Sp12to4
    port map (
            O => \N__10717\,
            I => \N__10709\
        );

    \I__2462\ : Span12Mux_v
    port map (
            O => \N__10714\,
            I => \N__10709\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__10709\,
            I => \DRA_c_5\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__10697\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__10688\,
            I => \N__10685\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__10682\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__10667\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__10658\,
            I => \N__10654\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10651\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__10654\,
            I => \N__10646\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10646\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__10646\,
            I => \N__10640\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__10645\,
            I => \N__10637\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10644\,
            I => \N__10634\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10631\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__10640\,
            I => \N__10628\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10625\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10634\,
            I => \N__10622\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10631\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__10628\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10625\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__10622\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2429\ : IoInMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__2427\ : IoSpan4Mux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2426\ : Span4Mux_s3_v
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__10598\,
            I => \CRCSn_c\
        );

    \I__2423\ : IoInMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10592\,
            I => \N__10589\
        );

    \I__2421\ : IoSpan4Mux
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__2420\ : Span4Mux_s2_v
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__10577\,
            I => \CASn_c\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__10574\,
            I => \N__10564\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10561\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10558\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__10571\,
            I => \N__10554\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \N__10550\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10545\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__10568\,
            I => \N__10536\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10531\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10527\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10524\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10521\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10518\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10512\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10512\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10505\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10505\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10505\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10502\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10497\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10497\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10542\,
            I => \N__10492\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10492\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__10540\,
            I => \N__10487\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10484\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10481\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10476\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10476\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10471\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10471\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10462\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10524\,
            I => \N__10462\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__10521\,
            I => \N__10462\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10462\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10457\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10512\,
            I => \N__10452\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10452\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__10502\,
            I => \N__10443\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10497\,
            I => \N__10443\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10492\,
            I => \N__10443\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10436\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10433\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10430\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10484\,
            I => \N__10425\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10425\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10476\,
            I => \N__10418\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10471\,
            I => \N__10418\
        );

    \I__2370\ : Span4Mux_h
    port map (
            O => \N__10462\,
            I => \N__10418\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10415\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10412\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10457\,
            I => \N__10409\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__10452\,
            I => \N__10406\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10401\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10401\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__10443\,
            I => \N__10398\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10393\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10393\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10388\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10388\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10436\,
            I => \N__10385\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10433\,
            I => \N__10374\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10374\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10425\,
            I => \N__10374\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10418\,
            I => \N__10374\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10415\,
            I => \N__10374\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10371\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__10409\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__10406\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10401\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__10398\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10393\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10388\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__10385\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__10374\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__10371\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10349\,
            I => \U712_CHIP_RAM.m158_xx_mm_0_2\
        );

    \I__2340\ : IoInMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__2338\ : Span4Mux_s2_h
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2336\ : Span12Mux_s11_v
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2335\ : Odrv12
    port map (
            O => \N__10331\,
            I => \CMA_c_3\
        );

    \I__2334\ : CEMux
    port map (
            O => \N__10328\,
            I => \N__10322\
        );

    \I__2333\ : CEMux
    port map (
            O => \N__10327\,
            I => \N__10316\
        );

    \I__2332\ : CEMux
    port map (
            O => \N__10326\,
            I => \N__10312\
        );

    \I__2331\ : CEMux
    port map (
            O => \N__10325\,
            I => \N__10309\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10322\,
            I => \N__10306\
        );

    \I__2329\ : CEMux
    port map (
            O => \N__10321\,
            I => \N__10303\
        );

    \I__2328\ : CEMux
    port map (
            O => \N__10320\,
            I => \N__10300\
        );

    \I__2327\ : CEMux
    port map (
            O => \N__10319\,
            I => \N__10297\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10294\
        );

    \I__2325\ : CEMux
    port map (
            O => \N__10315\,
            I => \N__10290\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10312\,
            I => \N__10287\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10309\,
            I => \N__10284\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__10306\,
            I => \N__10279\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10279\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10272\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10272\
        );

    \I__2318\ : Span4Mux_h
    port map (
            O => \N__10294\,
            I => \N__10272\
        );

    \I__2317\ : CEMux
    port map (
            O => \N__10293\,
            I => \N__10269\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10290\,
            I => \N__10266\
        );

    \I__2315\ : Span4Mux_v
    port map (
            O => \N__10287\,
            I => \N__10261\
        );

    \I__2314\ : Span4Mux_h
    port map (
            O => \N__10284\,
            I => \N__10261\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__10279\,
            I => \N__10258\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__10272\,
            I => \N__10255\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10269\,
            I => \U712_CHIP_RAM.N_168_0_0\
        );

    \I__2310\ : Odrv12
    port map (
            O => \N__10266\,
            I => \U712_CHIP_RAM.N_168_0_0\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__10261\,
            I => \U712_CHIP_RAM.N_168_0_0\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__10258\,
            I => \U712_CHIP_RAM.N_168_0_0\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__10255\,
            I => \U712_CHIP_RAM.N_168_0_0\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10238\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10235\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__10242\,
            I => \N__10229\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10221\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10238\,
            I => \N__10218\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10215\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10212\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10205\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10205\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10205\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10198\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10198\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10198\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10193\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10193\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10221\,
            I => \N__10188\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__10218\,
            I => \N__10188\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__10215\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10212\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10205\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__10198\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10193\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__10188\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__2283\ : IoInMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__2281\ : Span4Mux_s2_v
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__10157\,
            I => \CMA_c_10\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10150\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10147\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__10150\,
            I => \N__10140\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10140\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10137\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10134\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__10140\,
            I => \N__10131\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10128\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10134\,
            I => \N__10125\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__10131\,
            I => \N__10122\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__10128\,
            I => \N__10117\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__10125\,
            I => \N__10117\
        );

    \I__2264\ : Span12Mux_h
    port map (
            O => \N__10122\,
            I => \N__10114\
        );

    \I__2263\ : Sp12to4
    port map (
            O => \N__10117\,
            I => \N__10111\
        );

    \I__2262\ : Odrv12
    port map (
            O => \N__10114\,
            I => \DRA_c_8\
        );

    \I__2261\ : Odrv12
    port map (
            O => \N__10111\,
            I => \DRA_c_8\
        );

    \I__2260\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__2258\ : Odrv12
    port map (
            O => \N__10100\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10094\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10088\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__10082\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__2251\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10075\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10072\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__10075\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__10072\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__10055\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10049\,
            I => \U712_CHIP_RAM.m158_xx_mm_0_0\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \N__10042\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \N__10039\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10035\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10029\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10025\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10022\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10017\
        );

    \I__2233\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10012\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10012\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10009\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10006\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10025\,
            I => \N__10003\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__10022\,
            I => \N__10000\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10021\,
            I => \N__9997\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10020\,
            I => \N__9994\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__10017\,
            I => \N__9987\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10012\,
            I => \N__9987\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__10009\,
            I => \N__9987\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9980\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__10003\,
            I => \N__9980\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__10000\,
            I => \N__9980\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9997\,
            I => \U712_CHIP_RAM.m154_a2_0\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9994\,
            I => \U712_CHIP_RAM.m154_a2_0\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__9987\,
            I => \U712_CHIP_RAM.m154_a2_0\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__9980\,
            I => \U712_CHIP_RAM.m154_a2_0\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9965\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9962\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9959\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9956\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9965\,
            I => \N__9953\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9962\,
            I => \N__9946\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9959\,
            I => \N__9946\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9956\,
            I => \N__9946\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9953\,
            I => \N__9943\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__9943\,
            I => \N__9937\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__9940\,
            I => \N__9934\
        );

    \I__2203\ : Sp12to4
    port map (
            O => \N__9937\,
            I => \N__9929\
        );

    \I__2202\ : Sp12to4
    port map (
            O => \N__9934\,
            I => \N__9929\
        );

    \I__2201\ : Odrv12
    port map (
            O => \N__9929\,
            I => \DRA_c_7\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9923\,
            I => \N__9919\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9916\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__9919\,
            I => \N__9909\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9916\,
            I => \N__9909\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9906\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9903\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__9909\,
            I => \N__9898\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9906\,
            I => \N__9898\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9903\,
            I => \N__9895\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__9898\,
            I => \N__9892\
        );

    \I__2189\ : Sp12to4
    port map (
            O => \N__9895\,
            I => \N__9889\
        );

    \I__2188\ : Sp12to4
    port map (
            O => \N__9892\,
            I => \N__9886\
        );

    \I__2187\ : Span12Mux_v
    port map (
            O => \N__9889\,
            I => \N__9883\
        );

    \I__2186\ : Span12Mux_h
    port map (
            O => \N__9886\,
            I => \N__9880\
        );

    \I__2185\ : Odrv12
    port map (
            O => \N__9883\,
            I => \DRA_c_6\
        );

    \I__2184\ : Odrv12
    port map (
            O => \N__9880\,
            I => \DRA_c_6\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__9866\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9860\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9860\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9854\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__2173\ : Span4Mux_h
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__9842\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2169\ : Span4Mux_h
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2168\ : Span4Mux_h
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__9827\,
            I => \U712_CHIP_RAM.m228_0\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9818\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9818\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9818\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9810\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9806\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9813\,
            I => \N__9803\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9810\,
            I => \N__9800\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9797\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9794\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9803\,
            I => \N__9791\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__9800\,
            I => \N__9787\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9784\
        );

    \I__2154\ : Span12Mux_h
    port map (
            O => \N__9794\,
            I => \N__9778\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__9791\,
            I => \N__9775\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9772\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__9787\,
            I => \N__9767\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__9784\,
            I => \N__9767\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9762\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9762\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9759\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__9778\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9775\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9772\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__9767\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9762\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9759\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9743\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9743\,
            I => \N__9739\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__9733\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__9730\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2130\ : Sp12to4
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__2129\ : Span12Mux_h
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__9710\,
            I => \A_c_12\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__9698\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__9689\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9680\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9680\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9680\,
            I => \N__9663\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9660\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9655\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9655\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9652\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9647\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9647\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9642\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9642\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9635\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9635\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9635\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9629\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9626\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9623\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9663\,
            I => \N__9616\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9613\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9602\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9602\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9602\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9602\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9635\,
            I => \N__9602\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9595\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9595\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9595\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9629\,
            I => \N__9590\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9590\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9623\,
            I => \N__9587\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9580\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9580\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9580\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9577\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__9616\,
            I => \N__9570\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__9613\,
            I => \N__9570\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__9602\,
            I => \N__9570\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9595\,
            I => \N__9567\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__9590\,
            I => \N__9560\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__9587\,
            I => \N__9553\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9553\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9553\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__9570\,
            I => \N__9548\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__9567\,
            I => \N__9548\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9545\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9540\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9540\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9537\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__9560\,
            I => \N__9532\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__9553\,
            I => \N__9532\
        );

    \I__2070\ : Span4Mux_h
    port map (
            O => \N__9548\,
            I => \N__9529\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9520\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9540\,
            I => \N__9520\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9537\,
            I => \N__9520\
        );

    \I__2066\ : Sp12to4
    port map (
            O => \N__9532\,
            I => \N__9520\
        );

    \I__2065\ : Sp12to4
    port map (
            O => \N__9529\,
            I => \N__9515\
        );

    \I__2064\ : Span12Mux_h
    port map (
            O => \N__9520\,
            I => \N__9515\
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__9515\,
            I => \RESETn_c\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9505\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9496\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9496\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9496\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9496\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9505\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9496\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__9491\,
            I => \N__9487\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9483\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9478\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9478\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9483\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9478\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9468\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9463\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9463\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9457\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9463\,
            I => \N__9457\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9454\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__9457\,
            I => \N__9451\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9454\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9451\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__2040\ : IoInMux
    port map (
            O => \N__9446\,
            I => \N__9442\
        );

    \I__2039\ : IoInMux
    port map (
            O => \N__9445\,
            I => \N__9438\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9435\
        );

    \I__2037\ : IoInMux
    port map (
            O => \N__9441\,
            I => \N__9432\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9438\,
            I => \N__9429\
        );

    \I__2035\ : IoSpan4Mux
    port map (
            O => \N__9435\,
            I => \N__9426\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9423\
        );

    \I__2033\ : Span4Mux_s3_v
    port map (
            O => \N__9429\,
            I => \N__9420\
        );

    \I__2032\ : IoSpan4Mux
    port map (
            O => \N__9426\,
            I => \N__9417\
        );

    \I__2031\ : Span12Mux_s3_v
    port map (
            O => \N__9423\,
            I => \N__9413\
        );

    \I__2030\ : Sp12to4
    port map (
            O => \N__9420\,
            I => \N__9410\
        );

    \I__2029\ : Span4Mux_s2_h
    port map (
            O => \N__9417\,
            I => \N__9407\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9403\
        );

    \I__2027\ : Span12Mux_h
    port map (
            O => \N__9413\,
            I => \N__9398\
        );

    \I__2026\ : Span12Mux_h
    port map (
            O => \N__9410\,
            I => \N__9398\
        );

    \I__2025\ : Sp12to4
    port map (
            O => \N__9407\,
            I => \N__9395\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__9406\,
            I => \N__9392\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9389\
        );

    \I__2022\ : Span12Mux_v
    port map (
            O => \N__9398\,
            I => \N__9386\
        );

    \I__2021\ : Span12Mux_h
    port map (
            O => \N__9395\,
            I => \N__9383\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9380\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__9389\,
            I => \N__9377\
        );

    \I__2018\ : Odrv12
    port map (
            O => \N__9386\,
            I => \TACK_EN\
        );

    \I__2017\ : Odrv12
    port map (
            O => \N__9383\,
            I => \TACK_EN\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9380\,
            I => \TACK_EN\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__9377\,
            I => \TACK_EN\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9357\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9352\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9342\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9342\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9342\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9335\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__9357\,
            I => \N__9332\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9329\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9326\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9352\,
            I => \N__9323\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9316\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9316\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9316\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9342\,
            I => \N__9313\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9304\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9304\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9304\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9304\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9335\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__9332\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9329\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9326\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__9323\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9316\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__9313\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9304\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__1987\ : IoInMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__1985\ : Span4Mux_s2_v
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1983\ : Span4Mux_v
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__9269\,
            I => \ASn_c\
        );

    \I__1980\ : CEMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9263\,
            I => \U712_REG_SM.N_33_0_0\
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1976\ : IoSpan4Mux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__1975\ : Span4Mux_s3_v
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__9242\,
            I => \DMA_LATCH_EN_c\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9236\,
            I => \U712_CHIP_RAM.m160_xx_mm_0_2\
        );

    \I__1969\ : IoInMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9230\,
            I => \N__9227\
        );

    \I__1967\ : Span12Mux_s1_h
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__1966\ : Span12Mux_h
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__1965\ : Odrv12
    port map (
            O => \N__9221\,
            I => \CMA_c_6\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9215\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9209\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1958\ : Span12Mux_v
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__9194\,
            I => \A_c_14\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9188\,
            I => \U712_CHIP_RAM.m155_0_0\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9179\,
            I => \U712_CHIP_RAM.m155_0_2\
        );

    \I__1950\ : IoInMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9173\,
            I => \N__9169\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__1947\ : Span4Mux_s2_v
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9160\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__9160\,
            I => \N__9154\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__1942\ : Span12Mux_h
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__9151\,
            I => \N_68_0\
        );

    \I__1940\ : Odrv12
    port map (
            O => \N__9148\,
            I => \N_68_0\
        );

    \I__1939\ : IoInMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__1937\ : Span4Mux_s2_h
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__1936\ : Sp12to4
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__1935\ : Span12Mux_v
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1934\ : Span12Mux_h
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__1933\ : Odrv12
    port map (
            O => \N__9125\,
            I => \CUUBEn_c\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9118\
        );

    \I__1931\ : IoInMux
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__1927\ : Span12Mux_s10_v
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__9106\,
            I => \N__9100\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__9103\,
            I => \N_145_0\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__9100\,
            I => \N_145_0\
        );

    \I__1923\ : IoInMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__1921\ : IoSpan4Mux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1920\ : Span4Mux_s2_v
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1919\ : Sp12to4
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1918\ : Span12Mux_v
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__9077\,
            I => \CLLBEn_c\
        );

    \I__1916\ : IoInMux
    port map (
            O => \N__9074\,
            I => \N__9069\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9066\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9063\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9060\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9057\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9054\
        );

    \I__1910\ : Span12Mux_s4_v
    port map (
            O => \N__9060\,
            I => \N__9049\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__9057\,
            I => \N__9046\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__9054\,
            I => \N__9043\
        );

    \I__1907\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9038\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9038\
        );

    \I__1905\ : Span12Mux_v
    port map (
            O => \N__9049\,
            I => \N__9028\
        );

    \I__1904\ : Sp12to4
    port map (
            O => \N__9046\,
            I => \N__9028\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__9043\,
            I => \N__9028\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9038\,
            I => \N__9028\
        );

    \I__1901\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9025\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__9028\,
            I => \DBENn_c\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9025\,
            I => \DBENn_c\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9017\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9013\
        );

    \I__1896\ : IoInMux
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__9007\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__9004\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__9007\,
            I => \N__9001\
        );

    \I__1892\ : Span12Mux_s10_v
    port map (
            O => \N__9004\,
            I => \N__8998\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__9001\,
            I => \N__8995\
        );

    \I__1890\ : Odrv12
    port map (
            O => \N__8998\,
            I => \N_71_0\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__8995\,
            I => \N_71_0\
        );

    \I__1888\ : IoInMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__1886\ : Span4Mux_s2_h
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1885\ : Sp12to4
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1884\ : Span12Mux_v
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__1883\ : Span12Mux_h
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__8972\,
            I => \CUMBEn_c\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8966\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8959\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8953\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8959\,
            I => \N__8950\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__8958\,
            I => \N__8946\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__8957\,
            I => \N__8943\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__8956\,
            I => \N__8940\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8935\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__8950\,
            I => \N__8935\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8928\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8928\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8928\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8925\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__8935\,
            I => \N__8922\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8928\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8925\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__8922\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \U712_CYCLE_TERM.N_36_0_cascade_\
        );

    \I__1862\ : IoInMux
    port map (
            O => \N__8912\,
            I => \N__8908\
        );

    \I__1861\ : IoInMux
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1858\ : Span4Mux_s2_v
    port map (
            O => \N__8902\,
            I => \N__8895\
        );

    \I__1857\ : Span4Mux_s1_h
    port map (
            O => \N__8899\,
            I => \N__8892\
        );

    \I__1856\ : IoInMux
    port map (
            O => \N__8898\,
            I => \N__8889\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__8895\,
            I => \N__8886\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__8892\,
            I => \N__8883\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8889\,
            I => \N__8880\
        );

    \I__1852\ : Sp12to4
    port map (
            O => \N__8886\,
            I => \N__8877\
        );

    \I__1851\ : Sp12to4
    port map (
            O => \N__8883\,
            I => \N__8874\
        );

    \I__1850\ : Span12Mux_s10_v
    port map (
            O => \N__8880\,
            I => \N__8871\
        );

    \I__1849\ : Span12Mux_h
    port map (
            O => \N__8877\,
            I => \N__8868\
        );

    \I__1848\ : Span12Mux_v
    port map (
            O => \N__8874\,
            I => \N__8865\
        );

    \I__1847\ : Span12Mux_h
    port map (
            O => \N__8871\,
            I => \N__8861\
        );

    \I__1846\ : Span12Mux_v
    port map (
            O => \N__8868\,
            I => \N__8856\
        );

    \I__1845\ : Span12Mux_h
    port map (
            O => \N__8865\,
            I => \N__8856\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8853\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__8861\,
            I => \TACK_OUT\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8856\,
            I => \TACK_OUT\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8853\,
            I => \TACK_OUT\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8842\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8834\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8842\,
            I => \N__8831\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8828\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8840\,
            I => \N__8825\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8817\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8817\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8817\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8814\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__8831\,
            I => \N__8809\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8809\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8806\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8803\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8817\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__8814\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__8809\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8806\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8803\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8788\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__8782\,
            I => \DBR_SYNC_i_1\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__8779\,
            I => \DBR_SYNC_i_1\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8770\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8767\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8761\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8761\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8758\
        );

    \I__1811\ : Span4Mux_h
    port map (
            O => \N__8761\,
            I => \N__8755\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8758\,
            I => \N_33_0\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8755\,
            I => \N_33_0\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8745\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8749\,
            I => \N__8741\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8738\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8735\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__8744\,
            I => \N__8732\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8728\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8725\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__8735\,
            I => \N__8722\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8719\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8716\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8728\,
            I => \N__8711\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__8725\,
            I => \N__8711\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__8722\,
            I => \N__8706\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8706\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8716\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__8711\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__8706\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1791\ : IoInMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1789\ : IoSpan4Mux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1788\ : Sp12to4
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1787\ : Span12Mux_s9_v
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__8684\,
            I => \RASn_c\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1780\ : Span12Mux_h
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__8663\,
            I => \A_c_19\
        );

    \I__1778\ : IoInMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1776\ : IoSpan4Mux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1775\ : Span4Mux_s0_h
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1774\ : Sp12to4
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1773\ : Span12Mux_h
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__8642\,
            I => \CMA_c_9\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1769\ : Span4Mux_h
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8627\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8621\,
            I => \U712_CHIP_RAM.m160_xx_mm_0_0\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8613\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8610\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8607\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8613\,
            I => \U712_CHIP_RAM.m164_0\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8610\,
            I => \U712_CHIP_RAM.m164_0\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8607\,
            I => \U712_CHIP_RAM.m164_0\
        );

    \I__1758\ : IoInMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__1756\ : Span4Mux_s2_h
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1755\ : Sp12to4
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1754\ : Span12Mux_s10_v
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1753\ : Span12Mux_h
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__8582\,
            I => \CMA_c_5\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8573\,
            I => \U712_CHIP_RAM.m159_xx_mm_0_2\
        );

    \I__1748\ : IoInMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1746\ : Span4Mux_s3_h
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__1745\ : Sp12to4
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1744\ : Span12Mux_v
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__8555\,
            I => \CMA_c_4\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8546\,
            I => \U712_CHIP_RAM.m161_xx_mm_0_2\
        );

    \I__1739\ : IoInMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1737\ : IoSpan4Mux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1736\ : Span4Mux_s3_h
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1735\ : Sp12to4
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1734\ : Span12Mux_h
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1733\ : Odrv12
    port map (
            O => \N__8525\,
            I => \CMA_c_7\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8518\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8510\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8515\,
            I => \N__8510\
        );

    \I__1728\ : Odrv12
    port map (
            O => \N__8510\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8507\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8501\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8498\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8495\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8486\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8486\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8486\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__8477\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8471\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8459\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8459\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8459\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8450\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8441\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8441\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8435\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8426\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8426\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8420\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \U712_CHIP_RAM.m159_xx_mm_0_0_cascade_\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1692\ : Sp12to4
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__1691\ : Span12Mux_h
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1690\ : Odrv12
    port map (
            O => \N__8396\,
            I => \A_c_15\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8387\,
            I => \U712_CHIP_RAM.m156_xx_mm_0_2\
        );

    \I__1686\ : IoInMux
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1684\ : Span4Mux_s2_v
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1683\ : Sp12to4
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__1682\ : Span12Mux_h
    port map (
            O => \N__8372\,
            I => \N__8369\
        );

    \I__1681\ : Odrv12
    port map (
            O => \N__8369\,
            I => \CMA_c_0\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8363\,
            I => \N__8358\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8355\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__8361\,
            I => \N__8351\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__8358\,
            I => \N__8345\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8355\,
            I => \N__8345\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8342\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8339\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8336\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__8345\,
            I => \N__8333\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8330\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8339\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8336\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__8333\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__8330\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1665\ : IoInMux
    port map (
            O => \N__8321\,
            I => \N__8317\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8311\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8308\
        );

    \I__1661\ : Span12Mux_s4_v
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1659\ : Span12Mux_v
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1658\ : Sp12to4
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__1657\ : Span12Mux_h
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1656\ : Span12Mux_h
    port map (
            O => \N__8296\,
            I => \N__8290\
        );

    \I__1655\ : Odrv12
    port map (
            O => \N__8293\,
            I => \A_c_9\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__8290\,
            I => \A_c_9\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__8285\,
            I => \U712_CHIP_RAM.N_3_0_cascade_\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__8282\,
            I => \N__8279\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8276\,
            I => \U712_CHIP_RAM.m156_xx_mm_0_0\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1647\ : IoSpan4Mux
    port map (
            O => \N__8267\,
            I => \N__8263\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8260\
        );

    \I__1645\ : Span4Mux_s2_v
    port map (
            O => \N__8263\,
            I => \N__8257\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8254\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__8257\,
            I => \N__8251\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__8251\,
            I => \N__8243\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__8248\,
            I => \N__8243\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__8243\,
            I => \N_144_0\
        );

    \I__1638\ : IoInMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1636\ : Span4Mux_s3_h
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1635\ : Sp12to4
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1634\ : Span12Mux_v
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1633\ : Span12Mux_h
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__8222\,
            I => \CLMBEn_c\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8212\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1626\ : Span12Mux_h
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__8203\,
            I => \N__8197\
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__8200\,
            I => \DBRn_c_i\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__8197\,
            I => \DBRn_c_i\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8188\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8185\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8188\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8185\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8172\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8172\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8169\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8177\,
            I => \N__8166\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8172\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8169\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8166\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N_20_0\
        );

    \I__1608\ : IoInMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1606\ : IoSpan4Mux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1605\ : Sp12to4
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__1604\ : Span12Mux_v
    port map (
            O => \N__8138\,
            I => \N__8134\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__8134\,
            I => \PRnW_c\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__8131\,
            I => \PRnW_c\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8117\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__8124\,
            I => \N__8114\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__8123\,
            I => \N__8110\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8101\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8117\,
            I => \N__8101\
        );

    \I__1594\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8098\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \N__8091\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8088\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8085\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8078\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8078\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8078\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__8101\,
            I => \N__8073\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8073\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8068\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8068\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8061\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8061\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8061\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8088\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8085\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8078\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__8073\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8068\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8061\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8045\,
            I => \N__8041\
        );

    \I__1572\ : IoInMux
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1571\ : Span4Mux_s1_v
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1568\ : Span12Mux_s11_v
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__8029\,
            I => \N__8023\
        );

    \I__1566\ : Span12Mux_h
    port map (
            O => \N__8026\,
            I => \N__8020\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__8023\,
            I => \N__8017\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__8020\,
            I => \BLSn_c\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__8017\,
            I => \BLSn_c\
        );

    \I__1562\ : CEMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__8003\,
            I => \U712_REG_SM.N_20_0_0\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7997\,
            I => \N_172_0\
        );

    \I__1556\ : IoInMux
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1554\ : Span12Mux_s1_v
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1553\ : Span12Mux_h
    port map (
            O => \N__7985\,
            I => \N__7981\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7978\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7981\,
            I => \LDSn_c\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7978\,
            I => \LDSn_c\
        );

    \I__1549\ : IoInMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1547\ : Span12Mux_s3_v
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__7964\,
            I => \RESETn_c_i\
        );

    \I__1545\ : IoInMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1543\ : IoSpan4Mux
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__1542\ : IoSpan4Mux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__1541\ : Span4Mux_s2_h
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1540\ : Sp12to4
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1539\ : Span12Mux_h
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1538\ : Odrv12
    port map (
            O => \N__7940\,
            I => \WEn_c\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1535\ : Sp12to4
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1534\ : Span12Mux_v
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1533\ : Span12Mux_h
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1532\ : Odrv12
    port map (
            O => \N__7922\,
            I => \A_c_16\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7916\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \U712_CHIP_RAM.m161_xx_mm_0_0_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1525\ : Sp12to4
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1524\ : Span12Mux_h
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__7895\,
            I => \A_c_13\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1520\ : Span12Mux_v
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__7880\,
            I => \A_c_17\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__7868\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__7865\,
            I => \U712_CHIP_RAM.m162_xx_mm_0_0_cascade_\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__7862\,
            I => \U712_CHIP_RAM.m162_xx_mm_0_2_cascade_\
        );

    \I__1511\ : IoInMux
    port map (
            O => \N__7859\,
            I => \N__7856\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7856\,
            I => \N__7853\
        );

    \I__1509\ : IoSpan4Mux
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1508\ : Span4Mux_s3_h
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1507\ : Span4Mux_v
    port map (
            O => \N__7847\,
            I => \N__7844\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1505\ : Sp12to4
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__7838\,
            I => \CMA_c_8\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7832\,
            I => \U712_CHIP_RAM_m45_0\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7822\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7819\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7822\,
            I => \REG_TACK\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7819\,
            I => \REG_TACK\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7811\,
            I => \U712_REG_SM_REG_TACK_7_0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7797\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7792\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7792\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7785\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7785\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7785\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7797\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7792\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7785\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7770\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7770\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7765\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7765\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7770\,
            I => \U712_REG_SM_STATE_COUNT_3\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7765\,
            I => \U712_REG_SM_STATE_COUNT_3\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N_44_0\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7747\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7743\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7747\,
            I => \N__7740\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7737\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N_175_0\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__7740\,
            I => \N_175_0\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7737\,
            I => \N_175_0\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7726\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7723\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7720\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7717\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__1462\ : Sp12to4
    port map (
            O => \N__7714\,
            I => \N__7706\
        );

    \I__1461\ : Sp12to4
    port map (
            O => \N__7711\,
            I => \N__7706\
        );

    \I__1460\ : Span12Mux_h
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__7703\,
            I => \DBRn_c\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7697\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7697\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1456\ : IoInMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__1454\ : Span12Mux_s8_v
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__7685\,
            I => \CMA_c_1\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7679\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7679\,
            I => \U712_CHIP_RAM.m154_0_2\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7669\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7666\
        );

    \I__1447\ : Span4Mux_h
    port map (
            O => \N__7669\,
            I => \N__7663\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7666\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__7663\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7655\,
            I => \U712_CHIP_RAM.m154_0_0\
        );

    \I__1442\ : IoInMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1440\ : Span4Mux_s0_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__7643\,
            I => \N__7639\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7636\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__7639\,
            I => \N__7633\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7636\,
            I => \N__7630\
        );

    \I__1435\ : Sp12to4
    port map (
            O => \N__7633\,
            I => \N__7627\
        );

    \I__1434\ : Span4Mux_v
    port map (
            O => \N__7630\,
            I => \N__7624\
        );

    \I__1433\ : Span12Mux_h
    port map (
            O => \N__7627\,
            I => \N__7621\
        );

    \I__1432\ : Sp12to4
    port map (
            O => \N__7624\,
            I => \N__7618\
        );

    \I__1431\ : Span12Mux_v
    port map (
            O => \N__7621\,
            I => \N__7613\
        );

    \I__1430\ : Span12Mux_h
    port map (
            O => \N__7618\,
            I => \N__7613\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__7613\,
            I => \A_c_10\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7607\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1426\ : IoInMux
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1424\ : IoSpan4Mux
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__1423\ : Span4Mux_s2_v
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__1422\ : Sp12to4
    port map (
            O => \N__7592\,
            I => \N__7588\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7585\
        );

    \I__1420\ : Span12Mux_s8_v
    port map (
            O => \N__7588\,
            I => \N__7582\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__1418\ : Span12Mux_v
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1417\ : Span12Mux_v
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1416\ : Span12Mux_h
    port map (
            O => \N__7576\,
            I => \N__7570\
        );

    \I__1415\ : Span12Mux_h
    port map (
            O => \N__7573\,
            I => \N__7567\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__7570\,
            I => \A_c_11\
        );

    \I__1413\ : Odrv12
    port map (
            O => \N__7567\,
            I => \A_c_11\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__7553\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__7550\,
            I => \U712_CHIP_RAM.m157_xx_mm_0_0_cascade_\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7544\,
            I => \U712_CHIP_RAM.m157_xx_mm_0_2\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__7535\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7528\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7525\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7522\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7525\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__7522\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7513\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7507\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7510\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__7507\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7498\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7501\,
            I => \N__7495\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7498\,
            I => \U712_REG_SM_STATE_COUNT_2\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7495\,
            I => \U712_REG_SM_STATE_COUNT_2\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7484\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7484\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7484\,
            I => \U712_CHIP_RAM.N_37_0\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N_174_0\
        );

    \I__1383\ : IoInMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1381\ : Span12Mux_s5_v
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1380\ : Span12Mux_h
    port map (
            O => \N__7466\,
            I => \N__7462\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7459\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__7462\,
            I => \UDSn_c\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7459\,
            I => \UDSn_c\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7449\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7446\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7443\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7449\,
            I => \N__7437\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7446\,
            I => \N__7432\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7443\,
            I => \N__7432\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7429\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7426\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__7440\,
            I => \N__7423\
        );

    \I__1367\ : Span4Mux_v
    port map (
            O => \N__7437\,
            I => \N__7414\
        );

    \I__1366\ : Span4Mux_h
    port map (
            O => \N__7432\,
            I => \N__7414\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7414\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7414\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7411\
        );

    \I__1362\ : Span4Mux_h
    port map (
            O => \N__7414\,
            I => \N__7406\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7411\,
            I => \N__7406\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1358\ : Sp12to4
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1357\ : Span12Mux_h
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1356\ : Odrv12
    port map (
            O => \N__7394\,
            I => \SIZ_c_0\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__7391\,
            I => \N__7386\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__7390\,
            I => \N__7383\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7376\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7376\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7376\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7373\
        );

    \I__1349\ : Odrv12
    port map (
            O => \N__7373\,
            I => \U712_CHIP_RAM.N_326_mux\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7359\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7359\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7356\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7353\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7359\,
            I => \N__7346\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7356\,
            I => \N__7346\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7353\,
            I => \N__7346\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1339\ : Sp12to4
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1338\ : Span12Mux_h
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__7337\,
            I => \A_c_1\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7330\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7327\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7330\,
            I => \N__7324\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7321\
        );

    \I__1332\ : Span4Mux_h
    port map (
            O => \N__7324\,
            I => \N__7313\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7321\,
            I => \N__7313\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7310\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7307\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7304\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__7313\,
            I => \N__7300\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7293\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7307\,
            I => \N__7293\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7304\,
            I => \N__7293\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7290\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__7300\,
            I => \N__7287\
        );

    \I__1321\ : Sp12to4
    port map (
            O => \N__7293\,
            I => \N__7282\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7290\,
            I => \N__7282\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__7287\,
            I => \N__7277\
        );

    \I__1318\ : Span12Mux_v
    port map (
            O => \N__7282\,
            I => \N__7277\
        );

    \I__1317\ : Span12Mux_h
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__7274\,
            I => \SIZ_c_1\
        );

    \I__1315\ : IoInMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7264\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7261\
        );

    \I__1312\ : IoSpan4Mux
    port map (
            O => \N__7264\,
            I => \N__7258\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7255\
        );

    \I__1310\ : IoSpan4Mux
    port map (
            O => \N__7258\,
            I => \N__7252\
        );

    \I__1309\ : Span12Mux_h
    port map (
            O => \N__7255\,
            I => \N__7249\
        );

    \I__1308\ : IoSpan4Mux
    port map (
            O => \N__7252\,
            I => \N__7246\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__7249\,
            I => \C1_c\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__7246\,
            I => \C1_c\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__7235\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1302\ : ClkMux
    port map (
            O => \N__7232\,
            I => \N__7228\
        );

    \I__1301\ : ClkMux
    port map (
            O => \N__7231\,
            I => \N__7225\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7228\,
            I => \N__7222\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7219\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__7222\,
            I => \N__7216\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__7219\,
            I => \N__7213\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__7216\,
            I => \N__7210\
        );

    \I__1295\ : Sp12to4
    port map (
            O => \N__7213\,
            I => \N__7206\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__7210\,
            I => \N__7203\
        );

    \I__1293\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7200\
        );

    \I__1292\ : Span12Mux_h
    port map (
            O => \N__7206\,
            I => \N__7197\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__7203\,
            I => \N__7192\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__7200\,
            I => \N__7192\
        );

    \I__1289\ : Span12Mux_v
    port map (
            O => \N__7197\,
            I => \N__7189\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__7189\,
            I => \CLK40_PLL\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__7186\,
            I => \CLK40_PLL\
        );

    \I__1285\ : IoInMux
    port map (
            O => \N__7181\,
            I => \N__7177\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__7180\,
            I => \N__7173\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7177\,
            I => \N__7170\
        );

    \I__1282\ : IoInMux
    port map (
            O => \N__7176\,
            I => \N__7167\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7164\
        );

    \I__1280\ : Span4Mux_s1_v
    port map (
            O => \N__7170\,
            I => \N__7161\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7167\,
            I => \N__7158\
        );

    \I__1278\ : Span12Mux_s1_v
    port map (
            O => \N__7164\,
            I => \N__7155\
        );

    \I__1277\ : Sp12to4
    port map (
            O => \N__7161\,
            I => \N__7152\
        );

    \I__1276\ : Span4Mux_s2_h
    port map (
            O => \N__7158\,
            I => \N__7149\
        );

    \I__1275\ : Span12Mux_h
    port map (
            O => \N__7155\,
            I => \N__7146\
        );

    \I__1274\ : Span12Mux_h
    port map (
            O => \N__7152\,
            I => \N__7143\
        );

    \I__1273\ : Sp12to4
    port map (
            O => \N__7149\,
            I => \N__7140\
        );

    \I__1272\ : Span12Mux_v
    port map (
            O => \N__7146\,
            I => \N__7137\
        );

    \I__1271\ : Span12Mux_v
    port map (
            O => \N__7143\,
            I => \N__7134\
        );

    \I__1270\ : Span12Mux_v
    port map (
            O => \N__7140\,
            I => \N__7131\
        );

    \I__1269\ : Span12Mux_v
    port map (
            O => \N__7137\,
            I => \N__7128\
        );

    \I__1268\ : Span12Mux_v
    port map (
            O => \N__7134\,
            I => \N__7123\
        );

    \I__1267\ : Span12Mux_h
    port map (
            O => \N__7131\,
            I => \N__7123\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__7128\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__7123\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__7118\,
            I => \i66_mux_cascade_\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7112\,
            I => \U712_CHIP_RAM.m40_nsZ0Z_1\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7106\,
            I => \N_10_0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7100\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__7088\,
            I => \U712_REG_SM_STATE_COUNT_7\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7082\,
            I => \U712_CHIP_RAM.N_21_0\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__7079\,
            I => \U712_CHIP_RAM.N_21_0_cascade_\
        );

    \I__1250\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7073\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__7067\,
            I => \U712_CHIP_RAM.N_329\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__7064\,
            I => \N__7058\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7052\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7052\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7049\
        );

    \I__1242\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7044\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7044\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7052\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__7049\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7044\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \N_20_0_cascade_\
        );

    \I__1236\ : SRMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7031\,
            I => \U712_CYCLE_TERM.TACK_RST_0_i\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7025\,
            I => \N__7019\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7019\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7019\,
            I => \U712_REG_SM_STATE_COUNT_5\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7013\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__7010\,
            I => \N_10_0_cascade_\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7004\,
            I => \N__6999\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6996\
        );

    \I__1224\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6992\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__6999\,
            I => \N__6989\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6984\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6984\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6992\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__6989\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6984\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6977\,
            I => \U712_CHIP_RAM.N_84_0_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6968\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6965\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6960\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6960\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6968\,
            I => \U712_REG_SM_STATE_COUNT_0\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6965\,
            I => \U712_REG_SM_STATE_COUNT_0\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6960\,
            I => \U712_REG_SM_STATE_COUNT_0\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6953\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6950\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6947\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6944\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1205\ : ClkMux
    port map (
            O => \N__6941\,
            I => \N__6911\
        );

    \I__1204\ : ClkMux
    port map (
            O => \N__6940\,
            I => \N__6911\
        );

    \I__1203\ : ClkMux
    port map (
            O => \N__6939\,
            I => \N__6911\
        );

    \I__1202\ : ClkMux
    port map (
            O => \N__6938\,
            I => \N__6911\
        );

    \I__1201\ : ClkMux
    port map (
            O => \N__6937\,
            I => \N__6911\
        );

    \I__1200\ : ClkMux
    port map (
            O => \N__6936\,
            I => \N__6911\
        );

    \I__1199\ : ClkMux
    port map (
            O => \N__6935\,
            I => \N__6911\
        );

    \I__1198\ : ClkMux
    port map (
            O => \N__6934\,
            I => \N__6911\
        );

    \I__1197\ : ClkMux
    port map (
            O => \N__6933\,
            I => \N__6911\
        );

    \I__1196\ : ClkMux
    port map (
            O => \N__6932\,
            I => \N__6911\
        );

    \I__1195\ : GlobalMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1194\ : gio2CtrlBuf
    port map (
            O => \N__6908\,
            I => \C1_c_g\
        );

    \I__1193\ : SRMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1191\ : Span4Mux_h
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__6896\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6889\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6889\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6886\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6877\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6874\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6877\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6874\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__6869\,
            I => \N__6865\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6862\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6859\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6862\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6859\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6850\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6847\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6850\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6847\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6838\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6835\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6838\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6835\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6826\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6823\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6826\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6823\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6818\,
            I => \U712_CHIP_RAM.REFRESH5lt7_cascade_\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6811\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6808\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6811\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6808\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__6803\,
            I => \N__6799\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__6802\,
            I => \N__6795\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6791\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6788\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6785\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6782\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6778\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6771\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6771\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6782\,
            I => \N__6771\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6768\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__6778\,
            I => \N__6765\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__6771\,
            I => \N__6762\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6768\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__6765\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__6762\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6752\,
            I => \U712_CHIP_RAM.N_168_0\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6746\,
            I => \N__6742\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__6742\,
            I => \CPU_TACKm\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6739\,
            I => \CPU_TACKm\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__6734\,
            I => \U712_CHIP_RAM.N_66_0_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6727\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6724\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6727\,
            I => \N__6721\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__6721\,
            I => \N__6712\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__6718\,
            I => \N__6712\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__6717\,
            I => \N__6709\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__6712\,
            I => \N__6705\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6702\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6699\
        );

    \I__1125\ : Sp12to4
    port map (
            O => \N__6705\,
            I => \N__6692\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6702\,
            I => \N__6692\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6699\,
            I => \N__6692\
        );

    \I__1122\ : Span12Mux_h
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1121\ : Odrv12
    port map (
            O => \N__6689\,
            I => \A_c_0\
        );

    \I__1120\ : IoInMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1118\ : Span12Mux_s5_v
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1117\ : Odrv12
    port map (
            O => \N__6677\,
            I => \CMA_c_2\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6671\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6668\,
            I => \bfn_11_8_0_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6665\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6659\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6652\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6644\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6640\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6635\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6635\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6632\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6648\,
            I => \N__6629\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6626\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6623\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6620\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__6640\,
            I => \N__6612\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6635\,
            I => \N__6612\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6632\,
            I => \N__6612\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6609\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6606\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__6623\,
            I => \N__6601\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6620\,
            I => \N__6601\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6598\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__6612\,
            I => \N__6595\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__6606\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__6601\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6598\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__6595\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__6578\,
            I => \N__6573\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6568\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6568\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__6573\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1079\ : IoInMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6557\
        );

    \I__1077\ : IoSpan4Mux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1076\ : IoSpan4Mux
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1075\ : Span4Mux_s3_h
    port map (
            O => \N__6551\,
            I => \N__6547\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6544\,
            I => \N__6538\
        );

    \I__1071\ : Sp12to4
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__6538\,
            I => \N__6532\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__6535\,
            I => \N__6527\
        );

    \I__1068\ : Sp12to4
    port map (
            O => \N__6532\,
            I => \N__6527\
        );

    \I__1067\ : Span12Mux_h
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__6524\,
            I => \C3_c\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6518\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__6515\,
            I => \U712_CHIP_RAM.N_28_0_cascade_\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6509\,
            I => \U712_CHIP_RAM.N_16_0\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6506\,
            I => \U712_CHIP_RAM.N_16_0_cascade_\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__6503\,
            I => \N__6489\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6485\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__6501\,
            I => \N__6482\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__6500\,
            I => \N__6478\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6471\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6471\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6471\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6466\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6463\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6459\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6450\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6450\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6450\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6450\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6439\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6434\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6434\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6431\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6471\,
            I => \N__6428\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6425\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6422\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6417\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6417\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6414\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6459\,
            I => \N__6409\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6409\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6404\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6404\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6397\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6397\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6397\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6390\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6390\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6390\
        );

    \I__1025\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6381\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6381\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6381\
        );

    \I__1022\ : Span4Mux_v
    port map (
            O => \N__6428\,
            I => \N__6381\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6425\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__6417\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6414\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__6409\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6404\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6397\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6390\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__6381\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6357\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6361\,
            I => \N__6353\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6350\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6357\,
            I => \N__6347\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6344\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6341\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6338\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__6347\,
            I => \U712_CHIP_RAM.N_111_0\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6344\,
            I => \U712_CHIP_RAM.N_111_0\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6341\,
            I => \U712_CHIP_RAM.N_111_0\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__6338\,
            I => \U712_CHIP_RAM.N_111_0\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6319\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__6328\,
            I => \N__6313\
        );

    \I__999\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6304\
        );

    \I__998\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6304\
        );

    \I__997\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6304\
        );

    \I__996\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6301\
        );

    \I__995\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6296\
        );

    \I__994\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6296\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6292\
        );

    \I__992\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6280\
        );

    \I__991\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6280\
        );

    \I__990\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6280\
        );

    \I__989\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6270\
        );

    \I__988\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6270\
        );

    \I__987\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6270\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6304\,
            I => \N__6264\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6259\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6259\
        );

    \I__983\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6255\
        );

    \I__982\ : Span4Mux_h
    port map (
            O => \N__6292\,
            I => \N__6252\
        );

    \I__981\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6247\
        );

    \I__980\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6247\
        );

    \I__979\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6240\
        );

    \I__978\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6240\
        );

    \I__977\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6240\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__6280\,
            I => \N__6237\
        );

    \I__975\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6230\
        );

    \I__974\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6230\
        );

    \I__973\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6230\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6227\
        );

    \I__971\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6220\
        );

    \I__970\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6220\
        );

    \I__969\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6220\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__6264\,
            I => \N__6217\
        );

    \I__967\ : Span4Mux_h
    port map (
            O => \N__6259\,
            I => \N__6214\
        );

    \I__966\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6211\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6255\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__6252\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6247\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6240\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6230\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__6227\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__6220\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__6217\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6211\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__6188\,
            I => \U712_CHIP_RAM.N_359_cascade_\
        );

    \I__953\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6182\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6177\
        );

    \I__951\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6173\
        );

    \I__950\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6170\
        );

    \I__949\ : Span4Mux_h
    port map (
            O => \N__6177\,
            I => \N__6167\
        );

    \I__948\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6164\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6173\,
            I => \U712_CHIP_RAM.N_130_0\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.N_130_0\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__6167\,
            I => \U712_CHIP_RAM.N_130_0\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6164\,
            I => \U712_CHIP_RAM.N_130_0\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__6155\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__6146\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__6143\,
            I => \U712_CHIP_RAM.N_135_0_cascade_\
        );

    \I__938\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6137\,
            I => \U712_CHIP_RAM.N_125_0\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6134\,
            I => \N__6125\
        );

    \I__935\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6120\
        );

    \I__934\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6117\
        );

    \I__933\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6114\
        );

    \I__932\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6111\
        );

    \I__931\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6105\
        );

    \I__930\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6105\
        );

    \I__929\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6102\
        );

    \I__928\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6098\
        );

    \I__927\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6093\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6120\,
            I => \N__6086\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6086\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6114\,
            I => \N__6086\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6083\
        );

    \I__922\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6077\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__6105\,
            I => \N__6073\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6070\
        );

    \I__919\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6067\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6064\
        );

    \I__917\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6059\
        );

    \I__916\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6059\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6093\,
            I => \N__6052\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__6086\,
            I => \N__6052\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__6083\,
            I => \N__6052\
        );

    \I__912\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6045\
        );

    \I__911\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6045\
        );

    \I__910\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6045\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__6077\,
            I => \N__6042\
        );

    \I__908\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6039\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__6073\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__6070\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6067\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__6064\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__6052\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__6045\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__6042\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6039\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__898\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\
        );

    \I__896\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6011\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3\
        );

    \I__894\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6002\
        );

    \I__893\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5999\
        );

    \I__892\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5996\
        );

    \I__891\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5993\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5990\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5999\,
            I => \U712_CHIP_RAM.N_204_0\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5996\,
            I => \U712_CHIP_RAM.N_204_0\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5993\,
            I => \U712_CHIP_RAM.N_204_0\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__5990\,
            I => \U712_CHIP_RAM.N_204_0\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__5981\,
            I => \U712_CHIP_RAM.N_120_0_cascade_\
        );

    \I__884\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5975\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__882\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.m225_0\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5966\,
            I => \N__5962\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__878\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5949\
        );

    \I__877\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5949\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__5958\,
            I => \N__5944\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5957\,
            I => \N__5941\
        );

    \I__874\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5936\
        );

    \I__873\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5931\
        );

    \I__872\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5931\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5949\,
            I => \N__5928\
        );

    \I__870\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5925\
        );

    \I__869\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5920\
        );

    \I__868\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5917\
        );

    \I__867\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5910\
        );

    \I__866\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5910\
        );

    \I__865\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5910\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5905\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5905\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__5928\,
            I => \N__5900\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5900\
        );

    \I__860\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5895\
        );

    \I__859\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5895\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5920\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5917\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5910\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__5905\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__5900\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5895\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__5882\,
            I => \N__5876\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \N__5870\
        );

    \I__850\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5864\
        );

    \I__849\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5864\
        );

    \I__848\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5858\
        );

    \I__847\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5858\
        );

    \I__846\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5852\
        );

    \I__845\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5852\
        );

    \I__844\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5849\
        );

    \I__843\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5846\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5843\
        );

    \I__841\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5840\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5858\,
            I => \N__5837\
        );

    \I__839\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5834\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5852\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5849\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5846\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5840\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__5837\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5834\,
            I => \U712_CHIP_RAM.N_110_0\
        );

    \I__831\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5816\,
            I => \U712_CHIP_RAM.N_112_0\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5813\,
            I => \U712_CHIP_RAM.N_112_0_cascade_\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5810\,
            I => \N__5806\
        );

    \I__827\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5802\
        );

    \I__826\ : InMux
    port map (
            O => \N__5806\,
            I => \N__5793\
        );

    \I__825\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5790\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5787\
        );

    \I__823\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5780\
        );

    \I__822\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5780\
        );

    \I__821\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5780\
        );

    \I__820\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5775\
        );

    \I__819\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5775\
        );

    \I__818\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5772\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5793\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5787\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5772\,
            I => \U712_CHIP_RAM.N_94_0\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__810\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5749\
        );

    \I__808\ : IoInMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__807\ : Span12Mux_h
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__805\ : Span12Mux_v
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__804\ : IoSpan4Mux
    port map (
            O => \N__5740\,
            I => \N__5734\
        );

    \I__803\ : Odrv12
    port map (
            O => \N__5737\,
            I => \RAMENn_c\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__5734\,
            I => \RAMENn_c\
        );

    \I__801\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5723\
        );

    \I__800\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5720\
        );

    \I__799\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5715\
        );

    \I__798\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5715\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5723\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5720\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5715\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__794\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__792\ : Span4Mux_v
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__791\ : Sp12to4
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__790\ : Span12Mux_h
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__789\ : Span12Mux_v
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__5690\,
            I => \REGSPACEn_c\
        );

    \I__787\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5684\,
            I => \N__5680\
        );

    \I__785\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__784\ : Span4Mux_h
    port map (
            O => \N__5680\,
            I => \N__5672\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5672\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__780\ : Sp12to4
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__779\ : Span12Mux_h
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__778\ : Odrv12
    port map (
            O => \N__5660\,
            I => \TSn_c\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__776\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5648\
        );

    \I__775\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5648\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5648\,
            I => \U712_REG_SM_START_RST\
        );

    \I__773\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5636\
        );

    \I__772\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5636\
        );

    \I__771\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5636\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5629\
        );

    \I__769\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5626\
        );

    \I__768\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5623\
        );

    \I__767\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5620\
        );

    \I__766\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5617\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__5629\,
            I => \U712_CHIP_RAM.N_96_0\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.N_96_0\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5623\,
            I => \U712_CHIP_RAM.N_96_0\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5620\,
            I => \U712_CHIP_RAM.N_96_0\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5617\,
            I => \U712_CHIP_RAM.N_96_0\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5606\,
            I => \U712_CHIP_RAM.m123_0_cascade_\
        );

    \I__759\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5600\,
            I => \U712_CHIP_RAM.N_117_0\
        );

    \I__757\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5593\
        );

    \I__756\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5587\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5584\
        );

    \I__754\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5577\
        );

    \I__753\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5577\
        );

    \I__752\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5577\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__750\ : Odrv12
    port map (
            O => \N__5584\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5577\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5570\,
            I => \N__5566\
        );

    \I__747\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__746\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5552\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5552\
        );

    \I__743\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5545\
        );

    \I__742\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5545\
        );

    \I__741\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5545\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__5552\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5536\
        );

    \I__737\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5530\
        );

    \I__736\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__735\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5527\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5527\,
            I => \U712_CHIP_RAM.m92_0\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__5524\,
            I => \U712_CHIP_RAM.m92_0\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__5519\,
            I => \U712_CHIP_RAM.N_130_0_cascade_\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__5516\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_\
        );

    \I__729\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.m203_ns_1\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__5501\,
            I => \U712_CHIP_RAM.N_363_mux_cascade_\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__723\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__5489\,
            I => \N__5485\
        );

    \I__720\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__5485\,
            I => \U712_CHIP_RAM.m186_0\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5482\,
            I => \U712_CHIP_RAM.m186_0\
        );

    \I__717\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.m141_ns_1\
        );

    \I__715\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5465\
        );

    \I__714\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5465\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5465\,
            I => \U712_CHIP_RAM.N_140_0\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.N_140_0_cascade_\
        );

    \I__711\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5454\
        );

    \I__710\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5451\
        );

    \I__709\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5446\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5454\,
            I => \N__5443\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5451\,
            I => \N__5440\
        );

    \I__706\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5435\
        );

    \I__705\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5435\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5446\,
            I => \U712_CHIP_RAM.N_103_0\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__5443\,
            I => \U712_CHIP_RAM.N_103_0\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__5440\,
            I => \U712_CHIP_RAM.N_103_0\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5435\,
            I => \U712_CHIP_RAM.N_103_0\
        );

    \I__700\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5422\
        );

    \I__699\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5422\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5419\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__696\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5410\
        );

    \I__695\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5407\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5404\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5407\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__5404\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__691\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5395\
        );

    \I__690\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5392\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5395\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5392\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__687\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5383\
        );

    \I__686\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5380\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__683\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5367\
        );

    \I__682\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5367\
        );

    \I__681\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5364\
        );

    \I__680\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5361\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5358\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5364\,
            I => \N__5355\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5361\,
            I => \N__5352\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__5358\,
            I => \N__5349\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__5355\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__5352\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__672\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5337\
        );

    \I__671\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5334\
        );

    \I__670\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5331\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5337\,
            I => \U712_CHIP_RAM.N_188_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5334\,
            I => \U712_CHIP_RAM.N_188_0\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5331\,
            I => \U712_CHIP_RAM.N_188_0\
        );

    \I__666\ : CEMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__5315\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\
        );

    \I__662\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5309\,
            I => \N__5305\
        );

    \I__660\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5302\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__5305\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5302\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__5297\,
            I => \U712_CHIP_RAM.N_358_cascade_\
        );

    \I__656\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5291\,
            I => \U712_CHIP_RAM.m219_0\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__5288\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\
        );

    \I__653\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5282\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__650\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5269\
        );

    \I__648\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5266\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__5269\,
            I => \U712_CHIP_RAM.N_137_0\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5266\,
            I => \U712_CHIP_RAM.N_137_0\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__5261\,
            I => \U712_CHIP_RAM.N_142_0_cascade_\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__642\ : Span4Mux_s1_h
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__641\ : Sp12to4
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__640\ : Span12Mux_v
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__639\ : Span12Mux_h
    port map (
            O => \N__5243\,
            I => \N__5239\
        );

    \I__638\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5236\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__5239\,
            I => \CLK_EN_c\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5236\,
            I => \CLK_EN_c\
        );

    \I__635\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER43\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5225\,
            I => \U712_CHIP_RAM.m207_ns_1_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5219\,
            I => \U712_CHIP_RAM.N_206_0\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__629\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.N_208_0\
        );

    \I__625\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5197\
        );

    \I__624\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5194\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5197\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5194\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__621\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5185\
        );

    \I__620\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5182\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5177\,
            I => \U712_CHIP_RAM.m92_0_cascade_\
        );

    \I__616\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5171\,
            I => \U712_CHIP_RAM.N_190_0\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__5168\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__5165\,
            I => \N__5161\
        );

    \I__612\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5157\
        );

    \I__611\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5152\
        );

    \I__610\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5152\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5157\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__5147\,
            I => \U712_CHIP_RAM.N_222_0_cascade_\
        );

    \I__606\ : CEMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__603\ : CEMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__602\ : Span4Mux_v
    port map (
            O => \N__5134\,
            I => \N__5126\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5131\,
            I => \N__5126\
        );

    \I__600\ : Odrv4
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__599\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5119\
        );

    \I__598\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5111\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5108\
        );

    \I__595\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5102\
        );

    \I__594\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5102\
        );

    \I__593\ : Span4Mux_h
    port map (
            O => \N__5111\,
            I => \N__5099\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__5108\,
            I => \N__5096\
        );

    \I__591\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5093\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__5099\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__5096\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.N_111_0_cascade_\
        );

    \I__585\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5078\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__583\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__5069\,
            I => \U712_CHIP_RAM.m138_0\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \U712_CHIP_RAM.N_352_mux_cascade_\
        );

    \I__579\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5060\,
            I => \U712_CHIP_RAM.N_183_0\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__5057\,
            I => \U712_CHIP_RAM.N_137_0_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U712_CHIP_RAM.N_178_0\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__5048\,
            I => \U712_CHIP_RAM.N_94_0_cascade_\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__5045\,
            I => \U712_CHIP_RAM.N_96_0_cascade_\
        );

    \I__572\ : IoInMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__5039\,
            I => \N__5036\
        );

    \I__570\ : Span12Mux_s7_v
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__569\ : Odrv12
    port map (
            O => \N__5033\,
            I => \VBENn_c\
        );

    \I__568\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5027\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5027\,
            I => \N__5024\
        );

    \I__566\ : Span12Mux_h
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__565\ : Span12Mux_v
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__5018\,
            I => \A_c_2\
        );

    \I__563\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__559\ : Sp12to4
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__5000\,
            I => \A_c_5\
        );

    \I__557\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4982\,
            I => \A_c_6\
        );

    \I__551\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__549\ : Span4Mux_h
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__548\ : Sp12to4
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__547\ : Span12Mux_v
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__4964\,
            I => \A_c_3\
        );

    \I__545\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__543\ : Span12Mux_v
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__4952\,
            I => \A_c_7\
        );

    \I__541\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__538\ : Span4Mux_v
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__537\ : Span4Mux_h
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__4931\,
            I => \A_c_4\
        );

    \I__534\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4907\
        );

    \I__533\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4907\
        );

    \I__532\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4907\
        );

    \I__531\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4907\
        );

    \I__530\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4907\
        );

    \I__529\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4907\
        );

    \I__528\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4902\
        );

    \I__527\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4902\
        );

    \I__526\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4899\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4907\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4902\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4899\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__4892\,
            I => \U712_CHIP_RAM.N_206_0_cascade_\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__4889\,
            I => \U712_CHIP_RAM.N_214_0_cascade_\
        );

    \I__520\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4883\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4880\,
            I => \U712_CHIP_RAM.N_216_0_i_cascade_\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__4877\,
            I => \N__4873\
        );

    \I__516\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4870\
        );

    \I__515\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4867\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4870\,
            I => \N__4864\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4867\,
            I => \U712_CHIP_RAM.N_217_0\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4864\,
            I => \U712_CHIP_RAM.N_217_0\
        );

    \I__511\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4850\
        );

    \I__510\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4841\
        );

    \I__509\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4841\
        );

    \I__508\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4841\
        );

    \I__507\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4841\
        );

    \I__506\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4836\
        );

    \I__505\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4836\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4850\,
            I => \U712_CHIP_RAM.N_216_0_i\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4841\,
            I => \U712_CHIP_RAM.N_216_0_i\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4836\,
            I => \U712_CHIP_RAM.N_216_0_i\
        );

    \I__501\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4823\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \U712_CHIP_RAM.N_195_0_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U712_CHIP_RAM.N_213_0\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__494\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4801\
        );

    \I__492\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4798\
        );

    \I__491\ : Odrv4
    port map (
            O => \N__4801\,
            I => \U712_CHIP_RAM.N_189_0\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4798\,
            I => \U712_CHIP_RAM.N_189_0\
        );

    \I__489\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.N_195_0\
        );

    \I__487\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4783\
        );

    \I__486\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4780\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__483\ : InMux
    port map (
            O => \N__4775\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__482\ : InMux
    port map (
            O => \N__4772\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__481\ : InMux
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__480\ : InMux
    port map (
            O => \N__4766\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__479\ : InMux
    port map (
            O => \N__4763\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__478\ : InMux
    port map (
            O => \N__4760\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__477\ : InMux
    port map (
            O => \N__4757\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__476\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4751\,
            I => \U712_CHIP_RAM.N_233\
        );

    \I__474\ : IoInMux
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__472\ : Span4Mux_s3_v
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__471\ : Span4Mux_v
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__470\ : Span4Mux_v
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__469\ : Span4Mux_v
    port map (
            O => \N__4733\,
            I => \N__4729\
        );

    \I__468\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__4729\,
            I => \DBDIR_c\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4726\,
            I => \DBDIR_c\
        );

    \I__465\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__464\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4715\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__462\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4704\
        );

    \I__460\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4699\
        );

    \I__459\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4699\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__4704\,
            I => \N__4694\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4699\,
            I => \N__4694\
        );

    \I__456\ : Span4Mux_v
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__455\ : Span4Mux_v
    port map (
            O => \N__4691\,
            I => \N__4688\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__453\ : IoSpan4Mux
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__4682\,
            I => \AWEn_c\
        );

    \I__451\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__448\ : Sp12to4
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__447\ : Span12Mux_h
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__4661\,
            I => \A_c_18\
        );

    \I__444\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__442\ : Span4Mux_v
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__441\ : Span4Mux_v
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__440\ : Sp12to4
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__4643\,
            I => \A_c_20\
        );

    \I__438\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\
        );

    \I__436\ : IoInMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__434\ : Span4Mux_s3_v
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__433\ : Sp12to4
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__431\ : Span12Mux_v
    port map (
            O => \N__4619\,
            I => \N__4615\
        );

    \I__430\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4612\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__4615\,
            I => \CONSTANT_ONE_NET\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4612\,
            I => \CONSTANT_ONE_NET\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4607\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \U712_CHIP_RAM.m104_ns_1_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4601\,
            I => \U712_CHIP_RAM.N_105_0_cascade_\
        );

    \I__424\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4595\,
            I => \U712_CHIP_RAM.N_106_0\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4592\,
            I => \U712_CHIP_RAM.N_106_0_cascade_\
        );

    \I__421\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4586\,
            I => \U712_CHIP_RAM.DBENn_8_0\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__417\ : Span4Mux_s2_v
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__416\ : Span4Mux_v
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__4571\,
            I => \CLK80_PLL_i_i\
        );

    \I__414\ : IoInMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__4562\,
            I => \DBRn_c_i_0\
        );

    \I__411\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__409\ : Sp12to4
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__408\ : Span12Mux_v
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__4547\,
            I => \A_c_8\
        );

    \I__406\ : IoInMux
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__404\ : IoSpan4Mux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__403\ : Span4Mux_s2_v
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__402\ : Span4Mux_v
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__401\ : Sp12to4
    port map (
            O => \N__4529\,
            I => \N__4525\
        );

    \I__400\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__399\ : Odrv12
    port map (
            O => \N__4525\,
            I => \LATCH_CLK_c\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4522\,
            I => \LATCH_CLK_c\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__395\ : IoSpan4Mux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__394\ : Span4Mux_s2_v
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__393\ : Sp12to4
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__392\ : Span12Mux_v
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__4499\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__6935\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__6937\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__6940\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__6939\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__6941\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__6933\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__6934\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__6938\
        );

    \INVU712_CYCLE_TERM.TACK_ENC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            I => \N__7231\
        );

    \INVU712_CYCLE_TERM.TACK_OUTC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            I => \N__7232\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__6932\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7271\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7973\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4568\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6563\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8215\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11645\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4559\,
            in1 => \N__4787\,
            in2 => \_gnd_net_\,
            in3 => \N__4920\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12117\,
            ce => 'H',
            sr => \N__11605\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__4528\,
            in1 => \N__9790\,
            in2 => \N__6328\,
            in3 => \N__4640\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12117\,
            ce => 'H',
            sr => \N__11605\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4618\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10995\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6311\,
            lcout => \U712_CHIP_RAM.m138_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4712\,
            in1 => \N__11424\,
            in2 => \_gnd_net_\,
            in3 => \N__6656\,
            lcout => \U712_CHIP_RAM.N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5645\,
            in1 => \N__5374\,
            in2 => \_gnd_net_\,
            in3 => \N__6650\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__6128\,
            in1 => \N__9783\,
            in2 => \N__4607\,
            in3 => \N__4598\,
            lcout => \U712_CHIP_RAM.DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12123\,
            ce => 'H',
            sr => \N__11598\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5644\,
            in1 => \N__6469\,
            in2 => \_gnd_net_\,
            in3 => \N__10679\,
            lcout => \U712_CHIP_RAM.DBENn_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIMF791_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110111111"
        )
    port map (
            in0 => \N__6290\,
            in1 => \N__5114\,
            in2 => \N__5958\,
            in3 => \N__9782\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m104_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JFD6_0_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__5809\,
            in1 => \N__6291\,
            in2 => \N__4604\,
            in3 => \N__5458\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_105_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNINNJKA_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__6651\,
            in1 => \N__6495\,
            in2 => \N__4601\,
            in3 => \N__5643\,
            lcout => \U712_CHIP_RAM.N_106_0\,
            ltout => \U712_CHIP_RAM.N_106_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__9037\,
            in1 => \N__6129\,
            in2 => \N__4592\,
            in3 => \N__4589\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12123\,
            ce => 'H',
            sr => \N__11598\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__5375\,
            in1 => \N__4754\,
            in2 => \N__4877\,
            in3 => \N__5115\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12123\,
            ce => 'H',
            sr => \N__11598\
        );

    \U712_CHIP_RAM.DBDIR_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__4707\,
            in1 => \N__4720\,
            in2 => \_gnd_net_\,
            in3 => \N__4732\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12127\,
            ce => 'H',
            sr => \N__11591\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__4721\,
            in1 => \N__4708\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12127\,
            ce => 'H',
            sr => \N__11591\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4679\,
            in1 => \N__4921\,
            in2 => \_gnd_net_\,
            in3 => \N__7531\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__11606\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__4922\,
            in1 => \N__4658\,
            in2 => \N__11939\,
            in3 => \N__5413\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__11606\
        );

    \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5372\,
            in2 => \_gnd_net_\,
            in3 => \N__5341\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__6798\,
            in2 => \N__5498\,
            in3 => \N__5635\,
            lcout => \U712_CHIP_RAM.N_217_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6124\,
            in1 => \N__6470\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10994\,
            in1 => \N__4786\,
            in2 => \_gnd_net_\,
            in3 => \N__10491\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6324\,
            in2 => \_gnd_net_\,
            in3 => \N__4804\,
            lcout => \U712_CHIP_RAM.N_190_0\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__6462\,
            in2 => \_gnd_net_\,
            in3 => \N__4775\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5164\,
            in2 => \_gnd_net_\,
            in3 => \N__4772\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4856\,
            in1 => \N__5947\,
            in2 => \_gnd_net_\,
            in3 => \N__4769\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4853\,
            in1 => \N__5189\,
            in2 => \_gnd_net_\,
            in3 => \N__4766\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__5596\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__5569\,
            in2 => \_gnd_net_\,
            in3 => \N__4760\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4858\,
            in1 => \N__5201\,
            in2 => \_gnd_net_\,
            in3 => \N__4757\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12118\,
            ce => \N__5144\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIJB9Q7_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5450\,
            in1 => \N__9781\,
            in2 => \N__4811\,
            in3 => \N__6278\,
            lcout => \U712_CHIP_RAM.N_206_0\,
            ltout => \U712_CHIP_RAM.N_206_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOVP2B_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__6279\,
            in1 => \N__6449\,
            in2 => \N__4892\,
            in3 => \N__6185\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_214_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJR1UI_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__9685\,
            in1 => \N__6101\,
            in2 => \N__4889\,
            in3 => \N__4817\,
            lcout => \U712_CHIP_RAM.N_216_0_i\,
            ltout => \U712_CHIP_RAM.N_216_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__4886\,
            in1 => \N__5294\,
            in2 => \N__4880\,
            in3 => \N__4876\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12124\,
            ce => \N__5137\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__9686\,
            in1 => \N__4859\,
            in2 => \N__5216\,
            in3 => \N__4829\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12124\,
            ce => \N__5137\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6277\,
            in1 => \N__5956\,
            in2 => \_gnd_net_\,
            in3 => \N__5869\,
            lcout => \U712_CHIP_RAM.N_195_0\,
            ltout => \U712_CHIP_RAM.N_195_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__6448\,
            in1 => \N__5632\,
            in2 => \N__4820\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_213_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNICSPO4_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5857\,
            in1 => \N__5449\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \U712_CHIP_RAM.N_189_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__6123\,
            in1 => \N__6496\,
            in2 => \_gnd_net_\,
            in3 => \N__4793\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => 'H',
            sr => \N__11578\
        );

    \DBRn_ibuf_RNIBAB_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11170\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11044\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5030\,
            in1 => \N__5399\,
            in2 => \_gnd_net_\,
            in3 => \N__4923\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5015\,
            in1 => \N__5387\,
            in2 => \_gnd_net_\,
            in3 => \N__4926\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4927\,
            in1 => \N__4997\,
            in2 => \_gnd_net_\,
            in3 => \N__7516\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4979\,
            in1 => \N__7672\,
            in2 => \_gnd_net_\,
            in3 => \N__4924\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4928\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__8522\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4949\,
            in1 => \N__5426\,
            in2 => \_gnd_net_\,
            in3 => \N__4925\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \N__11599\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011111111"
        )
    port map (
            in0 => \N__6318\,
            in1 => \N__10973\,
            in2 => \N__6361\,
            in3 => \N__6447\,
            lcout => \U712_CHIP_RAM.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_3_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5939\,
            in2 => \_gnd_net_\,
            in3 => \N__5863\,
            lcout => \U712_CHIP_RAM.N_111_0\,
            ltout => \U712_CHIP_RAM.N_111_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000100000"
        )
    port map (
            in0 => \N__6317\,
            in1 => \N__6445\,
            in2 => \N__5084\,
            in3 => \N__5800\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__6745\,
            in1 => \N__5081\,
            in2 => \N__6134\,
            in3 => \N__5063\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12105\,
            ce => 'H',
            sr => \N__11592\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__5312\,
            in1 => \N__6356\,
            in2 => \N__5957\,
            in3 => \N__5801\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_352_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__6446\,
            in1 => \N__5075\,
            in2 => \N__5066\,
            in3 => \N__5272\,
            lcout => \U712_CHIP_RAM.N_183_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5940\,
            in1 => \N__5123\,
            in2 => \_gnd_net_\,
            in3 => \N__5799\,
            lcout => \U712_CHIP_RAM.N_137_0\,
            ltout => \U712_CHIP_RAM.N_137_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__9809\,
            in1 => \N__6316\,
            in2 => \N__5057\,
            in3 => \N__5457\,
            lcout => \U712_CHIP_RAM.N_178_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5559\,
            in1 => \N__5539\,
            in2 => \N__5165\,
            in3 => \N__5592\,
            lcout => \U712_CHIP_RAM.N_94_0\,
            ltout => \U712_CHIP_RAM.N_94_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_3_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__5924\,
            in1 => \_gnd_net_\,
            in2 => \N__5048\,
            in3 => \N__6258\,
            lcout => \U712_CHIP_RAM.N_96_0\,
            ltout => \U712_CHIP_RAM.N_96_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI50JL4_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6794\,
            in1 => \N__6649\,
            in2 => \N__5045\,
            in3 => \N__5488\,
            lcout => \U712_CHIP_RAM.N_188_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5NRT_7_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5200\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \U712_CHIP_RAM.m92_0\,
            ltout => \U712_CHIP_RAM.m92_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__5591\,
            in2 => \N__5177\,
            in3 => \N__5923\,
            lcout => \U712_CHIP_RAM.N_103_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__6110\,
            in1 => \N__5174\,
            in2 => \N__6500\,
            in3 => \N__5340\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5168\,
            in3 => \N__11644\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5590\,
            in1 => \N__5160\,
            in2 => \N__5540\,
            in3 => \N__5558\,
            lcout => \U712_CHIP_RAM.N_110_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIO7T54_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__6584\,
            in1 => \N__5633\,
            in2 => \N__6802\,
            in3 => \N__5728\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_222_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__6643\,
            in1 => \N__5972\,
            in2 => \N__5147\,
            in3 => \N__6096\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001000100"
        )
    port map (
            in0 => \N__6268\,
            in1 => \N__6176\,
            in2 => \N__5881\,
            in3 => \N__6443\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6267\,
            in2 => \_gnd_net_\,
            in3 => \N__5122\,
            lcout => \U712_CHIP_RAM.N_344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6442\,
            in2 => \_gnd_net_\,
            in3 => \N__6076\,
            lcout => \U712_CHIP_RAM.N_358\,
            ltout => \U712_CHIP_RAM.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5297\,
            in3 => \N__9668\,
            lcout => \U712_CHIP_RAM.m219_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__6269\,
            in1 => \N__5819\,
            in2 => \N__5810\,
            in3 => \N__6444\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6097\,
            in2 => \N__5288\,
            in3 => \N__5285\,
            lcout => \U712_CHIP_RAM.N_117_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001010000"
        )
    port map (
            in0 => \N__5477\,
            in1 => \N__5955\,
            in2 => \N__5279\,
            in3 => \N__6493\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_142_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__6082\,
            in1 => \N__5242\,
            in2 => \N__5261\,
            in3 => \N__5231\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12125\,
            ce => 'H',
            sr => \N__11577\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5471\,
            in1 => \N__6492\,
            in2 => \_gnd_net_\,
            in3 => \N__6295\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111010"
        )
    port map (
            in0 => \N__6360\,
            in1 => \N__5470\,
            in2 => \N__6503\,
            in3 => \N__6288\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m207_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101001000010"
        )
    port map (
            in0 => \N__6494\,
            in1 => \N__6081\,
            in2 => \N__5225\,
            in3 => \N__5222\,
            lcout => \U712_CHIP_RAM.N_208_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110101"
        )
    port map (
            in0 => \N__6488\,
            in1 => \N__11100\,
            in2 => \N__5882\,
            in3 => \N__6289\,
            lcout => \U712_CHIP_RAM.m141_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5954\,
            in2 => \_gnd_net_\,
            in3 => \N__5875\,
            lcout => \U712_CHIP_RAM.N_140_0\,
            ltout => \U712_CHIP_RAM.N_140_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBDIU5_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110111111"
        )
    port map (
            in0 => \N__6080\,
            in1 => \N__6287\,
            in2 => \N__5462\,
            in3 => \N__5459\,
            lcout => \U712_CHIP_RAM.m203_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5425\,
            in1 => \N__10960\,
            in2 => \_gnd_net_\,
            in3 => \N__10450\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10962\,
            in1 => \N__10440\,
            in2 => \_gnd_net_\,
            in3 => \N__5414\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5398\,
            in1 => \N__10961\,
            in2 => \_gnd_net_\,
            in3 => \N__10451\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10959\,
            in1 => \N__10439\,
            in2 => \_gnd_net_\,
            in3 => \N__5386\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5373\,
            in2 => \_gnd_net_\,
            in3 => \N__5342\,
            lcout => \U712_CHIP_RAM.CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12098\,
            ce => \N__5324\,
            sr => \N__11584\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6481\,
            in2 => \_gnd_net_\,
            in3 => \N__5308\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m123_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6131\,
            in1 => \N__5634\,
            in2 => \N__5606\,
            in3 => \N__5874\,
            lcout => \U712_CHIP_RAM.N_125_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111111111"
        )
    port map (
            in0 => \N__6005\,
            in1 => \N__5603\,
            in2 => \N__8749\,
            in3 => \N__9566\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_0_5_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__5948\,
            in2 => \N__5570\,
            in3 => \N__5535\,
            lcout => \U712_CHIP_RAM.N_130_0\,
            ltout => \U712_CHIP_RAM.N_130_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6322\,
            in2 => \N__5519\,
            in3 => \N__5796\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__6323\,
            in1 => \N__6180\,
            in2 => \N__6501\,
            in3 => \N__5873\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_3_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__6326\,
            in1 => \N__5798\,
            in2 => \N__5966\,
            in3 => \N__5880\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIU9G4C_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5978\,
            in2 => \N__5516\,
            in3 => \N__5513\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_363_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VCTI_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111000000"
        )
    port map (
            in0 => \N__5507\,
            in1 => \N__6130\,
            in2 => \N__5501\,
            in3 => \N__6499\,
            lcout => \U712_CHIP_RAM.N_204_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI4OCE_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5726\,
            lcout => \U712_CHIP_RAM.m186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__5727\,
            in1 => \N__6619\,
            in2 => \N__6803\,
            in3 => \N__6577\,
            lcout => \U712_CHIP_RAM.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIK0QU_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6497\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9667\,
            lcout => \U712_CHIP_RAM.m225_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_0_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__6325\,
            in1 => \N__5797\,
            in2 => \N__5965\,
            in3 => \N__5879\,
            lcout => \U712_CHIP_RAM.N_112_0\,
            ltout => \U712_CHIP_RAM.N_112_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__6498\,
            in1 => \N__6327\,
            in2 => \N__5813\,
            in3 => \N__5805\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__5687\,
            in1 => \N__10992\,
            in2 => \N__5759\,
            in3 => \N__5729\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12119\,
            ce => 'H',
            sr => \N__11573\
        );

    \U712_REG_SM.START_RST_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__5653\,
            in1 => \N__7746\,
            in2 => \_gnd_net_\,
            in3 => \N__7061\,
            lcout => \U712_REG_SM_START_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12126\,
            ce => 'H',
            sr => \N__11570\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010001"
        )
    port map (
            in0 => \N__5708\,
            in1 => \N__5683\,
            in2 => \N__5657\,
            in3 => \N__7002\,
            lcout => \U712_REG_SM_REG_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12126\,
            ce => 'H',
            sr => \N__11570\
        );

    \U712_CHIP_RAM.m69_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7441\,
            in1 => \N__6708\,
            in2 => \_gnd_net_\,
            in3 => \N__7318\,
            lcout => \U712_CHIP_RAM.N_326_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8354\,
            in1 => \N__10460\,
            in2 => \N__8744\,
            in3 => \N__10644\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001011"
        )
    port map (
            in0 => \N__8731\,
            in1 => \N__8350\,
            in2 => \N__10645\,
            in3 => \N__10441\,
            lcout => \U712_CHIP_RAM.N_168_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6502\,
            in1 => \N__6781\,
            in2 => \_gnd_net_\,
            in3 => \N__6647\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__6362\,
            in1 => \N__6329\,
            in2 => \N__6188\,
            in3 => \N__6181\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6132\,
            in2 => \N__6155\,
            in3 => \N__6152\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_135_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100111111"
        )
    port map (
            in0 => \N__10442\,
            in1 => \N__9679\,
            in2 => \N__6143\,
            in3 => \N__6008\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111111111"
        )
    port map (
            in0 => \N__6140\,
            in1 => \N__6007\,
            in2 => \N__8361\,
            in3 => \N__9564\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6133\,
            in1 => \N__6020\,
            in2 => \_gnd_net_\,
            in3 => \N__6014\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_120_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111101010111"
        )
    port map (
            in0 => \N__9565\,
            in1 => \N__6006\,
            in2 => \N__5981\,
            in3 => \N__10643\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__9839\,
            in1 => \N__9813\,
            in2 => \N__6648\,
            in3 => \N__8962\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12107\,
            ce => 'H',
            sr => \N__11574\
        );

    \U712_REG_SM.C3_SYNC_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6521\,
            lcout => \U712_REG_SM_C3_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \N__11571\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001110111"
        )
    port map (
            in0 => \N__8963\,
            in1 => \N__8483\,
            in2 => \_gnd_net_\,
            in3 => \N__8846\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \N__11571\
        );

    \U712_REG_SM.C3_SYNC_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \N__11571\
        );

    \U712_CHIP_RAM.m11_e_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6971\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6995\,
            lcout => \U712_CHIP_RAM.N_329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m174_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8096\,
            in1 => \N__9349\,
            in2 => \N__7003\,
            in3 => \N__6972\,
            lcout => \N_175_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m27_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__9351\,
            in1 => \N__7502\,
            in2 => \N__8123\,
            in3 => \N__8841\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_28_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__9678\,
            in1 => \N__6512\,
            in2 => \N__6515\,
            in3 => \N__7063\,
            lcout => \U712_REG_SM_STATE_COUNT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m15_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__9350\,
            in1 => \N__8097\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_16_0\,
            ltout => \U712_CHIP_RAM.N_16_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__9677\,
            in1 => \N__7750\,
            in2 => \N__6506\,
            in3 => \N__7062\,
            lcout => \U712_REG_SM_STATE_COUNT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m65_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__7454\,
            in1 => \N__7320\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_66_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m173_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__11411\,
            in1 => \N__6730\,
            in2 => \N__6734\,
            in3 => \N__9356\,
            lcout => \N_174_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m143_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__7365\,
            in1 => \N__7319\,
            in2 => \N__6717\,
            in3 => \N__7442\,
            lcout => \N_144_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m67_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__7303\,
            in1 => \N__7364\,
            in2 => \N__7440\,
            in3 => \N__6731\,
            lcout => \N_68_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__12347\,
            in1 => \N__10517\,
            in2 => \N__11125\,
            in3 => \N__7547\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12081\,
            ce => \N__10326\,
            sr => \N__11593\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6674\,
            in2 => \_gnd_net_\,
            in3 => \N__6668\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6854\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6881\,
            in2 => \_gnd_net_\,
            in3 => \N__6662\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6893\,
            in2 => \_gnd_net_\,
            in3 => \N__6659\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6868\,
            in2 => \_gnd_net_\,
            in3 => \N__6953\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6815\,
            in2 => \_gnd_net_\,
            in3 => \N__6950\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6830\,
            in2 => \_gnd_net_\,
            in3 => \N__6947\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6842\,
            in2 => \_gnd_net_\,
            in3 => \N__6944\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6936\,
            ce => 'H',
            sr => \N__6905\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__6892\,
            in1 => \N__6880\,
            in2 => \N__6869\,
            in3 => \N__6853\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH5lt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6841\,
            in1 => \N__6829\,
            in2 => \N__6818\,
            in3 => \N__6814\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12086\,
            ce => 'H',
            sr => \N__11579\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11643\,
            in2 => \_gnd_net_\,
            in3 => \N__6755\,
            lcout => \U712_CHIP_RAM.N_168_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_START_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7829\,
            in1 => \N__6749\,
            in2 => \_gnd_net_\,
            in3 => \N__9462\,
            lcout => \U712_CYCLE_TERM.TACK_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12092\,
            ce => 'H',
            sr => \N__7034\
        );

    \U712_CYCLE_TERM.TACK_START_RNO_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9563\,
            in2 => \_gnd_net_\,
            in3 => \N__9416\,
            lcout => \U712_CYCLE_TERM.TACK_RST_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9669\,
            in2 => \_gnd_net_\,
            in3 => \N__7103\,
            lcout => \U712_REG_SM_STATE_COUNT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7016\,
            lcout => \U712_REG_SM_STATE_COUNT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m45_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7024\,
            in2 => \_gnd_net_\,
            in3 => \N__6973\,
            lcout => \U712_CHIP_RAM_m45_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__9670\,
            in1 => \_gnd_net_\,
            in2 => \N__7028\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m9_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8107\,
            in2 => \_gnd_net_\,
            in3 => \N__9362\,
            lcout => \N_10_0\,
            ltout => \N_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__7490\,
            in1 => \N__9675\,
            in2 => \N__7010\,
            in3 => \N__7778\,
            lcout => \U712_REG_SM_STATE_COUNT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m83_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7007\,
            in1 => \N__9363\,
            in2 => \_gnd_net_\,
            in3 => \N__8108\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_84_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111110111011"
        )
    port map (
            in0 => \N__7076\,
            in1 => \N__9674\,
            in2 => \N__6977\,
            in3 => \N__6974\,
            lcout => \U712_REG_SM_STATE_COUNT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m40_ns_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000101"
        )
    port map (
            in0 => \N__11150\,
            in1 => \N__7115\,
            in2 => \N__7808\,
            in3 => \N__7489\,
            lcout => OPEN,
            ltout => \i66_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__9672\,
            in1 => \_gnd_net_\,
            in2 => \N__7118\,
            in3 => \N__11151\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m40_ns_1_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__8177\,
            in1 => \N__8106\,
            in2 => \_gnd_net_\,
            in3 => \N__9361\,
            lcout => \U712_CHIP_RAM.m40_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9673\,
            in1 => \N__7777\,
            in2 => \_gnd_net_\,
            in3 => \N__7109\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m32_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__7057\,
            in1 => \N__9338\,
            in2 => \N__8113\,
            in3 => \N__7800\,
            lcout => \N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__7802\,
            in1 => \N__9676\,
            in2 => \N__7097\,
            in3 => \N__7085\,
            lcout => \U712_REG_SM_STATE_COUNT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m20_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9340\,
            lcout => \U712_CHIP_RAM.N_21_0\,
            ltout => \U712_CHIP_RAM.N_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m30_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__7801\,
            in1 => \_gnd_net_\,
            in2 => \N__7079\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m19_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__7070\,
            in2 => \N__7064\,
            in3 => \N__9339\,
            lcout => \N_20_0\,
            ltout => \N_20_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_ess_RNO_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11642\,
            in1 => \_gnd_net_\,
            in2 => \N__7037\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_20_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m36_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7501\,
            in1 => \N__9341\,
            in2 => \N__8840\,
            in3 => \N__8109\,
            lcout => \U712_CHIP_RAM.N_37_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7241\,
            lcout => \U712_REG_SM_C1_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => 'H',
            sr => \N__11563\
        );

    \U712_REG_SM.UDSn_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__7465\,
            in1 => \N__7481\,
            in2 => \_gnd_net_\,
            in3 => \N__8766\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => 'H',
            sr => \N__11563\
        );

    \U712_CHIP_RAM.m144_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__7452\,
            in1 => \N__7366\,
            in2 => \N__7390\,
            in3 => \N__7333\,
            lcout => \N_145_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m171_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__11398\,
            in1 => \_gnd_net_\,
            in2 => \N__7391\,
            in3 => \N__9355\,
            lcout => \N_172_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m70_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010101100"
        )
    port map (
            in0 => \N__7453\,
            in1 => \N__7389\,
            in2 => \N__7370\,
            in3 => \N__7334\,
            lcout => \N_71_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12129\,
            ce => 'H',
            sr => \N__11557\
        );

    \CLK40_PLL_derived_clock_RNIIOT_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__8616\,
            in1 => \N__12203\,
            in2 => \N__11102\,
            in3 => \N__7682\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12078\,
            ce => \N__10320\,
            sr => \N__11590\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__10038\,
            in1 => \N__7658\,
            in2 => \N__9707\,
            in3 => \N__7610\,
            lcout => \U712_CHIP_RAM.m154_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111111"
        )
    port map (
            in0 => \N__10548\,
            in1 => \N__7676\,
            in2 => \N__11119\,
            in3 => \N__10232\,
            lcout => \U712_CHIP_RAM.m154_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11095\,
            in1 => \N__10549\,
            in2 => \N__10242\,
            in3 => \N__7642\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__7591\,
            in1 => \N__11096\,
            in2 => \N__10570\,
            in3 => \N__10233\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m157_xx_mm_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__7562\,
            in1 => \N__10034\,
            in2 => \N__7550\,
            in3 => \N__10766\,
            lcout => \U712_CHIP_RAM.m157_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__7541\,
            in1 => \N__10020\,
            in2 => \N__8282\,
            in3 => \N__10694\,
            lcout => \U712_CHIP_RAM.m156_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7532\,
            in1 => \N__11093\,
            in2 => \_gnd_net_\,
            in3 => \N__10542\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7517\,
            in1 => \N__11094\,
            in2 => \_gnd_net_\,
            in3 => \N__10541\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__10996\,
            in1 => \N__10234\,
            in2 => \N__10540\,
            in3 => \N__7892\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m162_xx_mm_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__10028\,
            in1 => \N__7877\,
            in2 => \N__7865\,
            in3 => \N__8191\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m162_xx_mm_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__10997\,
            in1 => \N__10106\,
            in2 => \N__7862\,
            in3 => \N__10490\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12085\,
            ce => \N__10293\,
            sr => \N__11572\
        );

    \U712_REG_SM.REG_TACK_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__7814\,
            in1 => \N__7835\,
            in2 => \N__7760\,
            in3 => \N__7825\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12094\,
            ce => 'H',
            sr => \N__11568\
        );

    \U712_CHIP_RAM.m35_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__7803\,
            in1 => \N__7776\,
            in2 => \_gnd_net_\,
            in3 => \N__8178\,
            lcout => \U712_REG_SM_REG_TACK_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m43_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000001000"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__9364\,
            in2 => \N__8124\,
            in3 => \N__7775\,
            lcout => \N_44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__11425\,
            in1 => \N__7751\,
            in2 => \_gnd_net_\,
            in3 => \N__8179\,
            lcout => \U712_REG_SM_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__11562\
        );

    \DBR_SYNC_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__11562\
        );

    \DBR_SYNC_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7700\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__11562\
        );

    \U712_REG_SM.PRnW_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110001011100"
        )
    port map (
            in0 => \N__8180\,
            in1 => \N__8137\,
            in2 => \N__8159\,
            in3 => \N__8126\,
            lcout => \PRnW_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__11562\
        );

    \U712_REG_SM.REGENn_ess_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8125\,
            in2 => \_gnd_net_\,
            in3 => \N__9360\,
            lcout => \BLSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12111\,
            ce => \N__8012\,
            sr => \N__11558\
        );

    \U712_REG_SM.LDSn_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__8000\,
            in1 => \N__7984\,
            in2 => \_gnd_net_\,
            in3 => \N__8774\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12116\,
            ce => 'H',
            sr => \N__11556\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9666\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8366\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12080\,
            ce => 'H',
            sr => \N__11600\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_1_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \U712_CHIP_RAM.m164_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__11065\,
            in1 => \N__10227\,
            in2 => \N__10568\,
            in3 => \N__7937\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m161_xx_mm_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__10032\,
            in1 => \N__7919\,
            in2 => \N__7913\,
            in3 => \N__9695\,
            lcout => \U712_CHIP_RAM.m161_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__10228\,
            in1 => \N__7910\,
            in2 => \N__10571\,
            in3 => \N__11066\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m159_xx_mm_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__8423\,
            in1 => \N__10033\,
            in2 => \N__8417\,
            in3 => \N__9851\,
            lcout => \U712_CHIP_RAM.m159_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__8414\,
            in1 => \N__10226\,
            in2 => \N__11108\,
            in3 => \N__10553\,
            lcout => \U712_CHIP_RAM.m160_xx_mm_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__11735\,
            in1 => \N__11114\,
            in2 => \N__8393\,
            in3 => \N__10544\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12087\,
            ce => \N__10315\,
            sr => \N__11580\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8748\,
            in2 => \_gnd_net_\,
            in3 => \N__8362\,
            lcout => \U712_CHIP_RAM.N_3_0\,
            ltout => \U712_CHIP_RAM.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__8320\,
            in1 => \N__11113\,
            in2 => \N__8285\,
            in3 => \N__10543\,
            lcout => \U712_CHIP_RAM.m156_xx_mm_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__8266\,
            in1 => \N__9746\,
            in2 => \N__11058\,
            in3 => \N__9072\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10993\,
            in2 => \_gnd_net_\,
            in3 => \N__10461\,
            lcout => \U712_CHIP_RAM.m154_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10837\,
            in1 => \N__11924\,
            in2 => \N__8219\,
            in3 => \N__8192\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11575\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__9619\,
            in1 => \N__8504\,
            in2 => \N__8956\,
            in3 => \N__8845\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8431\,
            in2 => \N__8791\,
            in3 => \N__8792\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8464\,
            in2 => \_gnd_net_\,
            in3 => \N__8507\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8491\,
            in2 => \_gnd_net_\,
            in3 => \N__8498\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8446\,
            in2 => \_gnd_net_\,
            in3 => \N__8495\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8447\,
            in1 => \N__8492\,
            in2 => \N__8468\,
            in3 => \N__8432\,
            lcout => \U712_CHIP_RAM.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__9621\,
            in1 => \N__8474\,
            in2 => \N__8958\,
            in3 => \N__8839\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__8837\,
            in1 => \N__9622\,
            in2 => \N__8456\,
            in3 => \N__8949\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__9620\,
            in1 => \N__8438\,
            in2 => \N__8957\,
            in3 => \N__8838\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8824\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11641\,
            in2 => \_gnd_net_\,
            in3 => \N__8773\,
            lcout => \U712_REG_SM.N_33_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8750\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => 'H',
            sr => \N__11619\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8618\,
            in1 => \N__8681\,
            in2 => \N__11103\,
            in3 => \N__10787\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12082\,
            ce => \N__10319\,
            sr => \N__11607\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__8624\,
            in2 => \N__10045\,
            in3 => \N__9218\,
            lcout => \U712_CHIP_RAM.m160_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__8617\,
            in1 => \N__9212\,
            in2 => \N__11131\,
            in3 => \N__9182\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12088\,
            ce => \N__10321\,
            sr => \N__11594\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__10775\,
            in1 => \N__11124\,
            in2 => \N__8579\,
            in3 => \N__10535\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12088\,
            ce => \N__10321\,
            sr => \N__11594\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__10534\,
            in1 => \N__11123\,
            in2 => \N__8552\,
            in3 => \N__9863\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12088\,
            ce => \N__10321\,
            sr => \N__11594\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010101"
        )
    port map (
            in0 => \N__10224\,
            in1 => \N__8521\,
            in2 => \N__11129\,
            in3 => \N__10530\,
            lcout => \U712_CHIP_RAM.m155_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9206\,
            in1 => \N__10225\,
            in2 => \N__10567\,
            in3 => \N__11112\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__10021\,
            in1 => \N__9191\,
            in2 => \N__9185\,
            in3 => \N__9857\,
            lcout => \U712_CHIP_RAM.m155_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__9073\,
            in1 => \N__9742\,
            in2 => \N__9172\,
            in3 => \N__11001\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__9824\,
            in1 => \N__9122\,
            in2 => \N__11130\,
            in3 => \N__9053\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__9052\,
            in1 => \N__9823\,
            in2 => \N__9020\,
            in3 => \N__11115\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__11286\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11224\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => 'H',
            sr => \N__11576\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8969\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => 'H',
            sr => \N__11576\
        );

    \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__9486\,
            in1 => \N__9508\,
            in2 => \_gnd_net_\,
            in3 => \N__9471\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_36_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__9511\,
            in1 => \N__9632\,
            in2 => \N__8915\,
            in3 => \N__8864\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__9633\,
            in1 => \N__9510\,
            in2 => \N__9491\,
            in3 => \N__9472\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9634\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__9512\,
            in1 => \N__9490\,
            in2 => \N__9406\,
            in3 => \N__9473\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            ce => 'H',
            sr => \N__11569\
        );

    \U712_REG_SM.ASn_ess_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12130\,
            ce => \N__9266\,
            sr => \N__11564\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11223\,
            in1 => \N__11293\,
            in2 => \_gnd_net_\,
            in3 => \N__11354\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__9875\,
            in1 => \N__11048\,
            in2 => \N__10574\,
            in3 => \N__9239\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__10328\,
            sr => \N__11615\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9970\,
            in1 => \N__11919\,
            in2 => \_gnd_net_\,
            in3 => \N__10154\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11689\,
            sr => \N__11608\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9926\,
            in1 => \N__11928\,
            in2 => \_gnd_net_\,
            in3 => \N__10750\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11723\,
            ce => \N__11687\,
            sr => \N__11601\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9969\,
            in1 => \N__11929\,
            in2 => \_gnd_net_\,
            in3 => \N__10153\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11723\,
            ce => \N__11687\,
            sr => \N__11601\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9968\,
            in1 => \N__11927\,
            in2 => \_gnd_net_\,
            in3 => \N__9922\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__11684\,
            sr => \N__11595\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10751\,
            in1 => \N__11926\,
            in2 => \_gnd_net_\,
            in3 => \N__9915\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11682\,
            sr => \N__11585\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10091\,
            in2 => \_gnd_net_\,
            in3 => \N__10078\,
            lcout => \U712_CHIP_RAM.m228_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11300\,
            lcout => \U712_CHIP_RAM.N_343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11234\,
            in2 => \_gnd_net_\,
            in3 => \N__9814\,
            lcout => \U712_CHIP_RAM.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__9725\,
            in1 => \N__10244\,
            in2 => \N__11101\,
            in3 => \N__10557\,
            lcout => \U712_CHIP_RAM.m158_xx_mm_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12338\,
            in1 => \N__11918\,
            in2 => \_gnd_net_\,
            in3 => \N__12242\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11692\,
            sr => \N__11616\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10145\,
            in1 => \N__11902\,
            in2 => \_gnd_net_\,
            in3 => \N__10838\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11690\,
            sr => \N__11609\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10243\,
            in1 => \N__10657\,
            in2 => \_gnd_net_\,
            in3 => \N__10569\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12102\,
            ce => \N__10325\,
            sr => \N__11602\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__11894\,
            in2 => \_gnd_net_\,
            in3 => \N__10146\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11718\,
            ce => \N__11685\,
            sr => \N__11596\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12146\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__11586\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10097\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__11586\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10079\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__11586\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10085\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__11586\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__10067\,
            in1 => \N__10052\,
            in2 => \N__10046\,
            in3 => \N__10706\,
            lcout => \U712_CHIP_RAM.m158_xx_mm_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11870\,
            in1 => \N__9971\,
            in2 => \_gnd_net_\,
            in3 => \N__9914\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11722\,
            ce => \N__11694\,
            sr => \N__11620\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10833\,
            in1 => \_gnd_net_\,
            in2 => \N__11923\,
            in3 => \N__12175\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11720\,
            ce => \N__11693\,
            sr => \N__11617\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10749\,
            in1 => \N__11895\,
            in2 => \_gnd_net_\,
            in3 => \N__12302\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11720\,
            ce => \N__11693\,
            sr => \N__11617\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11893\,
            in1 => \N__12301\,
            in2 => \_gnd_net_\,
            in3 => \N__12333\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11691\,
            sr => \N__11610\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12300\,
            in1 => \N__11892\,
            in2 => \_gnd_net_\,
            in3 => \N__10739\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11688\,
            sr => \N__11603\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12238\,
            in1 => \N__11817\,
            in2 => \_gnd_net_\,
            in3 => \N__11764\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11683\,
            sr => \N__11597\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11972\,
            in1 => \N__11816\,
            in2 => \_gnd_net_\,
            in3 => \N__11763\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11683\,
            sr => \N__11597\
        );

    \U712_CHIP_RAM.CRCSn_LC_18_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10664\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12084\,
            ce => 'H',
            sr => \N__11625\
        );

    \U712_CHIP_RAM.CASn_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10573\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12093\,
            ce => 'H',
            sr => \N__11624\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__12251\,
            in1 => \N__10572\,
            in2 => \N__11104\,
            in3 => \N__10352\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12096\,
            ce => \N__10327\,
            sr => \N__11623\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12234\,
            in1 => \N__11869\,
            in2 => \_gnd_net_\,
            in3 => \N__12332\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => \N__11696\,
            sr => \N__11622\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12334\,
            in1 => \_gnd_net_\,
            in2 => \N__11925\,
            in3 => \N__12299\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11719\,
            ce => \N__11695\,
            sr => \N__11621\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11768\,
            in1 => \N__11903\,
            in2 => \_gnd_net_\,
            in3 => \N__12233\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11719\,
            ce => \N__11695\,
            sr => \N__11621\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12188\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12176\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => 'H',
            sr => \N__11618\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12152\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12122\,
            ce => 'H',
            sr => \N__11611\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11971\,
            in1 => \N__11815\,
            in2 => \_gnd_net_\,
            in3 => \N__11754\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11717\,
            ce => \N__11686\,
            sr => \N__11604\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001111111"
        )
    port map (
            in0 => \N__11219\,
            in1 => \N__11280\,
            in2 => \N__11429\,
            in3 => \N__11353\,
            lcout => \N_323_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__11279\,
            in1 => \N__11218\,
            in2 => \N__11177\,
            in3 => \N__11132\,
            lcout => \N_333_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

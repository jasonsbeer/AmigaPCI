// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 19 2024 10:38:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    input C1;

    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9943;
    wire N__9942;
    wire N__9941;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9925;
    wire N__9924;
    wire N__9923;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9907;
    wire N__9906;
    wire N__9905;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9889;
    wire N__9888;
    wire N__9887;
    wire N__9880;
    wire N__9879;
    wire N__9878;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9862;
    wire N__9861;
    wire N__9860;
    wire N__9853;
    wire N__9852;
    wire N__9851;
    wire N__9844;
    wire N__9843;
    wire N__9842;
    wire N__9835;
    wire N__9834;
    wire N__9833;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9808;
    wire N__9807;
    wire N__9806;
    wire N__9799;
    wire N__9798;
    wire N__9797;
    wire N__9790;
    wire N__9789;
    wire N__9788;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9772;
    wire N__9771;
    wire N__9770;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9754;
    wire N__9753;
    wire N__9752;
    wire N__9745;
    wire N__9744;
    wire N__9743;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9718;
    wire N__9717;
    wire N__9716;
    wire N__9709;
    wire N__9708;
    wire N__9707;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9691;
    wire N__9690;
    wire N__9689;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9673;
    wire N__9672;
    wire N__9671;
    wire N__9664;
    wire N__9663;
    wire N__9662;
    wire N__9655;
    wire N__9654;
    wire N__9653;
    wire N__9646;
    wire N__9645;
    wire N__9644;
    wire N__9637;
    wire N__9636;
    wire N__9635;
    wire N__9628;
    wire N__9627;
    wire N__9626;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9601;
    wire N__9600;
    wire N__9599;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9574;
    wire N__9573;
    wire N__9572;
    wire N__9565;
    wire N__9564;
    wire N__9563;
    wire N__9556;
    wire N__9555;
    wire N__9554;
    wire N__9547;
    wire N__9546;
    wire N__9545;
    wire N__9538;
    wire N__9537;
    wire N__9536;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9520;
    wire N__9519;
    wire N__9518;
    wire N__9511;
    wire N__9510;
    wire N__9509;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9475;
    wire N__9474;
    wire N__9473;
    wire N__9466;
    wire N__9465;
    wire N__9464;
    wire N__9457;
    wire N__9456;
    wire N__9455;
    wire N__9448;
    wire N__9447;
    wire N__9446;
    wire N__9439;
    wire N__9438;
    wire N__9437;
    wire N__9430;
    wire N__9429;
    wire N__9428;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9385;
    wire N__9384;
    wire N__9383;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9331;
    wire N__9330;
    wire N__9329;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9286;
    wire N__9285;
    wire N__9284;
    wire N__9277;
    wire N__9276;
    wire N__9275;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9222;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9162;
    wire N__9159;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9154;
    wire N__9153;
    wire N__9152;
    wire N__9151;
    wire N__9150;
    wire N__9149;
    wire N__9148;
    wire N__9147;
    wire N__9146;
    wire N__9145;
    wire N__9142;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9133;
    wire N__9132;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9116;
    wire N__9115;
    wire N__9030;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8983;
    wire N__8982;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8975;
    wire N__8974;
    wire N__8973;
    wire N__8972;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8942;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8932;
    wire N__8931;
    wire N__8930;
    wire N__8929;
    wire N__8928;
    wire N__8927;
    wire N__8924;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8814;
    wire N__8813;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8744;
    wire N__8741;
    wire N__8734;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8719;
    wire N__8714;
    wire N__8711;
    wire N__8704;
    wire N__8701;
    wire N__8696;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8666;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8654;
    wire N__8651;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8639;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8620;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8573;
    wire N__8568;
    wire N__8565;
    wire N__8560;
    wire N__8559;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8539;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8531;
    wire N__8528;
    wire N__8523;
    wire N__8516;
    wire N__8513;
    wire N__8508;
    wire N__8505;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8467;
    wire N__8466;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8441;
    wire N__8438;
    wire N__8431;
    wire N__8424;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8162;
    wire N__8161;
    wire N__8160;
    wire N__8159;
    wire N__8158;
    wire N__8157;
    wire N__8156;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8144;
    wire N__8143;
    wire N__8142;
    wire N__8139;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8112;
    wire N__8105;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8087;
    wire N__8082;
    wire N__8077;
    wire N__8076;
    wire N__8075;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8044;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8026;
    wire N__8023;
    wire N__8016;
    wire N__8009;
    wire N__8004;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7839;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7572;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7560;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7523;
    wire N__7522;
    wire N__7521;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7503;
    wire N__7498;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7474;
    wire N__7473;
    wire N__7470;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7424;
    wire N__7421;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7391;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7377;
    wire N__7374;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7341;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7263;
    wire N__7260;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7143;
    wire N__7142;
    wire N__7141;
    wire N__7138;
    wire N__7133;
    wire N__7130;
    wire N__7125;
    wire N__7116;
    wire N__7115;
    wire N__7114;
    wire N__7109;
    wire N__7106;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7047;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6984;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6952;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6930;
    wire N__6927;
    wire N__6926;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6909;
    wire N__6908;
    wire N__6907;
    wire N__6904;
    wire N__6899;
    wire N__6894;
    wire N__6893;
    wire N__6892;
    wire N__6889;
    wire N__6884;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6860;
    wire N__6857;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6837;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6787;
    wire N__6780;
    wire N__6779;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6768;
    wire N__6767;
    wire N__6766;
    wire N__6759;
    wire N__6756;
    wire N__6751;
    wire N__6744;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6722;
    wire N__6721;
    wire N__6720;
    wire N__6717;
    wire N__6710;
    wire N__6705;
    wire N__6702;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6677;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6476;
    wire N__6475;
    wire N__6472;
    wire N__6467;
    wire N__6462;
    wire N__6459;
    wire N__6458;
    wire N__6455;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6443;
    wire N__6440;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6388;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6260;
    wire N__6259;
    wire N__6258;
    wire N__6255;
    wire N__6252;
    wire N__6247;
    wire N__6240;
    wire N__6237;
    wire N__6236;
    wire N__6235;
    wire N__6228;
    wire N__6225;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6213;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6153;
    wire N__6150;
    wire N__6149;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6132;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6103;
    wire N__6098;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6090;
    wire N__6087;
    wire N__6086;
    wire N__6085;
    wire N__6084;
    wire N__6079;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6054;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6047;
    wire N__6042;
    wire N__6039;
    wire N__6038;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6023;
    wire N__6018;
    wire N__6009;
    wire N__6008;
    wire N__6005;
    wire N__6002;
    wire N__5997;
    wire N__5994;
    wire N__5993;
    wire N__5990;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5943;
    wire N__5938;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5916;
    wire N__5913;
    wire N__5912;
    wire N__5911;
    wire N__5908;
    wire N__5903;
    wire N__5902;
    wire N__5897;
    wire N__5894;
    wire N__5889;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5853;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5828;
    wire N__5827;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5792;
    wire N__5791;
    wire N__5786;
    wire N__5785;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5779;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5757;
    wire N__5752;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5726;
    wire N__5725;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5711;
    wire N__5710;
    wire N__5709;
    wire N__5708;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5700;
    wire N__5699;
    wire N__5696;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5677;
    wire N__5676;
    wire N__5675;
    wire N__5674;
    wire N__5673;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5661;
    wire N__5654;
    wire N__5647;
    wire N__5638;
    wire N__5631;
    wire N__5628;
    wire N__5613;
    wire N__5610;
    wire N__5609;
    wire N__5608;
    wire N__5607;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5599;
    wire N__5594;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5586;
    wire N__5583;
    wire N__5582;
    wire N__5579;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5574;
    wire N__5573;
    wire N__5568;
    wire N__5565;
    wire N__5560;
    wire N__5557;
    wire N__5548;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5520;
    wire N__5519;
    wire N__5518;
    wire N__5515;
    wire N__5514;
    wire N__5511;
    wire N__5510;
    wire N__5509;
    wire N__5506;
    wire N__5505;
    wire N__5504;
    wire N__5503;
    wire N__5502;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5488;
    wire N__5485;
    wire N__5480;
    wire N__5473;
    wire N__5460;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5389;
    wire N__5384;
    wire N__5379;
    wire N__5376;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5289;
    wire N__5286;
    wire N__5277;
    wire N__5274;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5237;
    wire N__5234;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5219;
    wire N__5218;
    wire N__5217;
    wire N__5214;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5199;
    wire N__5194;
    wire N__5187;
    wire N__5186;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5179;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5158;
    wire N__5153;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5105;
    wire N__5102;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4892;
    wire N__4889;
    wire N__4888;
    wire N__4885;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4848;
    wire N__4845;
    wire N__4844;
    wire N__4839;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4788;
    wire N__4787;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4770;
    wire N__4767;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4748;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4730;
    wire N__4729;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4719;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4704;
    wire N__4701;
    wire N__4696;
    wire N__4693;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4674;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4633;
    wire N__4632;
    wire N__4627;
    wire N__4622;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4604;
    wire N__4601;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4582;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4570;
    wire N__4563;
    wire N__4560;
    wire N__4559;
    wire N__4556;
    wire N__4555;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4533;
    wire N__4532;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4512;
    wire N__4509;
    wire N__4508;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4497;
    wire N__4496;
    wire N__4495;
    wire N__4494;
    wire N__4487;
    wire N__4478;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4425;
    wire N__4422;
    wire N__4421;
    wire N__4420;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4392;
    wire N__4391;
    wire N__4390;
    wire N__4385;
    wire N__4382;
    wire N__4377;
    wire N__4374;
    wire N__4373;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4359;
    wire N__4358;
    wire N__4355;
    wire N__4354;
    wire N__4351;
    wire N__4346;
    wire N__4343;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4206;
    wire N__4203;
    wire N__4196;
    wire N__4191;
    wire N__4188;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4130;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4016;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4004;
    wire N__3999;
    wire N__3996;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3977;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3912;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3897;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3873;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3861;
    wire N__3858;
    wire N__3857;
    wire N__3854;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3807;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3779;
    wire N__3778;
    wire N__3777;
    wire N__3774;
    wire N__3767;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3746;
    wire N__3745;
    wire N__3744;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3725;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3662;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire bfn_7_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire TACK_EN_i_ess;
    wire N_888_i;
    wire \U712_BYTE_ENABLE.N_451_cascade_ ;
    wire N_48_i;
    wire SIZ_c_1;
    wire \U712_BYTE_ENABLE.N_352_cascade_ ;
    wire N_49_i;
    wire CLK40_OUT_i_i;
    wire A_c_1;
    wire \U712_BYTE_ENABLE.N_457 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_BYTE_ENABLE.N_455 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_459_cascade_ ;
    wire \U712_BYTE_ENABLE.N_352 ;
    wire N_47_i;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_362_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_362_i_0_en_0 ;
    wire VBENn_c;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_ ;
    wire A_c_16;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ;
    wire DBDIR_c;
    wire DRDDIR_i_0;
    wire DRDENn_c;
    wire \U712_REG_SM.N_343_cascade_ ;
    wire \U712_REG_SM.N_358_cascade_ ;
    wire REG_CYCLEm;
    wire REG_TACK;
    wire \U712_CHIP_RAM.N_563_cascade_ ;
    wire \U712_CHIP_RAM.N_215_cascade_ ;
    wire \U712_CHIP_RAM.N_565 ;
    wire \U712_CHIP_RAM.N_565_cascade_ ;
    wire \U712_CHIP_RAM.N_563 ;
    wire \U712_CHIP_RAM.N_445_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_333_cascade_ ;
    wire \U712_CHIP_RAM.N_564 ;
    wire \U712_CHIP_RAM.N_471_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_447_cascade_ ;
    wire \U712_CHIP_RAM.N_333 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_330_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.N_554_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0 ;
    wire \U712_CHIP_RAM.N_332_cascade_ ;
    wire \U712_CHIP_RAM.N_493 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_351 ;
    wire \U712_CHIP_RAM.N_351_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1 ;
    wire \U712_CHIP_RAM.N_402 ;
    wire \U712_CHIP_RAM.N_341 ;
    wire \U712_CHIP_RAM.N_341_cascade_ ;
    wire \U712_CHIP_RAM.N_560 ;
    wire \U712_CHIP_RAM.N_450_cascade_ ;
    wire \U712_CHIP_RAM.N_326_cascade_ ;
    wire \U712_CHIP_RAM.N_326 ;
    wire DBENn_c;
    wire \U712_CHIP_RAM.N_450 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_450_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_7 ;
    wire \U712_REG_SM.N_338 ;
    wire \U712_REG_SM.N_338_cascade_ ;
    wire \U712_REG_SM.N_354_cascade_ ;
    wire REGSPACEn_c;
    wire CASUn_c;
    wire CASLn_c;
    wire \U712_REG_SM.N_431 ;
    wire \U712_REG_SM.N_358 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_71 ;
    wire CMA_c_2;
    wire CONSTANT_ONE_NET;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.N_369 ;
    wire \U712_CHIP_RAM.N_445 ;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_CHIP_RAM.N_492 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_ ;
    wire \U712_CHIP_RAM.N_331 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire \U712_CHIP_RAM.N_222 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ;
    wire \U712_CHIP_RAM.N_332 ;
    wire \U712_CHIP_RAM.N_346 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0 ;
    wire \U712_CHIP_RAM.N_330 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3 ;
    wire \U712_CHIP_RAM.N_52 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire TSn_c;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire DMA_CYCLEm;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_361 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire DBRn_c;
    wire U712_REG_SM_DBR_SYNC_0;
    wire U712_REG_SM_DBR_SYNC_1;
    wire C1_c;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_347_cascade_ ;
    wire \U712_REG_SM.N_559 ;
    wire \U712_REG_SM.N_559_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire ASn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ;
    wire \U712_REG_SM.N_186_0 ;
    wire \U712_REG_SM.N_348_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_364_cascade_ ;
    wire \U712_REG_SM.N_343 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.N_370 ;
    wire CMA_c_3;
    wire CMA_c_1;
    wire A_c_3;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_368 ;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2 ;
    wire \U712_CHIP_RAM.un1_CMA31_0_i ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.N_374 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_BYTE_ENABLE.N_453 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_451 ;
    wire N_50_i;
    wire \U712_REG_SM.N_354 ;
    wire \U712_REG_SM.N_394 ;
    wire \U712_REG_SM.N_364 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire A_c_0;
    wire \U712_REG_SM.N_395 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_REG_SM.N_348 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_347 ;
    wire \U712_REG_SM.N_433 ;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire RnW_c;
    wire SIZ_c_0;
    wire \U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0 ;
    wire CMA_c_10;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_5_i_0_8 ;
    wire A_c_17;
    wire CMA_c_8;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.N_367_cascade_ ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire A_c_14;
    wire A_c_7;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.N_371 ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire CASn_c;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire RASn_c;
    wire \U712_CHIP_RAM.N_373 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.N_372 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire _gnd_net_;
    wire CLK80_OUT;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3540),
            .RESETB(N__5061),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__9952),
            .DIN(N__9951),
            .DOUT(N__9950),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__9952),
            .PADOUT(N__9951),
            .PADIN(N__9950),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4740),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__9943),
            .DIN(N__9942),
            .DOUT(N__9941),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__9943),
            .PADOUT(N__9942),
            .PADIN(N__9941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__9934),
            .DIN(N__9933),
            .DOUT(N__9932),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__9934),
            .PADOUT(N__9933),
            .PADIN(N__9932),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7890),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__9925),
            .DIN(N__9924),
            .DOUT(N__9923),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__9925),
            .PADOUT(N__9924),
            .PADIN(N__9923),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__9916),
            .DIN(N__9915),
            .DOUT(N__9914),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__9916),
            .PADOUT(N__9915),
            .PADIN(N__9914),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__9907),
            .DIN(N__9906),
            .DOUT(N__9905),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__9907),
            .PADOUT(N__9906),
            .PADIN(N__9905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__9898),
            .DIN(N__9897),
            .DOUT(N__9896),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__9898),
            .PADOUT(N__9897),
            .PADIN(N__9896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__9889),
            .DIN(N__9888),
            .DOUT(N__9887),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__9889),
            .PADOUT(N__9888),
            .PADIN(N__9887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__9880),
            .DIN(N__9879),
            .DOUT(N__9878),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__9880),
            .PADOUT(N__9879),
            .PADIN(N__9878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__9871),
            .DIN(N__9870),
            .DOUT(N__9869),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__9871),
            .PADOUT(N__9870),
            .PADIN(N__9869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__9862),
            .DIN(N__9861),
            .DOUT(N__9860),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__9862),
            .PADOUT(N__9861),
            .PADIN(N__9860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__9853),
            .DIN(N__9852),
            .DOUT(N__9851),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__9853),
            .PADOUT(N__9852),
            .PADIN(N__9851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5330),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__9844),
            .DIN(N__9843),
            .DOUT(N__9842),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__9844),
            .PADOUT(N__9843),
            .PADIN(N__9842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9835),
            .DIN(N__9834),
            .DOUT(N__9833),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9835),
            .PADOUT(N__9834),
            .PADIN(N__9833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__9826),
            .DIN(N__9825),
            .DOUT(N__9824),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__9826),
            .PADOUT(N__9825),
            .PADIN(N__9824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3948),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__9817),
            .DIN(N__9816),
            .DOUT(N__9815),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__9817),
            .PADOUT(N__9816),
            .PADIN(N__9815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__9808),
            .DIN(N__9807),
            .DOUT(N__9806),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__9808),
            .PADOUT(N__9807),
            .PADIN(N__9806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__9799),
            .DIN(N__9798),
            .DOUT(N__9797),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__9799),
            .PADOUT(N__9798),
            .PADIN(N__9797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7173),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__9790),
            .DIN(N__9789),
            .DOUT(N__9788),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__9790),
            .PADOUT(N__9789),
            .PADIN(N__9788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__9781),
            .DIN(N__9780),
            .DOUT(N__9779),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__9781),
            .PADOUT(N__9780),
            .PADIN(N__9779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7812),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__9772),
            .DIN(N__9771),
            .DOUT(N__9770),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__9772),
            .PADOUT(N__9771),
            .PADIN(N__9770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__9763),
            .DIN(N__9762),
            .DOUT(N__9761),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__9763),
            .PADOUT(N__9762),
            .PADIN(N__9761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__9754),
            .DIN(N__9753),
            .DOUT(N__9752),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__9754),
            .PADOUT(N__9753),
            .PADIN(N__9752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__9745),
            .DIN(N__9744),
            .DOUT(N__9743),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__9745),
            .PADOUT(N__9744),
            .PADIN(N__9743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__9736),
            .DIN(N__9735),
            .DOUT(N__9734),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__9736),
            .PADOUT(N__9735),
            .PADIN(N__9734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9727),
            .DIN(N__9726),
            .DOUT(N__9725),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9727),
            .PADOUT(N__9726),
            .PADIN(N__9725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4446),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9718),
            .DIN(N__9717),
            .DOUT(N__9716),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9718),
            .PADOUT(N__9717),
            .PADIN(N__9716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__9709),
            .DIN(N__9708),
            .DOUT(N__9707),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__9709),
            .PADOUT(N__9708),
            .PADIN(N__9707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__9700),
            .DIN(N__9699),
            .DOUT(N__9698),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__9700),
            .PADOUT(N__9699),
            .PADIN(N__9698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__9691),
            .DIN(N__9690),
            .DOUT(N__9689),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__9691),
            .PADOUT(N__9690),
            .PADIN(N__9689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__9682),
            .DIN(N__9681),
            .DOUT(N__9680),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__9682),
            .PADOUT(N__9681),
            .PADIN(N__9680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__9673),
            .DIN(N__9672),
            .DOUT(N__9671),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__9673),
            .PADOUT(N__9672),
            .PADIN(N__9671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7773),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__9664),
            .DIN(N__9663),
            .DOUT(N__9662),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__9664),
            .PADOUT(N__9663),
            .PADIN(N__9662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9655),
            .DIN(N__9654),
            .DOUT(N__9653),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9655),
            .PADOUT(N__9654),
            .PADIN(N__9653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9646),
            .DIN(N__9645),
            .DOUT(N__9644),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9646),
            .PADOUT(N__9645),
            .PADIN(N__9644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9637),
            .DIN(N__9636),
            .DOUT(N__9635),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9637),
            .PADOUT(N__9636),
            .PADIN(N__9635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__9628),
            .DIN(N__9627),
            .DOUT(N__9626),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__9628),
            .PADOUT(N__9627),
            .PADIN(N__9626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3675),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9619),
            .DIN(N__9618),
            .DOUT(N__9617),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9619),
            .PADOUT(N__9618),
            .PADIN(N__9617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6825),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9610),
            .DIN(N__9609),
            .DOUT(N__9608),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9610),
            .PADOUT(N__9609),
            .PADIN(N__9608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9601),
            .DIN(N__9600),
            .DOUT(N__9599),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9601),
            .PADOUT(N__9600),
            .PADIN(N__9599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9592),
            .DIN(N__9591),
            .DOUT(N__9590),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9592),
            .PADOUT(N__9591),
            .PADIN(N__9590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9583),
            .DIN(N__9582),
            .DOUT(N__9581),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9583),
            .PADOUT(N__9582),
            .PADIN(N__9581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9574),
            .DIN(N__9573),
            .DOUT(N__9572),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9574),
            .PADOUT(N__9573),
            .PADIN(N__9572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9565),
            .DIN(N__9564),
            .DOUT(N__9563),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9565),
            .PADOUT(N__9564),
            .PADIN(N__9563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9556),
            .DIN(N__9555),
            .DOUT(N__9554),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9556),
            .PADOUT(N__9555),
            .PADIN(N__9554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9547),
            .DIN(N__9546),
            .DOUT(N__9545),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9547),
            .PADOUT(N__9546),
            .PADIN(N__9545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6360),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9538),
            .DIN(N__9537),
            .DOUT(N__9536),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9538),
            .PADOUT(N__9537),
            .PADIN(N__9536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9529),
            .DIN(N__9528),
            .DOUT(N__9527),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9529),
            .PADOUT(N__9528),
            .PADIN(N__9527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9520),
            .DIN(N__9519),
            .DOUT(N__9518),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9520),
            .PADOUT(N__9519),
            .PADIN(N__9518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9511),
            .DIN(N__9510),
            .DOUT(N__9509),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9511),
            .PADOUT(N__9510),
            .PADIN(N__9509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7323),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9502),
            .DIN(N__9501),
            .DOUT(N__9500),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9502),
            .PADOUT(N__9501),
            .PADIN(N__9500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9493),
            .DIN(N__9492),
            .DOUT(N__9491),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9493),
            .PADOUT(N__9492),
            .PADIN(N__9491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7302),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9484),
            .DIN(N__9483),
            .DOUT(N__9482),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9484),
            .PADOUT(N__9483),
            .PADIN(N__9482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9475),
            .DIN(N__9474),
            .DOUT(N__9473),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9475),
            .PADOUT(N__9474),
            .PADIN(N__9473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9466),
            .DIN(N__9465),
            .DOUT(N__9464),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9466),
            .PADOUT(N__9465),
            .PADIN(N__9464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9457),
            .DIN(N__9456),
            .DOUT(N__9455),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9457),
            .PADOUT(N__9456),
            .PADIN(N__9455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6212),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9448),
            .DIN(N__9447),
            .DOUT(N__9446),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9448),
            .PADOUT(N__9447),
            .PADIN(N__9446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9439),
            .DIN(N__9438),
            .DOUT(N__9437),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9439),
            .PADOUT(N__9438),
            .PADIN(N__9437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9430),
            .DIN(N__9429),
            .DOUT(N__9428),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9430),
            .PADOUT(N__9429),
            .PADIN(N__9428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9421),
            .DIN(N__9420),
            .DOUT(N__9419),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9421),
            .PADOUT(N__9420),
            .PADIN(N__9419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9412),
            .DIN(N__9411),
            .DOUT(N__9410),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9412),
            .PADOUT(N__9411),
            .PADIN(N__9410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9403),
            .DIN(N__9402),
            .DOUT(N__9401),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9403),
            .PADOUT(N__9402),
            .PADIN(N__9401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3699),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9394),
            .DIN(N__9393),
            .DOUT(N__9392),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9394),
            .PADOUT(N__9393),
            .PADIN(N__9392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9385),
            .DIN(N__9384),
            .DOUT(N__9383),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9385),
            .PADOUT(N__9384),
            .PADIN(N__9383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9376),
            .DIN(N__9375),
            .DOUT(N__9374),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9376),
            .PADOUT(N__9375),
            .PADIN(N__9374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9367),
            .DIN(N__9366),
            .DOUT(N__9365),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9367),
            .PADOUT(N__9366),
            .PADIN(N__9365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9358),
            .DIN(N__9357),
            .DOUT(N__9356),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9358),
            .PADOUT(N__9357),
            .PADIN(N__9356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6336),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9349),
            .DIN(N__9348),
            .DOUT(N__9347),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9349),
            .PADOUT(N__9348),
            .PADIN(N__9347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9340),
            .DIN(N__9339),
            .DOUT(N__9338),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9340),
            .PADOUT(N__9339),
            .PADIN(N__9338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7023),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9331),
            .DIN(N__9330),
            .DOUT(N__9329),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9331),
            .PADOUT(N__9330),
            .PADIN(N__9329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3606),
            .DIN0(),
            .DOUT0(N__3837),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9322),
            .DIN(N__9321),
            .DOUT(N__9320),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9322),
            .PADOUT(N__9321),
            .PADIN(N__9320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9313),
            .DIN(N__9312),
            .DOUT(N__9311),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9313),
            .PADOUT(N__9312),
            .PADIN(N__9311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9304),
            .DIN(N__9303),
            .DOUT(N__9302),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9304),
            .PADOUT(N__9303),
            .PADIN(N__9302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9295),
            .DIN(N__9294),
            .DOUT(N__9293),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9295),
            .PADOUT(N__9294),
            .PADIN(N__9293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9286),
            .DIN(N__9285),
            .DOUT(N__9284),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9286),
            .PADOUT(N__9285),
            .PADIN(N__9284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9277),
            .DIN(N__9276),
            .DOUT(N__9275),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9277),
            .PADOUT(N__9276),
            .PADIN(N__9275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9268),
            .DIN(N__9267),
            .DOUT(N__9266),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9268),
            .PADOUT(N__9267),
            .PADIN(N__9266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9259),
            .DIN(N__9258),
            .DOUT(N__9257),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9259),
            .PADOUT(N__9258),
            .PADIN(N__9257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9250),
            .DIN(N__9249),
            .DOUT(N__9248),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9250),
            .PADOUT(N__9249),
            .PADIN(N__9248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8490),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9241),
            .DIN(N__9240),
            .DOUT(N__9239),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9241),
            .PADOUT(N__9240),
            .PADIN(N__9239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2198 (
            .O(N__9222),
            .I(N__9218));
    InMux I__2197 (
            .O(N__9221),
            .I(N__9215));
    LocalMux I__2196 (
            .O(N__9218),
            .I(N__9212));
    LocalMux I__2195 (
            .O(N__9215),
            .I(N__9209));
    Span4Mux_v I__2194 (
            .O(N__9212),
            .I(N__9206));
    Span12Mux_v I__2193 (
            .O(N__9209),
            .I(N__9203));
    Span4Mux_h I__2192 (
            .O(N__9206),
            .I(N__9200));
    Span12Mux_h I__2191 (
            .O(N__9203),
            .I(N__9197));
    Span4Mux_h I__2190 (
            .O(N__9200),
            .I(N__9194));
    Odrv12 I__2189 (
            .O(N__9197),
            .I(RAS0n_c));
    Odrv4 I__2188 (
            .O(N__9194),
            .I(RAS0n_c));
    InMux I__2187 (
            .O(N__9189),
            .I(N__9186));
    LocalMux I__2186 (
            .O(N__9186),
            .I(N__9183));
    Span4Mux_v I__2185 (
            .O(N__9183),
            .I(N__9180));
    Sp12to4 I__2184 (
            .O(N__9180),
            .I(N__9177));
    Odrv12 I__2183 (
            .O(N__9177),
            .I(RAS1n_c));
    InMux I__2182 (
            .O(N__9174),
            .I(N__9170));
    InMux I__2181 (
            .O(N__9173),
            .I(N__9167));
    LocalMux I__2180 (
            .O(N__9170),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    LocalMux I__2179 (
            .O(N__9167),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2178 (
            .O(N__9162),
            .I(N__9159));
    LocalMux I__2177 (
            .O(N__9159),
            .I(N__9142));
    ClkMux I__2176 (
            .O(N__9158),
            .I(N__9030));
    ClkMux I__2175 (
            .O(N__9157),
            .I(N__9030));
    ClkMux I__2174 (
            .O(N__9156),
            .I(N__9030));
    ClkMux I__2173 (
            .O(N__9155),
            .I(N__9030));
    ClkMux I__2172 (
            .O(N__9154),
            .I(N__9030));
    ClkMux I__2171 (
            .O(N__9153),
            .I(N__9030));
    ClkMux I__2170 (
            .O(N__9152),
            .I(N__9030));
    ClkMux I__2169 (
            .O(N__9151),
            .I(N__9030));
    ClkMux I__2168 (
            .O(N__9150),
            .I(N__9030));
    ClkMux I__2167 (
            .O(N__9149),
            .I(N__9030));
    ClkMux I__2166 (
            .O(N__9148),
            .I(N__9030));
    ClkMux I__2165 (
            .O(N__9147),
            .I(N__9030));
    ClkMux I__2164 (
            .O(N__9146),
            .I(N__9030));
    ClkMux I__2163 (
            .O(N__9145),
            .I(N__9030));
    Glb2LocalMux I__2162 (
            .O(N__9142),
            .I(N__9030));
    ClkMux I__2161 (
            .O(N__9141),
            .I(N__9030));
    ClkMux I__2160 (
            .O(N__9140),
            .I(N__9030));
    ClkMux I__2159 (
            .O(N__9139),
            .I(N__9030));
    ClkMux I__2158 (
            .O(N__9138),
            .I(N__9030));
    ClkMux I__2157 (
            .O(N__9137),
            .I(N__9030));
    ClkMux I__2156 (
            .O(N__9136),
            .I(N__9030));
    ClkMux I__2155 (
            .O(N__9135),
            .I(N__9030));
    ClkMux I__2154 (
            .O(N__9134),
            .I(N__9030));
    ClkMux I__2153 (
            .O(N__9133),
            .I(N__9030));
    ClkMux I__2152 (
            .O(N__9132),
            .I(N__9030));
    ClkMux I__2151 (
            .O(N__9131),
            .I(N__9030));
    ClkMux I__2150 (
            .O(N__9130),
            .I(N__9030));
    ClkMux I__2149 (
            .O(N__9129),
            .I(N__9030));
    ClkMux I__2148 (
            .O(N__9128),
            .I(N__9030));
    ClkMux I__2147 (
            .O(N__9127),
            .I(N__9030));
    ClkMux I__2146 (
            .O(N__9126),
            .I(N__9030));
    ClkMux I__2145 (
            .O(N__9125),
            .I(N__9030));
    ClkMux I__2144 (
            .O(N__9124),
            .I(N__9030));
    ClkMux I__2143 (
            .O(N__9123),
            .I(N__9030));
    ClkMux I__2142 (
            .O(N__9122),
            .I(N__9030));
    ClkMux I__2141 (
            .O(N__9121),
            .I(N__9030));
    ClkMux I__2140 (
            .O(N__9120),
            .I(N__9030));
    ClkMux I__2139 (
            .O(N__9119),
            .I(N__9030));
    ClkMux I__2138 (
            .O(N__9118),
            .I(N__9030));
    ClkMux I__2137 (
            .O(N__9117),
            .I(N__9030));
    ClkMux I__2136 (
            .O(N__9116),
            .I(N__9030));
    ClkMux I__2135 (
            .O(N__9115),
            .I(N__9030));
    GlobalMux I__2134 (
            .O(N__9030),
            .I(CLK80_OUT));
    InMux I__2133 (
            .O(N__9027),
            .I(N__9013));
    InMux I__2132 (
            .O(N__9026),
            .I(N__9010));
    InMux I__2131 (
            .O(N__9025),
            .I(N__9007));
    InMux I__2130 (
            .O(N__9024),
            .I(N__9000));
    InMux I__2129 (
            .O(N__9023),
            .I(N__9000));
    InMux I__2128 (
            .O(N__9022),
            .I(N__9000));
    InMux I__2127 (
            .O(N__9021),
            .I(N__8997));
    InMux I__2126 (
            .O(N__9020),
            .I(N__8994));
    InMux I__2125 (
            .O(N__9019),
            .I(N__8991));
    InMux I__2124 (
            .O(N__9018),
            .I(N__8988));
    InMux I__2123 (
            .O(N__9017),
            .I(N__8983));
    InMux I__2122 (
            .O(N__9016),
            .I(N__8983));
    LocalMux I__2121 (
            .O(N__9013),
            .I(N__8975));
    LocalMux I__2120 (
            .O(N__9010),
            .I(N__8969));
    LocalMux I__2119 (
            .O(N__9007),
            .I(N__8961));
    LocalMux I__2118 (
            .O(N__9000),
            .I(N__8958));
    LocalMux I__2117 (
            .O(N__8997),
            .I(N__8955));
    LocalMux I__2116 (
            .O(N__8994),
            .I(N__8948));
    LocalMux I__2115 (
            .O(N__8991),
            .I(N__8945));
    LocalMux I__2114 (
            .O(N__8988),
            .I(N__8939));
    LocalMux I__2113 (
            .O(N__8983),
            .I(N__8924));
    SRMux I__2112 (
            .O(N__8982),
            .I(N__8832));
    SRMux I__2111 (
            .O(N__8981),
            .I(N__8832));
    SRMux I__2110 (
            .O(N__8980),
            .I(N__8832));
    SRMux I__2109 (
            .O(N__8979),
            .I(N__8832));
    SRMux I__2108 (
            .O(N__8978),
            .I(N__8832));
    Glb2LocalMux I__2107 (
            .O(N__8975),
            .I(N__8832));
    SRMux I__2106 (
            .O(N__8974),
            .I(N__8832));
    SRMux I__2105 (
            .O(N__8973),
            .I(N__8832));
    SRMux I__2104 (
            .O(N__8972),
            .I(N__8832));
    Glb2LocalMux I__2103 (
            .O(N__8969),
            .I(N__8832));
    SRMux I__2102 (
            .O(N__8968),
            .I(N__8832));
    SRMux I__2101 (
            .O(N__8967),
            .I(N__8832));
    SRMux I__2100 (
            .O(N__8966),
            .I(N__8832));
    SRMux I__2099 (
            .O(N__8965),
            .I(N__8832));
    SRMux I__2098 (
            .O(N__8964),
            .I(N__8832));
    Glb2LocalMux I__2097 (
            .O(N__8961),
            .I(N__8832));
    Glb2LocalMux I__2096 (
            .O(N__8958),
            .I(N__8832));
    Glb2LocalMux I__2095 (
            .O(N__8955),
            .I(N__8832));
    SRMux I__2094 (
            .O(N__8954),
            .I(N__8832));
    SRMux I__2093 (
            .O(N__8953),
            .I(N__8832));
    SRMux I__2092 (
            .O(N__8952),
            .I(N__8832));
    SRMux I__2091 (
            .O(N__8951),
            .I(N__8832));
    Glb2LocalMux I__2090 (
            .O(N__8948),
            .I(N__8832));
    Glb2LocalMux I__2089 (
            .O(N__8945),
            .I(N__8832));
    SRMux I__2088 (
            .O(N__8944),
            .I(N__8832));
    SRMux I__2087 (
            .O(N__8943),
            .I(N__8832));
    SRMux I__2086 (
            .O(N__8942),
            .I(N__8832));
    Glb2LocalMux I__2085 (
            .O(N__8939),
            .I(N__8832));
    SRMux I__2084 (
            .O(N__8938),
            .I(N__8832));
    SRMux I__2083 (
            .O(N__8937),
            .I(N__8832));
    SRMux I__2082 (
            .O(N__8936),
            .I(N__8832));
    SRMux I__2081 (
            .O(N__8935),
            .I(N__8832));
    SRMux I__2080 (
            .O(N__8934),
            .I(N__8832));
    SRMux I__2079 (
            .O(N__8933),
            .I(N__8832));
    SRMux I__2078 (
            .O(N__8932),
            .I(N__8832));
    SRMux I__2077 (
            .O(N__8931),
            .I(N__8832));
    SRMux I__2076 (
            .O(N__8930),
            .I(N__8832));
    SRMux I__2075 (
            .O(N__8929),
            .I(N__8832));
    SRMux I__2074 (
            .O(N__8928),
            .I(N__8832));
    SRMux I__2073 (
            .O(N__8927),
            .I(N__8832));
    Glb2LocalMux I__2072 (
            .O(N__8924),
            .I(N__8832));
    SRMux I__2071 (
            .O(N__8923),
            .I(N__8832));
    SRMux I__2070 (
            .O(N__8922),
            .I(N__8832));
    SRMux I__2069 (
            .O(N__8921),
            .I(N__8832));
    GlobalMux I__2068 (
            .O(N__8832),
            .I(N__8829));
    gio2CtrlBuf I__2067 (
            .O(N__8829),
            .I(RESETn_c_i_g));
    InMux I__2066 (
            .O(N__8826),
            .I(N__8823));
    LocalMux I__2065 (
            .O(N__8823),
            .I(\U712_CHIP_RAM.N_372 ));
    CascadeMux I__2064 (
            .O(N__8820),
            .I(N__8814));
    InMux I__2063 (
            .O(N__8819),
            .I(N__8809));
    CascadeMux I__2062 (
            .O(N__8818),
            .I(N__8806));
    CascadeMux I__2061 (
            .O(N__8817),
            .I(N__8803));
    InMux I__2060 (
            .O(N__8814),
            .I(N__8797));
    CascadeMux I__2059 (
            .O(N__8813),
            .I(N__8794));
    InMux I__2058 (
            .O(N__8812),
            .I(N__8791));
    LocalMux I__2057 (
            .O(N__8809),
            .I(N__8785));
    InMux I__2056 (
            .O(N__8806),
            .I(N__8782));
    InMux I__2055 (
            .O(N__8803),
            .I(N__8779));
    CascadeMux I__2054 (
            .O(N__8802),
            .I(N__8776));
    CascadeMux I__2053 (
            .O(N__8801),
            .I(N__8773));
    CascadeMux I__2052 (
            .O(N__8800),
            .I(N__8770));
    LocalMux I__2051 (
            .O(N__8797),
            .I(N__8765));
    InMux I__2050 (
            .O(N__8794),
            .I(N__8762));
    LocalMux I__2049 (
            .O(N__8791),
            .I(N__8759));
    CascadeMux I__2048 (
            .O(N__8790),
            .I(N__8755));
    CascadeMux I__2047 (
            .O(N__8789),
            .I(N__8752));
    InMux I__2046 (
            .O(N__8788),
            .I(N__8749));
    Span4Mux_v I__2045 (
            .O(N__8785),
            .I(N__8744));
    LocalMux I__2044 (
            .O(N__8782),
            .I(N__8744));
    LocalMux I__2043 (
            .O(N__8779),
            .I(N__8741));
    InMux I__2042 (
            .O(N__8776),
            .I(N__8734));
    InMux I__2041 (
            .O(N__8773),
            .I(N__8734));
    InMux I__2040 (
            .O(N__8770),
            .I(N__8734));
    CascadeMux I__2039 (
            .O(N__8769),
            .I(N__8730));
    InMux I__2038 (
            .O(N__8768),
            .I(N__8727));
    Span4Mux_v I__2037 (
            .O(N__8765),
            .I(N__8724));
    LocalMux I__2036 (
            .O(N__8762),
            .I(N__8719));
    Span4Mux_h I__2035 (
            .O(N__8759),
            .I(N__8719));
    InMux I__2034 (
            .O(N__8758),
            .I(N__8714));
    InMux I__2033 (
            .O(N__8755),
            .I(N__8714));
    InMux I__2032 (
            .O(N__8752),
            .I(N__8711));
    LocalMux I__2031 (
            .O(N__8749),
            .I(N__8704));
    Span4Mux_h I__2030 (
            .O(N__8744),
            .I(N__8704));
    Span4Mux_h I__2029 (
            .O(N__8741),
            .I(N__8704));
    LocalMux I__2028 (
            .O(N__8734),
            .I(N__8701));
    InMux I__2027 (
            .O(N__8733),
            .I(N__8696));
    InMux I__2026 (
            .O(N__8730),
            .I(N__8696));
    LocalMux I__2025 (
            .O(N__8727),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2024 (
            .O(N__8724),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2023 (
            .O(N__8719),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2022 (
            .O(N__8714),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2021 (
            .O(N__8711),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2020 (
            .O(N__8704),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2019 (
            .O(N__8701),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2018 (
            .O(N__8696),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2017 (
            .O(N__8679),
            .I(N__8666));
    InMux I__2016 (
            .O(N__8678),
            .I(N__8666));
    InMux I__2015 (
            .O(N__8677),
            .I(N__8661));
    InMux I__2014 (
            .O(N__8676),
            .I(N__8661));
    CascadeMux I__2013 (
            .O(N__8675),
            .I(N__8658));
    CascadeMux I__2012 (
            .O(N__8674),
            .I(N__8655));
    InMux I__2011 (
            .O(N__8673),
            .I(N__8651));
    InMux I__2010 (
            .O(N__8672),
            .I(N__8647));
    InMux I__2009 (
            .O(N__8671),
            .I(N__8644));
    LocalMux I__2008 (
            .O(N__8666),
            .I(N__8639));
    LocalMux I__2007 (
            .O(N__8661),
            .I(N__8639));
    InMux I__2006 (
            .O(N__8658),
            .I(N__8634));
    InMux I__2005 (
            .O(N__8655),
            .I(N__8634));
    InMux I__2004 (
            .O(N__8654),
            .I(N__8631));
    LocalMux I__2003 (
            .O(N__8651),
            .I(N__8628));
    InMux I__2002 (
            .O(N__8650),
            .I(N__8625));
    LocalMux I__2001 (
            .O(N__8647),
            .I(N__8620));
    LocalMux I__2000 (
            .O(N__8644),
            .I(N__8620));
    Span4Mux_v I__1999 (
            .O(N__8639),
            .I(N__8615));
    LocalMux I__1998 (
            .O(N__8634),
            .I(N__8615));
    LocalMux I__1997 (
            .O(N__8631),
            .I(N__8610));
    Span12Mux_s9_v I__1996 (
            .O(N__8628),
            .I(N__8607));
    LocalMux I__1995 (
            .O(N__8625),
            .I(N__8600));
    Span4Mux_v I__1994 (
            .O(N__8620),
            .I(N__8600));
    Span4Mux_h I__1993 (
            .O(N__8615),
            .I(N__8600));
    InMux I__1992 (
            .O(N__8614),
            .I(N__8597));
    InMux I__1991 (
            .O(N__8613),
            .I(N__8594));
    Odrv4 I__1990 (
            .O(N__8610),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv12 I__1989 (
            .O(N__8607),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__1988 (
            .O(N__8600),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__1987 (
            .O(N__8597),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__1986 (
            .O(N__8594),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    InMux I__1985 (
            .O(N__8583),
            .I(N__8573));
    InMux I__1984 (
            .O(N__8582),
            .I(N__8568));
    InMux I__1983 (
            .O(N__8581),
            .I(N__8568));
    InMux I__1982 (
            .O(N__8580),
            .I(N__8565));
    InMux I__1981 (
            .O(N__8579),
            .I(N__8560));
    InMux I__1980 (
            .O(N__8578),
            .I(N__8560));
    InMux I__1979 (
            .O(N__8577),
            .I(N__8555));
    InMux I__1978 (
            .O(N__8576),
            .I(N__8552));
    LocalMux I__1977 (
            .O(N__8573),
            .I(N__8549));
    LocalMux I__1976 (
            .O(N__8568),
            .I(N__8546));
    LocalMux I__1975 (
            .O(N__8565),
            .I(N__8543));
    LocalMux I__1974 (
            .O(N__8560),
            .I(N__8540));
    InMux I__1973 (
            .O(N__8559),
            .I(N__8531));
    InMux I__1972 (
            .O(N__8558),
            .I(N__8531));
    LocalMux I__1971 (
            .O(N__8555),
            .I(N__8528));
    LocalMux I__1970 (
            .O(N__8552),
            .I(N__8523));
    Span4Mux_h I__1969 (
            .O(N__8549),
            .I(N__8523));
    Span4Mux_h I__1968 (
            .O(N__8546),
            .I(N__8516));
    Span4Mux_v I__1967 (
            .O(N__8543),
            .I(N__8516));
    Span4Mux_v I__1966 (
            .O(N__8540),
            .I(N__8516));
    InMux I__1965 (
            .O(N__8539),
            .I(N__8513));
    InMux I__1964 (
            .O(N__8538),
            .I(N__8508));
    InMux I__1963 (
            .O(N__8537),
            .I(N__8508));
    InMux I__1962 (
            .O(N__8536),
            .I(N__8505));
    LocalMux I__1961 (
            .O(N__8531),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1960 (
            .O(N__8528),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1959 (
            .O(N__8523),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1958 (
            .O(N__8516),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__1957 (
            .O(N__8513),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__1956 (
            .O(N__8508),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__1955 (
            .O(N__8505),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    IoInMux I__1954 (
            .O(N__8490),
            .I(N__8487));
    LocalMux I__1953 (
            .O(N__8487),
            .I(N__8484));
    Span12Mux_s1_h I__1952 (
            .O(N__8484),
            .I(N__8481));
    Span12Mux_h I__1951 (
            .O(N__8481),
            .I(N__8478));
    Odrv12 I__1950 (
            .O(N__8478),
            .I(CMA_c_5));
    CEMux I__1949 (
            .O(N__8475),
            .I(N__8471));
    CEMux I__1948 (
            .O(N__8474),
            .I(N__8468));
    LocalMux I__1947 (
            .O(N__8471),
            .I(N__8461));
    LocalMux I__1946 (
            .O(N__8468),
            .I(N__8458));
    CEMux I__1945 (
            .O(N__8467),
            .I(N__8455));
    CEMux I__1944 (
            .O(N__8466),
            .I(N__8452));
    CEMux I__1943 (
            .O(N__8465),
            .I(N__8449));
    CEMux I__1942 (
            .O(N__8464),
            .I(N__8446));
    Span4Mux_v I__1941 (
            .O(N__8461),
            .I(N__8441));
    Span4Mux_h I__1940 (
            .O(N__8458),
            .I(N__8441));
    LocalMux I__1939 (
            .O(N__8455),
            .I(N__8438));
    LocalMux I__1938 (
            .O(N__8452),
            .I(N__8431));
    LocalMux I__1937 (
            .O(N__8449),
            .I(N__8431));
    LocalMux I__1936 (
            .O(N__8446),
            .I(N__8431));
    Odrv4 I__1935 (
            .O(N__8441),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv12 I__1934 (
            .O(N__8438),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1933 (
            .O(N__8431),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    InMux I__1932 (
            .O(N__8424),
            .I(N__8420));
    InMux I__1931 (
            .O(N__8423),
            .I(N__8417));
    LocalMux I__1930 (
            .O(N__8420),
            .I(N__8414));
    LocalMux I__1929 (
            .O(N__8417),
            .I(N__8411));
    Sp12to4 I__1928 (
            .O(N__8414),
            .I(N__8408));
    Span12Mux_v I__1927 (
            .O(N__8411),
            .I(N__8405));
    Span12Mux_v I__1926 (
            .O(N__8408),
            .I(N__8402));
    Span12Mux_h I__1925 (
            .O(N__8405),
            .I(N__8399));
    Span12Mux_h I__1924 (
            .O(N__8402),
            .I(N__8396));
    Odrv12 I__1923 (
            .O(N__8399),
            .I(DRA_c_4));
    Odrv12 I__1922 (
            .O(N__8396),
            .I(DRA_c_4));
    InMux I__1921 (
            .O(N__8391),
            .I(N__8388));
    LocalMux I__1920 (
            .O(N__8388),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1919 (
            .O(N__8385),
            .I(N__8382));
    LocalMux I__1918 (
            .O(N__8382),
            .I(N__8378));
    InMux I__1917 (
            .O(N__8381),
            .I(N__8375));
    Span4Mux_h I__1916 (
            .O(N__8378),
            .I(N__8370));
    LocalMux I__1915 (
            .O(N__8375),
            .I(N__8370));
    Span4Mux_v I__1914 (
            .O(N__8370),
            .I(N__8367));
    Sp12to4 I__1913 (
            .O(N__8367),
            .I(N__8364));
    Span12Mux_h I__1912 (
            .O(N__8364),
            .I(N__8361));
    Odrv12 I__1911 (
            .O(N__8361),
            .I(DRA_c_8));
    CascadeMux I__1910 (
            .O(N__8358),
            .I(N__8355));
    InMux I__1909 (
            .O(N__8355),
            .I(N__8352));
    LocalMux I__1908 (
            .O(N__8352),
            .I(N__8349));
    Span4Mux_v I__1907 (
            .O(N__8349),
            .I(N__8346));
    Odrv4 I__1906 (
            .O(N__8346),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1905 (
            .O(N__8343),
            .I(N__8340));
    LocalMux I__1904 (
            .O(N__8340),
            .I(N__8336));
    InMux I__1903 (
            .O(N__8339),
            .I(N__8333));
    Span4Mux_v I__1902 (
            .O(N__8336),
            .I(N__8330));
    LocalMux I__1901 (
            .O(N__8333),
            .I(N__8327));
    Sp12to4 I__1900 (
            .O(N__8330),
            .I(N__8324));
    Span12Mux_v I__1899 (
            .O(N__8327),
            .I(N__8321));
    Span12Mux_h I__1898 (
            .O(N__8324),
            .I(N__8318));
    Span12Mux_h I__1897 (
            .O(N__8321),
            .I(N__8313));
    Span12Mux_v I__1896 (
            .O(N__8318),
            .I(N__8313));
    Odrv12 I__1895 (
            .O(N__8313),
            .I(DRA_c_5));
    InMux I__1894 (
            .O(N__8310),
            .I(N__8307));
    LocalMux I__1893 (
            .O(N__8307),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1892 (
            .O(N__8304),
            .I(N__8300));
    InMux I__1891 (
            .O(N__8303),
            .I(N__8297));
    LocalMux I__1890 (
            .O(N__8300),
            .I(N__8292));
    LocalMux I__1889 (
            .O(N__8297),
            .I(N__8292));
    Span4Mux_h I__1888 (
            .O(N__8292),
            .I(N__8289));
    Sp12to4 I__1887 (
            .O(N__8289),
            .I(N__8286));
    Span12Mux_v I__1886 (
            .O(N__8286),
            .I(N__8283));
    Odrv12 I__1885 (
            .O(N__8283),
            .I(DRA_c_6));
    InMux I__1884 (
            .O(N__8280),
            .I(N__8277));
    LocalMux I__1883 (
            .O(N__8277),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1882 (
            .O(N__8274),
            .I(N__8271));
    LocalMux I__1881 (
            .O(N__8271),
            .I(N__8267));
    InMux I__1880 (
            .O(N__8270),
            .I(N__8264));
    Span4Mux_h I__1879 (
            .O(N__8267),
            .I(N__8261));
    LocalMux I__1878 (
            .O(N__8264),
            .I(N__8258));
    Span4Mux_v I__1877 (
            .O(N__8261),
            .I(N__8255));
    Sp12to4 I__1876 (
            .O(N__8258),
            .I(N__8252));
    Sp12to4 I__1875 (
            .O(N__8255),
            .I(N__8247));
    Span12Mux_v I__1874 (
            .O(N__8252),
            .I(N__8247));
    Span12Mux_h I__1873 (
            .O(N__8247),
            .I(N__8244));
    Odrv12 I__1872 (
            .O(N__8244),
            .I(DRA_c_7));
    InMux I__1871 (
            .O(N__8241),
            .I(N__8238));
    LocalMux I__1870 (
            .O(N__8238),
            .I(N__8235));
    Odrv12 I__1869 (
            .O(N__8235),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1868 (
            .O(N__8232),
            .I(N__8228));
    InMux I__1867 (
            .O(N__8231),
            .I(N__8225));
    LocalMux I__1866 (
            .O(N__8228),
            .I(N__8222));
    LocalMux I__1865 (
            .O(N__8225),
            .I(N__8219));
    Span4Mux_v I__1864 (
            .O(N__8222),
            .I(N__8214));
    Span4Mux_h I__1863 (
            .O(N__8219),
            .I(N__8214));
    Sp12to4 I__1862 (
            .O(N__8214),
            .I(N__8211));
    Span12Mux_v I__1861 (
            .O(N__8211),
            .I(N__8208));
    Span12Mux_h I__1860 (
            .O(N__8208),
            .I(N__8205));
    Odrv12 I__1859 (
            .O(N__8205),
            .I(DRA_c_0));
    InMux I__1858 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1857 (
            .O(N__8199),
            .I(N__8196));
    Odrv4 I__1856 (
            .O(N__8196),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    CEMux I__1855 (
            .O(N__8193),
            .I(N__8190));
    LocalMux I__1854 (
            .O(N__8190),
            .I(N__8187));
    Span4Mux_h I__1853 (
            .O(N__8187),
            .I(N__8182));
    CEMux I__1852 (
            .O(N__8186),
            .I(N__8179));
    CEMux I__1851 (
            .O(N__8185),
            .I(N__8176));
    Odrv4 I__1850 (
            .O(N__8182),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__1849 (
            .O(N__8179),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__1848 (
            .O(N__8176),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__1847 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__1846 (
            .O(N__8166),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    CascadeMux I__1845 (
            .O(N__8163),
            .I(N__8148));
    InMux I__1844 (
            .O(N__8162),
            .I(N__8145));
    InMux I__1843 (
            .O(N__8161),
            .I(N__8139));
    InMux I__1842 (
            .O(N__8160),
            .I(N__8132));
    InMux I__1841 (
            .O(N__8159),
            .I(N__8132));
    InMux I__1840 (
            .O(N__8158),
            .I(N__8132));
    InMux I__1839 (
            .O(N__8157),
            .I(N__8125));
    InMux I__1838 (
            .O(N__8156),
            .I(N__8125));
    InMux I__1837 (
            .O(N__8155),
            .I(N__8122));
    InMux I__1836 (
            .O(N__8154),
            .I(N__8119));
    InMux I__1835 (
            .O(N__8153),
            .I(N__8112));
    InMux I__1834 (
            .O(N__8152),
            .I(N__8105));
    InMux I__1833 (
            .O(N__8151),
            .I(N__8105));
    InMux I__1832 (
            .O(N__8148),
            .I(N__8105));
    LocalMux I__1831 (
            .O(N__8145),
            .I(N__8101));
    InMux I__1830 (
            .O(N__8144),
            .I(N__8098));
    InMux I__1829 (
            .O(N__8143),
            .I(N__8095));
    InMux I__1828 (
            .O(N__8142),
            .I(N__8092));
    LocalMux I__1827 (
            .O(N__8139),
            .I(N__8087));
    LocalMux I__1826 (
            .O(N__8132),
            .I(N__8087));
    InMux I__1825 (
            .O(N__8131),
            .I(N__8082));
    InMux I__1824 (
            .O(N__8130),
            .I(N__8082));
    LocalMux I__1823 (
            .O(N__8125),
            .I(N__8077));
    LocalMux I__1822 (
            .O(N__8122),
            .I(N__8077));
    LocalMux I__1821 (
            .O(N__8119),
            .I(N__8071));
    InMux I__1820 (
            .O(N__8118),
            .I(N__8068));
    InMux I__1819 (
            .O(N__8117),
            .I(N__8065));
    InMux I__1818 (
            .O(N__8116),
            .I(N__8060));
    InMux I__1817 (
            .O(N__8115),
            .I(N__8060));
    LocalMux I__1816 (
            .O(N__8112),
            .I(N__8057));
    LocalMux I__1815 (
            .O(N__8105),
            .I(N__8054));
    InMux I__1814 (
            .O(N__8104),
            .I(N__8051));
    Span4Mux_v I__1813 (
            .O(N__8101),
            .I(N__8044));
    LocalMux I__1812 (
            .O(N__8098),
            .I(N__8044));
    LocalMux I__1811 (
            .O(N__8095),
            .I(N__8044));
    LocalMux I__1810 (
            .O(N__8092),
            .I(N__8037));
    Span4Mux_h I__1809 (
            .O(N__8087),
            .I(N__8037));
    LocalMux I__1808 (
            .O(N__8082),
            .I(N__8037));
    Span4Mux_v I__1807 (
            .O(N__8077),
            .I(N__8034));
    InMux I__1806 (
            .O(N__8076),
            .I(N__8031));
    InMux I__1805 (
            .O(N__8075),
            .I(N__8026));
    InMux I__1804 (
            .O(N__8074),
            .I(N__8026));
    Span4Mux_h I__1803 (
            .O(N__8071),
            .I(N__8023));
    LocalMux I__1802 (
            .O(N__8068),
            .I(N__8016));
    LocalMux I__1801 (
            .O(N__8065),
            .I(N__8016));
    LocalMux I__1800 (
            .O(N__8060),
            .I(N__8016));
    Span4Mux_v I__1799 (
            .O(N__8057),
            .I(N__8009));
    Span4Mux_h I__1798 (
            .O(N__8054),
            .I(N__8009));
    LocalMux I__1797 (
            .O(N__8051),
            .I(N__8009));
    Span4Mux_v I__1796 (
            .O(N__8044),
            .I(N__8004));
    Span4Mux_v I__1795 (
            .O(N__8037),
            .I(N__8004));
    Odrv4 I__1794 (
            .O(N__8034),
            .I(CPU_CYCLEm));
    LocalMux I__1793 (
            .O(N__8031),
            .I(CPU_CYCLEm));
    LocalMux I__1792 (
            .O(N__8026),
            .I(CPU_CYCLEm));
    Odrv4 I__1791 (
            .O(N__8023),
            .I(CPU_CYCLEm));
    Odrv4 I__1790 (
            .O(N__8016),
            .I(CPU_CYCLEm));
    Odrv4 I__1789 (
            .O(N__8009),
            .I(CPU_CYCLEm));
    Odrv4 I__1788 (
            .O(N__8004),
            .I(CPU_CYCLEm));
    InMux I__1787 (
            .O(N__7989),
            .I(N__7986));
    LocalMux I__1786 (
            .O(N__7986),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6 ));
    InMux I__1785 (
            .O(N__7983),
            .I(N__7980));
    LocalMux I__1784 (
            .O(N__7980),
            .I(N__7977));
    Span4Mux_h I__1783 (
            .O(N__7977),
            .I(N__7973));
    InMux I__1782 (
            .O(N__7976),
            .I(N__7970));
    Span4Mux_v I__1781 (
            .O(N__7973),
            .I(N__7967));
    LocalMux I__1780 (
            .O(N__7970),
            .I(N__7964));
    Sp12to4 I__1779 (
            .O(N__7967),
            .I(N__7959));
    Span12Mux_v I__1778 (
            .O(N__7964),
            .I(N__7959));
    Span12Mux_h I__1777 (
            .O(N__7959),
            .I(N__7956));
    Span12Mux_v I__1776 (
            .O(N__7956),
            .I(N__7953));
    Odrv12 I__1775 (
            .O(N__7953),
            .I(DRA_c_1));
    InMux I__1774 (
            .O(N__7950),
            .I(N__7947));
    LocalMux I__1773 (
            .O(N__7947),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1772 (
            .O(N__7944),
            .I(N__7941));
    LocalMux I__1771 (
            .O(N__7941),
            .I(N__7938));
    Odrv4 I__1770 (
            .O(N__7938),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    CEMux I__1769 (
            .O(N__7935),
            .I(N__7932));
    LocalMux I__1768 (
            .O(N__7932),
            .I(N__7928));
    CEMux I__1767 (
            .O(N__7931),
            .I(N__7925));
    Span4Mux_v I__1766 (
            .O(N__7928),
            .I(N__7920));
    LocalMux I__1765 (
            .O(N__7925),
            .I(N__7917));
    CEMux I__1764 (
            .O(N__7924),
            .I(N__7914));
    CEMux I__1763 (
            .O(N__7923),
            .I(N__7911));
    Span4Mux_h I__1762 (
            .O(N__7920),
            .I(N__7904));
    Span4Mux_v I__1761 (
            .O(N__7917),
            .I(N__7904));
    LocalMux I__1760 (
            .O(N__7914),
            .I(N__7904));
    LocalMux I__1759 (
            .O(N__7911),
            .I(N__7901));
    Span4Mux_h I__1758 (
            .O(N__7904),
            .I(N__7898));
    Span4Mux_h I__1757 (
            .O(N__7901),
            .I(N__7895));
    Odrv4 I__1756 (
            .O(N__7898),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__1755 (
            .O(N__7895),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    IoInMux I__1754 (
            .O(N__7890),
            .I(N__7887));
    LocalMux I__1753 (
            .O(N__7887),
            .I(N__7884));
    Span4Mux_s2_v I__1752 (
            .O(N__7884),
            .I(N__7881));
    Span4Mux_v I__1751 (
            .O(N__7881),
            .I(N__7878));
    Sp12to4 I__1750 (
            .O(N__7878),
            .I(N__7875));
    Odrv12 I__1749 (
            .O(N__7875),
            .I(CASn_c));
    IoInMux I__1748 (
            .O(N__7872),
            .I(N__7869));
    LocalMux I__1747 (
            .O(N__7869),
            .I(N__7866));
    Span12Mux_s1_h I__1746 (
            .O(N__7866),
            .I(N__7863));
    Span12Mux_h I__1745 (
            .O(N__7863),
            .I(N__7860));
    Odrv12 I__1744 (
            .O(N__7860),
            .I(WEn_c));
    InMux I__1743 (
            .O(N__7857),
            .I(N__7854));
    LocalMux I__1742 (
            .O(N__7854),
            .I(N__7850));
    InMux I__1741 (
            .O(N__7853),
            .I(N__7847));
    Span4Mux_h I__1740 (
            .O(N__7850),
            .I(N__7843));
    LocalMux I__1739 (
            .O(N__7847),
            .I(N__7840));
    InMux I__1738 (
            .O(N__7846),
            .I(N__7835));
    Span4Mux_h I__1737 (
            .O(N__7843),
            .I(N__7832));
    Span4Mux_h I__1736 (
            .O(N__7840),
            .I(N__7829));
    InMux I__1735 (
            .O(N__7839),
            .I(N__7826));
    InMux I__1734 (
            .O(N__7838),
            .I(N__7823));
    LocalMux I__1733 (
            .O(N__7835),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1732 (
            .O(N__7832),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1731 (
            .O(N__7829),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1730 (
            .O(N__7826),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1729 (
            .O(N__7823),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1728 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__1727 (
            .O(N__7809),
            .I(N__7806));
    Span4Mux_s3_v I__1726 (
            .O(N__7806),
            .I(N__7803));
    Span4Mux_h I__1725 (
            .O(N__7803),
            .I(N__7800));
    Odrv4 I__1724 (
            .O(N__7800),
            .I(CRCSn_c));
    IoInMux I__1723 (
            .O(N__7797),
            .I(N__7794));
    LocalMux I__1722 (
            .O(N__7794),
            .I(N__7791));
    Span4Mux_s3_v I__1721 (
            .O(N__7791),
            .I(N__7788));
    Span4Mux_v I__1720 (
            .O(N__7788),
            .I(N__7785));
    Span4Mux_h I__1719 (
            .O(N__7785),
            .I(N__7782));
    Odrv4 I__1718 (
            .O(N__7782),
            .I(RASn_c));
    InMux I__1717 (
            .O(N__7779),
            .I(N__7776));
    LocalMux I__1716 (
            .O(N__7776),
            .I(\U712_CHIP_RAM.N_373 ));
    IoInMux I__1715 (
            .O(N__7773),
            .I(N__7770));
    LocalMux I__1714 (
            .O(N__7770),
            .I(N__7767));
    Span4Mux_s2_h I__1713 (
            .O(N__7767),
            .I(N__7764));
    Span4Mux_v I__1712 (
            .O(N__7764),
            .I(N__7761));
    Sp12to4 I__1711 (
            .O(N__7761),
            .I(N__7758));
    Span12Mux_h I__1710 (
            .O(N__7758),
            .I(N__7755));
    Odrv12 I__1709 (
            .O(N__7755),
            .I(CMA_c_6));
    InMux I__1708 (
            .O(N__7752),
            .I(N__7749));
    LocalMux I__1707 (
            .O(N__7749),
            .I(N__7746));
    Odrv12 I__1706 (
            .O(N__7746),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1705 (
            .O(N__7743),
            .I(N__7740));
    LocalMux I__1704 (
            .O(N__7740),
            .I(N__7737));
    Span4Mux_h I__1703 (
            .O(N__7737),
            .I(N__7734));
    Odrv4 I__1702 (
            .O(N__7734),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1701 (
            .O(N__7731),
            .I(N__7728));
    LocalMux I__1700 (
            .O(N__7728),
            .I(N__7725));
    Span12Mux_v I__1699 (
            .O(N__7725),
            .I(N__7722));
    Span12Mux_h I__1698 (
            .O(N__7722),
            .I(N__7719));
    Odrv12 I__1697 (
            .O(N__7719),
            .I(A_c_14));
    InMux I__1696 (
            .O(N__7716),
            .I(N__7713));
    LocalMux I__1695 (
            .O(N__7713),
            .I(N__7710));
    Span4Mux_h I__1694 (
            .O(N__7710),
            .I(N__7707));
    Sp12to4 I__1693 (
            .O(N__7707),
            .I(N__7704));
    Span12Mux_v I__1692 (
            .O(N__7704),
            .I(N__7701));
    Span12Mux_h I__1691 (
            .O(N__7701),
            .I(N__7698));
    Odrv12 I__1690 (
            .O(N__7698),
            .I(A_c_7));
    InMux I__1689 (
            .O(N__7695),
            .I(N__7692));
    LocalMux I__1688 (
            .O(N__7692),
            .I(N__7689));
    Span4Mux_v I__1687 (
            .O(N__7689),
            .I(N__7686));
    Sp12to4 I__1686 (
            .O(N__7686),
            .I(N__7683));
    Span12Mux_h I__1685 (
            .O(N__7683),
            .I(N__7680));
    Odrv12 I__1684 (
            .O(N__7680),
            .I(A_c_13));
    CascadeMux I__1683 (
            .O(N__7677),
            .I(N__7674));
    InMux I__1682 (
            .O(N__7674),
            .I(N__7671));
    LocalMux I__1681 (
            .O(N__7671),
            .I(N__7668));
    Span4Mux_v I__1680 (
            .O(N__7668),
            .I(N__7665));
    Sp12to4 I__1679 (
            .O(N__7665),
            .I(N__7662));
    Span12Mux_h I__1678 (
            .O(N__7662),
            .I(N__7659));
    Span12Mux_v I__1677 (
            .O(N__7659),
            .I(N__7656));
    Odrv12 I__1676 (
            .O(N__7656),
            .I(A_c_6));
    InMux I__1675 (
            .O(N__7653),
            .I(N__7650));
    LocalMux I__1674 (
            .O(N__7650),
            .I(\U712_CHIP_RAM.N_371 ));
    InMux I__1673 (
            .O(N__7647),
            .I(N__7644));
    LocalMux I__1672 (
            .O(N__7644),
            .I(N__7641));
    Span4Mux_v I__1671 (
            .O(N__7641),
            .I(N__7638));
    Sp12to4 I__1670 (
            .O(N__7638),
            .I(N__7635));
    Span12Mux_h I__1669 (
            .O(N__7635),
            .I(N__7632));
    Odrv12 I__1668 (
            .O(N__7632),
            .I(A_c_15));
    CascadeMux I__1667 (
            .O(N__7629),
            .I(N__7626));
    InMux I__1666 (
            .O(N__7626),
            .I(N__7623));
    LocalMux I__1665 (
            .O(N__7623),
            .I(N__7620));
    Span12Mux_v I__1664 (
            .O(N__7620),
            .I(N__7617));
    Span12Mux_h I__1663 (
            .O(N__7617),
            .I(N__7614));
    Odrv12 I__1662 (
            .O(N__7614),
            .I(A_c_8));
    InMux I__1661 (
            .O(N__7611),
            .I(N__7608));
    LocalMux I__1660 (
            .O(N__7608),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5 ));
    InMux I__1659 (
            .O(N__7605),
            .I(N__7602));
    LocalMux I__1658 (
            .O(N__7602),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1657 (
            .O(N__7599),
            .I(N__7596));
    LocalMux I__1656 (
            .O(N__7596),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4 ));
    InMux I__1655 (
            .O(N__7593),
            .I(N__7590));
    LocalMux I__1654 (
            .O(N__7590),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1653 (
            .O(N__7587),
            .I(N__7584));
    LocalMux I__1652 (
            .O(N__7584),
            .I(N__7580));
    InMux I__1651 (
            .O(N__7583),
            .I(N__7577));
    Odrv4 I__1650 (
            .O(N__7580),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__1649 (
            .O(N__7577),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    InMux I__1648 (
            .O(N__7572),
            .I(N__7568));
    InMux I__1647 (
            .O(N__7571),
            .I(N__7565));
    LocalMux I__1646 (
            .O(N__7568),
            .I(N__7560));
    LocalMux I__1645 (
            .O(N__7565),
            .I(N__7560));
    Span4Mux_v I__1644 (
            .O(N__7560),
            .I(N__7556));
    InMux I__1643 (
            .O(N__7559),
            .I(N__7553));
    Odrv4 I__1642 (
            .O(N__7556),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__1641 (
            .O(N__7553),
            .I(\U712_REG_SM.DS_ENZ0 ));
    IoInMux I__1640 (
            .O(N__7548),
            .I(N__7545));
    LocalMux I__1639 (
            .O(N__7545),
            .I(N__7542));
    Span4Mux_s2_v I__1638 (
            .O(N__7542),
            .I(N__7539));
    Span4Mux_v I__1637 (
            .O(N__7539),
            .I(N__7536));
    Sp12to4 I__1636 (
            .O(N__7536),
            .I(N__7533));
    Span12Mux_h I__1635 (
            .O(N__7533),
            .I(N__7530));
    Odrv12 I__1634 (
            .O(N__7530),
            .I(U712_REG_SM_un1_UDSn_i));
    CascadeMux I__1633 (
            .O(N__7527),
            .I(N__7524));
    InMux I__1632 (
            .O(N__7524),
            .I(N__7513));
    InMux I__1631 (
            .O(N__7523),
            .I(N__7513));
    InMux I__1630 (
            .O(N__7522),
            .I(N__7510));
    InMux I__1629 (
            .O(N__7521),
            .I(N__7507));
    InMux I__1628 (
            .O(N__7520),
            .I(N__7504));
    InMux I__1627 (
            .O(N__7519),
            .I(N__7498));
    InMux I__1626 (
            .O(N__7518),
            .I(N__7498));
    LocalMux I__1625 (
            .O(N__7513),
            .I(N__7491));
    LocalMux I__1624 (
            .O(N__7510),
            .I(N__7491));
    LocalMux I__1623 (
            .O(N__7507),
            .I(N__7491));
    LocalMux I__1622 (
            .O(N__7504),
            .I(N__7488));
    InMux I__1621 (
            .O(N__7503),
            .I(N__7485));
    LocalMux I__1620 (
            .O(N__7498),
            .I(N__7482));
    Span4Mux_h I__1619 (
            .O(N__7491),
            .I(N__7479));
    Span4Mux_v I__1618 (
            .O(N__7488),
            .I(N__7474));
    LocalMux I__1617 (
            .O(N__7485),
            .I(N__7474));
    Span4Mux_v I__1616 (
            .O(N__7482),
            .I(N__7470));
    Span4Mux_v I__1615 (
            .O(N__7479),
            .I(N__7465));
    Span4Mux_h I__1614 (
            .O(N__7474),
            .I(N__7465));
    InMux I__1613 (
            .O(N__7473),
            .I(N__7462));
    Span4Mux_v I__1612 (
            .O(N__7470),
            .I(N__7459));
    Sp12to4 I__1611 (
            .O(N__7465),
            .I(N__7454));
    LocalMux I__1610 (
            .O(N__7462),
            .I(N__7454));
    Sp12to4 I__1609 (
            .O(N__7459),
            .I(N__7451));
    Span12Mux_v I__1608 (
            .O(N__7454),
            .I(N__7448));
    Span12Mux_h I__1607 (
            .O(N__7451),
            .I(N__7445));
    Span12Mux_h I__1606 (
            .O(N__7448),
            .I(N__7442));
    Odrv12 I__1605 (
            .O(N__7445),
            .I(RESETn_c));
    Odrv12 I__1604 (
            .O(N__7442),
            .I(RESETn_c));
    IoInMux I__1603 (
            .O(N__7437),
            .I(N__7434));
    LocalMux I__1602 (
            .O(N__7434),
            .I(N__7431));
    Span12Mux_s5_v I__1601 (
            .O(N__7431),
            .I(N__7428));
    Odrv12 I__1600 (
            .O(N__7428),
            .I(RESETn_c_i));
    InMux I__1599 (
            .O(N__7425),
            .I(N__7421));
    CascadeMux I__1598 (
            .O(N__7424),
            .I(N__7417));
    LocalMux I__1597 (
            .O(N__7421),
            .I(N__7414));
    InMux I__1596 (
            .O(N__7420),
            .I(N__7410));
    InMux I__1595 (
            .O(N__7417),
            .I(N__7407));
    Span4Mux_v I__1594 (
            .O(N__7414),
            .I(N__7404));
    InMux I__1593 (
            .O(N__7413),
            .I(N__7401));
    LocalMux I__1592 (
            .O(N__7410),
            .I(N__7398));
    LocalMux I__1591 (
            .O(N__7407),
            .I(N__7391));
    Sp12to4 I__1590 (
            .O(N__7404),
            .I(N__7391));
    LocalMux I__1589 (
            .O(N__7401),
            .I(N__7391));
    Sp12to4 I__1588 (
            .O(N__7398),
            .I(N__7388));
    Span12Mux_h I__1587 (
            .O(N__7391),
            .I(N__7385));
    Span12Mux_v I__1586 (
            .O(N__7388),
            .I(N__7382));
    Span12Mux_v I__1585 (
            .O(N__7385),
            .I(N__7377));
    Span12Mux_h I__1584 (
            .O(N__7382),
            .I(N__7377));
    Odrv12 I__1583 (
            .O(N__7377),
            .I(RnW_c));
    InMux I__1582 (
            .O(N__7374),
            .I(N__7370));
    InMux I__1581 (
            .O(N__7373),
            .I(N__7367));
    LocalMux I__1580 (
            .O(N__7370),
            .I(N__7364));
    LocalMux I__1579 (
            .O(N__7367),
            .I(N__7361));
    Span4Mux_v I__1578 (
            .O(N__7364),
            .I(N__7358));
    Span12Mux_h I__1577 (
            .O(N__7361),
            .I(N__7355));
    Sp12to4 I__1576 (
            .O(N__7358),
            .I(N__7352));
    Span12Mux_v I__1575 (
            .O(N__7355),
            .I(N__7349));
    Span12Mux_v I__1574 (
            .O(N__7352),
            .I(N__7346));
    Odrv12 I__1573 (
            .O(N__7349),
            .I(SIZ_c_0));
    Odrv12 I__1572 (
            .O(N__7346),
            .I(SIZ_c_0));
    CascadeMux I__1571 (
            .O(N__7341),
            .I(N__7337));
    CascadeMux I__1570 (
            .O(N__7340),
            .I(N__7334));
    InMux I__1569 (
            .O(N__7337),
            .I(N__7329));
    InMux I__1568 (
            .O(N__7334),
            .I(N__7329));
    LocalMux I__1567 (
            .O(N__7329),
            .I(N__7326));
    Odrv4 I__1566 (
            .O(N__7326),
            .I(\U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0 ));
    IoInMux I__1565 (
            .O(N__7323),
            .I(N__7320));
    LocalMux I__1564 (
            .O(N__7320),
            .I(N__7317));
    Span4Mux_s0_v I__1563 (
            .O(N__7317),
            .I(N__7314));
    Span4Mux_v I__1562 (
            .O(N__7314),
            .I(N__7311));
    Span4Mux_v I__1561 (
            .O(N__7311),
            .I(N__7308));
    Span4Mux_h I__1560 (
            .O(N__7308),
            .I(N__7305));
    Odrv4 I__1559 (
            .O(N__7305),
            .I(CMA_c_10));
    IoInMux I__1558 (
            .O(N__7302),
            .I(N__7299));
    LocalMux I__1557 (
            .O(N__7299),
            .I(N__7296));
    IoSpan4Mux I__1556 (
            .O(N__7296),
            .I(N__7293));
    IoSpan4Mux I__1555 (
            .O(N__7293),
            .I(N__7290));
    Span4Mux_s2_h I__1554 (
            .O(N__7290),
            .I(N__7287));
    Sp12to4 I__1553 (
            .O(N__7287),
            .I(N__7284));
    Odrv12 I__1552 (
            .O(N__7284),
            .I(CMA_c_4));
    InMux I__1551 (
            .O(N__7281),
            .I(N__7277));
    InMux I__1550 (
            .O(N__7280),
            .I(N__7274));
    LocalMux I__1549 (
            .O(N__7277),
            .I(N__7271));
    LocalMux I__1548 (
            .O(N__7274),
            .I(N__7268));
    Odrv4 I__1547 (
            .O(N__7271),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    Odrv4 I__1546 (
            .O(N__7268),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    InMux I__1545 (
            .O(N__7263),
            .I(N__7260));
    LocalMux I__1544 (
            .O(N__7260),
            .I(N__7257));
    Span4Mux_v I__1543 (
            .O(N__7257),
            .I(N__7254));
    Sp12to4 I__1542 (
            .O(N__7254),
            .I(N__7251));
    Span12Mux_h I__1541 (
            .O(N__7251),
            .I(N__7248));
    Odrv12 I__1540 (
            .O(N__7248),
            .I(A_c_17));
    IoInMux I__1539 (
            .O(N__7245),
            .I(N__7242));
    LocalMux I__1538 (
            .O(N__7242),
            .I(N__7239));
    Span4Mux_s2_h I__1537 (
            .O(N__7239),
            .I(N__7236));
    Span4Mux_v I__1536 (
            .O(N__7236),
            .I(N__7233));
    Span4Mux_h I__1535 (
            .O(N__7233),
            .I(N__7230));
    Sp12to4 I__1534 (
            .O(N__7230),
            .I(N__7227));
    Odrv12 I__1533 (
            .O(N__7227),
            .I(CMA_c_8));
    InMux I__1532 (
            .O(N__7224),
            .I(N__7221));
    LocalMux I__1531 (
            .O(N__7221),
            .I(N__7218));
    Span4Mux_v I__1530 (
            .O(N__7218),
            .I(N__7215));
    Span4Mux_v I__1529 (
            .O(N__7215),
            .I(N__7212));
    Sp12to4 I__1528 (
            .O(N__7212),
            .I(N__7209));
    Span12Mux_h I__1527 (
            .O(N__7209),
            .I(N__7206));
    Odrv12 I__1526 (
            .O(N__7206),
            .I(A_c_9));
    CascadeMux I__1525 (
            .O(N__7203),
            .I(N__7200));
    InMux I__1524 (
            .O(N__7200),
            .I(N__7197));
    LocalMux I__1523 (
            .O(N__7197),
            .I(N__7194));
    Span4Mux_h I__1522 (
            .O(N__7194),
            .I(N__7191));
    Span4Mux_v I__1521 (
            .O(N__7191),
            .I(N__7188));
    Sp12to4 I__1520 (
            .O(N__7188),
            .I(N__7185));
    Span12Mux_h I__1519 (
            .O(N__7185),
            .I(N__7182));
    Span12Mux_v I__1518 (
            .O(N__7182),
            .I(N__7179));
    Odrv12 I__1517 (
            .O(N__7179),
            .I(A_c_2));
    CascadeMux I__1516 (
            .O(N__7176),
            .I(\U712_CHIP_RAM.N_367_cascade_ ));
    IoInMux I__1515 (
            .O(N__7173),
            .I(N__7170));
    LocalMux I__1514 (
            .O(N__7170),
            .I(N__7167));
    Span4Mux_s3_v I__1513 (
            .O(N__7167),
            .I(N__7164));
    Span4Mux_v I__1512 (
            .O(N__7164),
            .I(N__7161));
    Span4Mux_h I__1511 (
            .O(N__7161),
            .I(N__7158));
    Odrv4 I__1510 (
            .O(N__7158),
            .I(CMA_c_0));
    InMux I__1509 (
            .O(N__7155),
            .I(N__7152));
    LocalMux I__1508 (
            .O(N__7152),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0 ));
    InMux I__1507 (
            .O(N__7149),
            .I(N__7143));
    InMux I__1506 (
            .O(N__7148),
            .I(N__7138));
    InMux I__1505 (
            .O(N__7147),
            .I(N__7133));
    InMux I__1504 (
            .O(N__7146),
            .I(N__7133));
    LocalMux I__1503 (
            .O(N__7143),
            .I(N__7130));
    InMux I__1502 (
            .O(N__7142),
            .I(N__7125));
    InMux I__1501 (
            .O(N__7141),
            .I(N__7125));
    LocalMux I__1500 (
            .O(N__7138),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1499 (
            .O(N__7133),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1498 (
            .O(N__7130),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1497 (
            .O(N__7125),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1496 (
            .O(N__7116),
            .I(N__7109));
    InMux I__1495 (
            .O(N__7115),
            .I(N__7109));
    InMux I__1494 (
            .O(N__7114),
            .I(N__7106));
    LocalMux I__1493 (
            .O(N__7109),
            .I(N__7101));
    LocalMux I__1492 (
            .O(N__7106),
            .I(N__7101));
    Span4Mux_h I__1491 (
            .O(N__7101),
            .I(N__7096));
    InMux I__1490 (
            .O(N__7100),
            .I(N__7093));
    InMux I__1489 (
            .O(N__7099),
            .I(N__7090));
    Odrv4 I__1488 (
            .O(N__7096),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__1487 (
            .O(N__7093),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__1486 (
            .O(N__7090),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__1485 (
            .O(N__7083),
            .I(N__7080));
    LocalMux I__1484 (
            .O(N__7080),
            .I(N__7077));
    Span4Mux_v I__1483 (
            .O(N__7077),
            .I(N__7074));
    Odrv4 I__1482 (
            .O(N__7074),
            .I(\U712_BYTE_ENABLE.N_453 ));
    CascadeMux I__1481 (
            .O(N__7071),
            .I(N__7068));
    InMux I__1480 (
            .O(N__7068),
            .I(N__7065));
    LocalMux I__1479 (
            .O(N__7065),
            .I(N__7062));
    Span4Mux_h I__1478 (
            .O(N__7062),
            .I(N__7059));
    Span4Mux_h I__1477 (
            .O(N__7059),
            .I(N__7055));
    InMux I__1476 (
            .O(N__7058),
            .I(N__7052));
    Odrv4 I__1475 (
            .O(N__7055),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0 ));
    LocalMux I__1474 (
            .O(N__7052),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0 ));
    InMux I__1473 (
            .O(N__7047),
            .I(N__7043));
    InMux I__1472 (
            .O(N__7046),
            .I(N__7040));
    LocalMux I__1471 (
            .O(N__7043),
            .I(N__7036));
    LocalMux I__1470 (
            .O(N__7040),
            .I(N__7033));
    InMux I__1469 (
            .O(N__7039),
            .I(N__7030));
    Odrv12 I__1468 (
            .O(N__7036),
            .I(\U712_BYTE_ENABLE.N_451 ));
    Odrv4 I__1467 (
            .O(N__7033),
            .I(\U712_BYTE_ENABLE.N_451 ));
    LocalMux I__1466 (
            .O(N__7030),
            .I(\U712_BYTE_ENABLE.N_451 ));
    IoInMux I__1465 (
            .O(N__7023),
            .I(N__7020));
    LocalMux I__1464 (
            .O(N__7020),
            .I(N__7017));
    IoSpan4Mux I__1463 (
            .O(N__7017),
            .I(N__7014));
    IoSpan4Mux I__1462 (
            .O(N__7014),
            .I(N__7011));
    Span4Mux_s3_h I__1461 (
            .O(N__7011),
            .I(N__7008));
    Sp12to4 I__1460 (
            .O(N__7008),
            .I(N__7005));
    Odrv12 I__1459 (
            .O(N__7005),
            .I(N_50_i));
    InMux I__1458 (
            .O(N__7002),
            .I(N__6998));
    InMux I__1457 (
            .O(N__7001),
            .I(N__6995));
    LocalMux I__1456 (
            .O(N__6998),
            .I(N__6992));
    LocalMux I__1455 (
            .O(N__6995),
            .I(N__6989));
    Odrv4 I__1454 (
            .O(N__6992),
            .I(\U712_REG_SM.N_354 ));
    Odrv4 I__1453 (
            .O(N__6989),
            .I(\U712_REG_SM.N_354 ));
    InMux I__1452 (
            .O(N__6984),
            .I(N__6980));
    InMux I__1451 (
            .O(N__6983),
            .I(N__6977));
    LocalMux I__1450 (
            .O(N__6980),
            .I(\U712_REG_SM.N_394 ));
    LocalMux I__1449 (
            .O(N__6977),
            .I(\U712_REG_SM.N_394 ));
    InMux I__1448 (
            .O(N__6972),
            .I(N__6969));
    LocalMux I__1447 (
            .O(N__6969),
            .I(\U712_REG_SM.N_364 ));
    InMux I__1446 (
            .O(N__6966),
            .I(N__6962));
    InMux I__1445 (
            .O(N__6965),
            .I(N__6959));
    LocalMux I__1444 (
            .O(N__6962),
            .I(N__6956));
    LocalMux I__1443 (
            .O(N__6959),
            .I(N__6953));
    Span4Mux_h I__1442 (
            .O(N__6956),
            .I(N__6948));
    Span4Mux_h I__1441 (
            .O(N__6953),
            .I(N__6945));
    InMux I__1440 (
            .O(N__6952),
            .I(N__6942));
    InMux I__1439 (
            .O(N__6951),
            .I(N__6939));
    Odrv4 I__1438 (
            .O(N__6948),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__1437 (
            .O(N__6945),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__1436 (
            .O(N__6942),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__1435 (
            .O(N__6939),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__1434 (
            .O(N__6930),
            .I(N__6927));
    InMux I__1433 (
            .O(N__6927),
            .I(N__6922));
    InMux I__1432 (
            .O(N__6926),
            .I(N__6919));
    InMux I__1431 (
            .O(N__6925),
            .I(N__6916));
    LocalMux I__1430 (
            .O(N__6922),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__1429 (
            .O(N__6919),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__1428 (
            .O(N__6916),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__1427 (
            .O(N__6909),
            .I(N__6904));
    InMux I__1426 (
            .O(N__6908),
            .I(N__6899));
    InMux I__1425 (
            .O(N__6907),
            .I(N__6899));
    LocalMux I__1424 (
            .O(N__6904),
            .I(N__6894));
    LocalMux I__1423 (
            .O(N__6899),
            .I(N__6894));
    Span4Mux_v I__1422 (
            .O(N__6894),
            .I(N__6889));
    InMux I__1421 (
            .O(N__6893),
            .I(N__6884));
    InMux I__1420 (
            .O(N__6892),
            .I(N__6884));
    Span4Mux_h I__1419 (
            .O(N__6889),
            .I(N__6879));
    LocalMux I__1418 (
            .O(N__6884),
            .I(N__6879));
    Sp12to4 I__1417 (
            .O(N__6879),
            .I(N__6876));
    Span12Mux_v I__1416 (
            .O(N__6876),
            .I(N__6873));
    Odrv12 I__1415 (
            .O(N__6873),
            .I(A_c_0));
    CascadeMux I__1414 (
            .O(N__6870),
            .I(N__6867));
    InMux I__1413 (
            .O(N__6867),
            .I(N__6864));
    LocalMux I__1412 (
            .O(N__6864),
            .I(N__6857));
    InMux I__1411 (
            .O(N__6863),
            .I(N__6852));
    InMux I__1410 (
            .O(N__6862),
            .I(N__6852));
    InMux I__1409 (
            .O(N__6861),
            .I(N__6849));
    InMux I__1408 (
            .O(N__6860),
            .I(N__6846));
    Odrv4 I__1407 (
            .O(N__6857),
            .I(\U712_REG_SM.N_395 ));
    LocalMux I__1406 (
            .O(N__6852),
            .I(\U712_REG_SM.N_395 ));
    LocalMux I__1405 (
            .O(N__6849),
            .I(\U712_REG_SM.N_395 ));
    LocalMux I__1404 (
            .O(N__6846),
            .I(\U712_REG_SM.N_395 ));
    InMux I__1403 (
            .O(N__6837),
            .I(N__6833));
    InMux I__1402 (
            .O(N__6836),
            .I(N__6830));
    LocalMux I__1401 (
            .O(N__6833),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__1400 (
            .O(N__6830),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__1399 (
            .O(N__6825),
            .I(N__6822));
    LocalMux I__1398 (
            .O(N__6822),
            .I(N__6819));
    Span12Mux_s5_v I__1397 (
            .O(N__6819),
            .I(N__6816));
    Span12Mux_h I__1396 (
            .O(N__6816),
            .I(N__6813));
    Odrv12 I__1395 (
            .O(N__6813),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__1394 (
            .O(N__6810),
            .I(N__6804));
    InMux I__1393 (
            .O(N__6809),
            .I(N__6801));
    InMux I__1392 (
            .O(N__6808),
            .I(N__6798));
    InMux I__1391 (
            .O(N__6807),
            .I(N__6795));
    LocalMux I__1390 (
            .O(N__6804),
            .I(N__6792));
    LocalMux I__1389 (
            .O(N__6801),
            .I(N__6787));
    LocalMux I__1388 (
            .O(N__6798),
            .I(N__6787));
    LocalMux I__1387 (
            .O(N__6795),
            .I(\U712_REG_SM.N_348 ));
    Odrv4 I__1386 (
            .O(N__6792),
            .I(\U712_REG_SM.N_348 ));
    Odrv4 I__1385 (
            .O(N__6787),
            .I(\U712_REG_SM.N_348 ));
    InMux I__1384 (
            .O(N__6780),
            .I(N__6775));
    InMux I__1383 (
            .O(N__6779),
            .I(N__6772));
    InMux I__1382 (
            .O(N__6778),
            .I(N__6769));
    LocalMux I__1381 (
            .O(N__6775),
            .I(N__6759));
    LocalMux I__1380 (
            .O(N__6772),
            .I(N__6759));
    LocalMux I__1379 (
            .O(N__6769),
            .I(N__6759));
    InMux I__1378 (
            .O(N__6768),
            .I(N__6756));
    InMux I__1377 (
            .O(N__6767),
            .I(N__6751));
    InMux I__1376 (
            .O(N__6766),
            .I(N__6751));
    Odrv4 I__1375 (
            .O(N__6759),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1374 (
            .O(N__6756),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1373 (
            .O(N__6751),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__1372 (
            .O(N__6744),
            .I(N__6740));
    CascadeMux I__1371 (
            .O(N__6743),
            .I(N__6737));
    InMux I__1370 (
            .O(N__6740),
            .I(N__6734));
    InMux I__1369 (
            .O(N__6737),
            .I(N__6729));
    LocalMux I__1368 (
            .O(N__6734),
            .I(N__6726));
    InMux I__1367 (
            .O(N__6733),
            .I(N__6723));
    InMux I__1366 (
            .O(N__6732),
            .I(N__6717));
    LocalMux I__1365 (
            .O(N__6729),
            .I(N__6710));
    Span4Mux_h I__1364 (
            .O(N__6726),
            .I(N__6710));
    LocalMux I__1363 (
            .O(N__6723),
            .I(N__6710));
    InMux I__1362 (
            .O(N__6722),
            .I(N__6705));
    InMux I__1361 (
            .O(N__6721),
            .I(N__6705));
    InMux I__1360 (
            .O(N__6720),
            .I(N__6702));
    LocalMux I__1359 (
            .O(N__6717),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__1358 (
            .O(N__6710),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1357 (
            .O(N__6705),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1356 (
            .O(N__6702),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__1355 (
            .O(N__6693),
            .I(N__6688));
    InMux I__1354 (
            .O(N__6692),
            .I(N__6685));
    InMux I__1353 (
            .O(N__6691),
            .I(N__6682));
    LocalMux I__1352 (
            .O(N__6688),
            .I(N__6677));
    LocalMux I__1351 (
            .O(N__6685),
            .I(N__6677));
    LocalMux I__1350 (
            .O(N__6682),
            .I(\U712_REG_SM.N_347 ));
    Odrv4 I__1349 (
            .O(N__6677),
            .I(\U712_REG_SM.N_347 ));
    InMux I__1348 (
            .O(N__6672),
            .I(N__6669));
    LocalMux I__1347 (
            .O(N__6669),
            .I(\U712_REG_SM.N_433 ));
    InMux I__1346 (
            .O(N__6666),
            .I(N__6663));
    LocalMux I__1345 (
            .O(N__6663),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i ));
    InMux I__1344 (
            .O(N__6660),
            .I(N__6657));
    LocalMux I__1343 (
            .O(N__6657),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1342 (
            .O(N__6654),
            .I(N__6651));
    LocalMux I__1341 (
            .O(N__6651),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1340 (
            .O(N__6648),
            .I(N__6645));
    LocalMux I__1339 (
            .O(N__6645),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    CascadeMux I__1338 (
            .O(N__6642),
            .I(N__6639));
    InMux I__1337 (
            .O(N__6639),
            .I(N__6636));
    LocalMux I__1336 (
            .O(N__6636),
            .I(N__6633));
    Span12Mux_v I__1335 (
            .O(N__6633),
            .I(N__6630));
    Span12Mux_h I__1334 (
            .O(N__6630),
            .I(N__6627));
    Odrv12 I__1333 (
            .O(N__6627),
            .I(A_c_19));
    IoInMux I__1332 (
            .O(N__6624),
            .I(N__6621));
    LocalMux I__1331 (
            .O(N__6621),
            .I(N__6618));
    Span4Mux_s3_h I__1330 (
            .O(N__6618),
            .I(N__6615));
    Span4Mux_v I__1329 (
            .O(N__6615),
            .I(N__6612));
    Sp12to4 I__1328 (
            .O(N__6612),
            .I(N__6609));
    Span12Mux_h I__1327 (
            .O(N__6609),
            .I(N__6606));
    Odrv12 I__1326 (
            .O(N__6606),
            .I(CMA_c_9));
    InMux I__1325 (
            .O(N__6603),
            .I(N__6600));
    LocalMux I__1324 (
            .O(N__6600),
            .I(N__6597));
    Odrv4 I__1323 (
            .O(N__6597),
            .I(\U712_CHIP_RAM.N_374 ));
    IoInMux I__1322 (
            .O(N__6594),
            .I(N__6591));
    LocalMux I__1321 (
            .O(N__6591),
            .I(N__6588));
    IoSpan4Mux I__1320 (
            .O(N__6588),
            .I(N__6585));
    IoSpan4Mux I__1319 (
            .O(N__6585),
            .I(N__6582));
    Sp12to4 I__1318 (
            .O(N__6582),
            .I(N__6579));
    Span12Mux_s7_h I__1317 (
            .O(N__6579),
            .I(N__6576));
    Odrv12 I__1316 (
            .O(N__6576),
            .I(CMA_c_7));
    InMux I__1315 (
            .O(N__6573),
            .I(N__6570));
    LocalMux I__1314 (
            .O(N__6570),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1313 (
            .O(N__6567),
            .I(N__6563));
    InMux I__1312 (
            .O(N__6566),
            .I(N__6560));
    LocalMux I__1311 (
            .O(N__6563),
            .I(N__6555));
    LocalMux I__1310 (
            .O(N__6560),
            .I(N__6555));
    Span4Mux_v I__1309 (
            .O(N__6555),
            .I(N__6552));
    Sp12to4 I__1308 (
            .O(N__6552),
            .I(N__6549));
    Span12Mux_h I__1307 (
            .O(N__6549),
            .I(N__6546));
    Span12Mux_v I__1306 (
            .O(N__6546),
            .I(N__6543));
    Odrv12 I__1305 (
            .O(N__6543),
            .I(DRA_c_3));
    InMux I__1304 (
            .O(N__6540),
            .I(N__6537));
    LocalMux I__1303 (
            .O(N__6537),
            .I(N__6534));
    Odrv12 I__1302 (
            .O(N__6534),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1301 (
            .O(N__6531),
            .I(N__6528));
    LocalMux I__1300 (
            .O(N__6528),
            .I(N__6524));
    InMux I__1299 (
            .O(N__6527),
            .I(N__6521));
    Span4Mux_v I__1298 (
            .O(N__6524),
            .I(N__6518));
    LocalMux I__1297 (
            .O(N__6521),
            .I(N__6515));
    Sp12to4 I__1296 (
            .O(N__6518),
            .I(N__6512));
    Span12Mux_h I__1295 (
            .O(N__6515),
            .I(N__6509));
    Span12Mux_h I__1294 (
            .O(N__6512),
            .I(N__6506));
    Span12Mux_v I__1293 (
            .O(N__6509),
            .I(N__6503));
    Span12Mux_v I__1292 (
            .O(N__6506),
            .I(N__6500));
    Odrv12 I__1291 (
            .O(N__6503),
            .I(DRA_c_2));
    Odrv12 I__1290 (
            .O(N__6500),
            .I(DRA_c_2));
    CascadeMux I__1289 (
            .O(N__6495),
            .I(N__6492));
    InMux I__1288 (
            .O(N__6492),
            .I(N__6489));
    LocalMux I__1287 (
            .O(N__6489),
            .I(N__6486));
    Odrv12 I__1286 (
            .O(N__6486),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1285 (
            .O(N__6483),
            .I(N__6480));
    LocalMux I__1284 (
            .O(N__6480),
            .I(N__6477));
    Span4Mux_h I__1283 (
            .O(N__6477),
            .I(N__6472));
    InMux I__1282 (
            .O(N__6476),
            .I(N__6467));
    InMux I__1281 (
            .O(N__6475),
            .I(N__6467));
    Odrv4 I__1280 (
            .O(N__6472),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1279 (
            .O(N__6467),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1278 (
            .O(N__6462),
            .I(\U712_REG_SM.N_364_cascade_ ));
    InMux I__1277 (
            .O(N__6459),
            .I(N__6455));
    CascadeMux I__1276 (
            .O(N__6458),
            .I(N__6451));
    LocalMux I__1275 (
            .O(N__6455),
            .I(N__6448));
    InMux I__1274 (
            .O(N__6454),
            .I(N__6443));
    InMux I__1273 (
            .O(N__6451),
            .I(N__6443));
    Span4Mux_h I__1272 (
            .O(N__6448),
            .I(N__6440));
    LocalMux I__1271 (
            .O(N__6443),
            .I(\U712_REG_SM.N_343 ));
    Odrv4 I__1270 (
            .O(N__6440),
            .I(\U712_REG_SM.N_343 ));
    InMux I__1269 (
            .O(N__6435),
            .I(N__6432));
    LocalMux I__1268 (
            .O(N__6432),
            .I(N__6429));
    Span4Mux_h I__1267 (
            .O(N__6429),
            .I(N__6425));
    InMux I__1266 (
            .O(N__6428),
            .I(N__6422));
    Odrv4 I__1265 (
            .O(N__6425),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__1264 (
            .O(N__6422),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    InMux I__1263 (
            .O(N__6417),
            .I(N__6414));
    LocalMux I__1262 (
            .O(N__6414),
            .I(N__6411));
    Span12Mux_h I__1261 (
            .O(N__6411),
            .I(N__6408));
    Span12Mux_v I__1260 (
            .O(N__6408),
            .I(N__6405));
    Odrv12 I__1259 (
            .O(N__6405),
            .I(C3_c));
    CascadeMux I__1258 (
            .O(N__6402),
            .I(N__6399));
    InMux I__1257 (
            .O(N__6399),
            .I(N__6395));
    InMux I__1256 (
            .O(N__6398),
            .I(N__6392));
    LocalMux I__1255 (
            .O(N__6395),
            .I(N__6388));
    LocalMux I__1254 (
            .O(N__6392),
            .I(N__6384));
    InMux I__1253 (
            .O(N__6391),
            .I(N__6381));
    Span4Mux_v I__1252 (
            .O(N__6388),
            .I(N__6378));
    InMux I__1251 (
            .O(N__6387),
            .I(N__6375));
    Odrv12 I__1250 (
            .O(N__6384),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1249 (
            .O(N__6381),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__1248 (
            .O(N__6378),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1247 (
            .O(N__6375),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1246 (
            .O(N__6366),
            .I(N__6363));
    LocalMux I__1245 (
            .O(N__6363),
            .I(\U712_CHIP_RAM.N_370 ));
    IoInMux I__1244 (
            .O(N__6360),
            .I(N__6357));
    LocalMux I__1243 (
            .O(N__6357),
            .I(N__6354));
    Span4Mux_s3_h I__1242 (
            .O(N__6354),
            .I(N__6351));
    Span4Mux_v I__1241 (
            .O(N__6351),
            .I(N__6348));
    Span4Mux_h I__1240 (
            .O(N__6348),
            .I(N__6345));
    Span4Mux_h I__1239 (
            .O(N__6345),
            .I(N__6342));
    Span4Mux_h I__1238 (
            .O(N__6342),
            .I(N__6339));
    Odrv4 I__1237 (
            .O(N__6339),
            .I(CMA_c_3));
    IoInMux I__1236 (
            .O(N__6336),
            .I(N__6333));
    LocalMux I__1235 (
            .O(N__6333),
            .I(N__6330));
    Odrv12 I__1234 (
            .O(N__6330),
            .I(CMA_c_1));
    InMux I__1233 (
            .O(N__6327),
            .I(N__6324));
    LocalMux I__1232 (
            .O(N__6324),
            .I(N__6321));
    Span4Mux_v I__1231 (
            .O(N__6321),
            .I(N__6318));
    Sp12to4 I__1230 (
            .O(N__6318),
            .I(N__6315));
    Span12Mux_h I__1229 (
            .O(N__6315),
            .I(N__6312));
    Span12Mux_v I__1228 (
            .O(N__6312),
            .I(N__6309));
    Odrv12 I__1227 (
            .O(N__6309),
            .I(A_c_3));
    InMux I__1226 (
            .O(N__6306),
            .I(N__6303));
    LocalMux I__1225 (
            .O(N__6303),
            .I(N__6300));
    Span4Mux_v I__1224 (
            .O(N__6300),
            .I(N__6297));
    Sp12to4 I__1223 (
            .O(N__6297),
            .I(N__6294));
    Span12Mux_h I__1222 (
            .O(N__6294),
            .I(N__6291));
    Odrv12 I__1221 (
            .O(N__6291),
            .I(A_c_10));
    CascadeMux I__1220 (
            .O(N__6288),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_ ));
    InMux I__1219 (
            .O(N__6285),
            .I(N__6282));
    LocalMux I__1218 (
            .O(N__6282),
            .I(\U712_CHIP_RAM.N_368 ));
    InMux I__1217 (
            .O(N__6279),
            .I(N__6276));
    LocalMux I__1216 (
            .O(N__6276),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2 ));
    CascadeMux I__1215 (
            .O(N__6273),
            .I(\U712_REG_SM.N_347_cascade_ ));
    InMux I__1214 (
            .O(N__6270),
            .I(N__6267));
    LocalMux I__1213 (
            .O(N__6267),
            .I(\U712_REG_SM.N_559 ));
    CascadeMux I__1212 (
            .O(N__6264),
            .I(\U712_REG_SM.N_559_cascade_ ));
    InMux I__1211 (
            .O(N__6261),
            .I(N__6255));
    InMux I__1210 (
            .O(N__6260),
            .I(N__6252));
    InMux I__1209 (
            .O(N__6259),
            .I(N__6247));
    InMux I__1208 (
            .O(N__6258),
            .I(N__6247));
    LocalMux I__1207 (
            .O(N__6255),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1206 (
            .O(N__6252),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1205 (
            .O(N__6247),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__1204 (
            .O(N__6240),
            .I(N__6237));
    InMux I__1203 (
            .O(N__6237),
            .I(N__6228));
    InMux I__1202 (
            .O(N__6236),
            .I(N__6228));
    InMux I__1201 (
            .O(N__6235),
            .I(N__6228));
    LocalMux I__1200 (
            .O(N__6228),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__1199 (
            .O(N__6225),
            .I(N__6221));
    InMux I__1198 (
            .O(N__6224),
            .I(N__6218));
    LocalMux I__1197 (
            .O(N__6221),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    LocalMux I__1196 (
            .O(N__6218),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    IoInMux I__1195 (
            .O(N__6213),
            .I(N__6209));
    IoInMux I__1194 (
            .O(N__6212),
            .I(N__6206));
    LocalMux I__1193 (
            .O(N__6209),
            .I(N__6203));
    LocalMux I__1192 (
            .O(N__6206),
            .I(N__6200));
    IoSpan4Mux I__1191 (
            .O(N__6203),
            .I(N__6197));
    IoSpan4Mux I__1190 (
            .O(N__6200),
            .I(N__6194));
    Span4Mux_s2_v I__1189 (
            .O(N__6197),
            .I(N__6191));
    Span4Mux_s2_v I__1188 (
            .O(N__6194),
            .I(N__6188));
    Sp12to4 I__1187 (
            .O(N__6191),
            .I(N__6185));
    Sp12to4 I__1186 (
            .O(N__6188),
            .I(N__6182));
    Span12Mux_s8_v I__1185 (
            .O(N__6185),
            .I(N__6179));
    Span12Mux_s8_v I__1184 (
            .O(N__6182),
            .I(N__6176));
    Span12Mux_h I__1183 (
            .O(N__6179),
            .I(N__6171));
    Span12Mux_h I__1182 (
            .O(N__6176),
            .I(N__6171));
    Odrv12 I__1181 (
            .O(N__6171),
            .I(ASn_c));
    InMux I__1180 (
            .O(N__6168),
            .I(N__6165));
    LocalMux I__1179 (
            .O(N__6165),
            .I(N__6161));
    InMux I__1178 (
            .O(N__6164),
            .I(N__6158));
    Odrv4 I__1177 (
            .O(N__6161),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1176 (
            .O(N__6158),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1175 (
            .O(N__6153),
            .I(N__6150));
    LocalMux I__1174 (
            .O(N__6150),
            .I(N__6145));
    InMux I__1173 (
            .O(N__6149),
            .I(N__6142));
    InMux I__1172 (
            .O(N__6148),
            .I(N__6139));
    Odrv4 I__1171 (
            .O(N__6145),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1170 (
            .O(N__6142),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1169 (
            .O(N__6139),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1168 (
            .O(N__6132),
            .I(N__6128));
    InMux I__1167 (
            .O(N__6131),
            .I(N__6125));
    LocalMux I__1166 (
            .O(N__6128),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ));
    LocalMux I__1165 (
            .O(N__6125),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ));
    CEMux I__1164 (
            .O(N__6120),
            .I(N__6117));
    LocalMux I__1163 (
            .O(N__6117),
            .I(\U712_REG_SM.N_186_0 ));
    CascadeMux I__1162 (
            .O(N__6114),
            .I(\U712_REG_SM.N_348_cascade_ ));
    InMux I__1161 (
            .O(N__6111),
            .I(N__6103));
    InMux I__1160 (
            .O(N__6110),
            .I(N__6103));
    InMux I__1159 (
            .O(N__6109),
            .I(N__6098));
    InMux I__1158 (
            .O(N__6108),
            .I(N__6098));
    LocalMux I__1157 (
            .O(N__6103),
            .I(N__6094));
    LocalMux I__1156 (
            .O(N__6098),
            .I(N__6091));
    CascadeMux I__1155 (
            .O(N__6097),
            .I(N__6087));
    Span4Mux_v I__1154 (
            .O(N__6094),
            .I(N__6079));
    Span4Mux_v I__1153 (
            .O(N__6091),
            .I(N__6079));
    InMux I__1152 (
            .O(N__6090),
            .I(N__6074));
    InMux I__1151 (
            .O(N__6087),
            .I(N__6074));
    InMux I__1150 (
            .O(N__6086),
            .I(N__6071));
    InMux I__1149 (
            .O(N__6085),
            .I(N__6068));
    InMux I__1148 (
            .O(N__6084),
            .I(N__6065));
    Odrv4 I__1147 (
            .O(N__6079),
            .I(DMA_CYCLEm));
    LocalMux I__1146 (
            .O(N__6074),
            .I(DMA_CYCLEm));
    LocalMux I__1145 (
            .O(N__6071),
            .I(DMA_CYCLEm));
    LocalMux I__1144 (
            .O(N__6068),
            .I(DMA_CYCLEm));
    LocalMux I__1143 (
            .O(N__6065),
            .I(DMA_CYCLEm));
    CascadeMux I__1142 (
            .O(N__6054),
            .I(N__6047));
    InMux I__1141 (
            .O(N__6053),
            .I(N__6042));
    InMux I__1140 (
            .O(N__6052),
            .I(N__6042));
    CascadeMux I__1139 (
            .O(N__6051),
            .I(N__6039));
    CascadeMux I__1138 (
            .O(N__6050),
            .I(N__6034));
    InMux I__1137 (
            .O(N__6047),
            .I(N__6031));
    LocalMux I__1136 (
            .O(N__6042),
            .I(N__6028));
    InMux I__1135 (
            .O(N__6039),
            .I(N__6023));
    InMux I__1134 (
            .O(N__6038),
            .I(N__6023));
    InMux I__1133 (
            .O(N__6037),
            .I(N__6018));
    InMux I__1132 (
            .O(N__6034),
            .I(N__6018));
    LocalMux I__1131 (
            .O(N__6031),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1130 (
            .O(N__6028),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1129 (
            .O(N__6023),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1128 (
            .O(N__6018),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1127 (
            .O(N__6009),
            .I(N__6005));
    InMux I__1126 (
            .O(N__6008),
            .I(N__6002));
    LocalMux I__1125 (
            .O(N__6005),
            .I(\U712_REG_SM.N_361 ));
    LocalMux I__1124 (
            .O(N__6002),
            .I(\U712_REG_SM.N_361 ));
    CascadeMux I__1123 (
            .O(N__5997),
            .I(N__5994));
    InMux I__1122 (
            .O(N__5994),
            .I(N__5990));
    InMux I__1121 (
            .O(N__5993),
            .I(N__5986));
    LocalMux I__1120 (
            .O(N__5990),
            .I(N__5983));
    InMux I__1119 (
            .O(N__5989),
            .I(N__5980));
    LocalMux I__1118 (
            .O(N__5986),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    Odrv4 I__1117 (
            .O(N__5983),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1116 (
            .O(N__5980),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__1115 (
            .O(N__5973),
            .I(N__5970));
    LocalMux I__1114 (
            .O(N__5970),
            .I(N__5967));
    Span4Mux_v I__1113 (
            .O(N__5967),
            .I(N__5964));
    Sp12to4 I__1112 (
            .O(N__5964),
            .I(N__5961));
    Span12Mux_h I__1111 (
            .O(N__5961),
            .I(N__5958));
    Span12Mux_v I__1110 (
            .O(N__5958),
            .I(N__5955));
    Odrv12 I__1109 (
            .O(N__5955),
            .I(DBRn_c));
    InMux I__1108 (
            .O(N__5952),
            .I(N__5949));
    LocalMux I__1107 (
            .O(N__5949),
            .I(N__5943));
    InMux I__1106 (
            .O(N__5948),
            .I(N__5938));
    InMux I__1105 (
            .O(N__5947),
            .I(N__5938));
    InMux I__1104 (
            .O(N__5946),
            .I(N__5934));
    Span4Mux_h I__1103 (
            .O(N__5943),
            .I(N__5931));
    LocalMux I__1102 (
            .O(N__5938),
            .I(N__5928));
    InMux I__1101 (
            .O(N__5937),
            .I(N__5925));
    LocalMux I__1100 (
            .O(N__5934),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__1099 (
            .O(N__5931),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__1098 (
            .O(N__5928),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__1097 (
            .O(N__5925),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__1096 (
            .O(N__5916),
            .I(N__5913));
    LocalMux I__1095 (
            .O(N__5913),
            .I(N__5908));
    InMux I__1094 (
            .O(N__5912),
            .I(N__5903));
    InMux I__1093 (
            .O(N__5911),
            .I(N__5903));
    Span4Mux_h I__1092 (
            .O(N__5908),
            .I(N__5897));
    LocalMux I__1091 (
            .O(N__5903),
            .I(N__5897));
    InMux I__1090 (
            .O(N__5902),
            .I(N__5894));
    Odrv4 I__1089 (
            .O(N__5897),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__1088 (
            .O(N__5894),
            .I(U712_REG_SM_DBR_SYNC_1));
    InMux I__1087 (
            .O(N__5889),
            .I(N__5885));
    IoInMux I__1086 (
            .O(N__5888),
            .I(N__5882));
    LocalMux I__1085 (
            .O(N__5885),
            .I(N__5879));
    LocalMux I__1084 (
            .O(N__5882),
            .I(N__5876));
    Sp12to4 I__1083 (
            .O(N__5879),
            .I(N__5873));
    Span4Mux_s3_h I__1082 (
            .O(N__5876),
            .I(N__5870));
    Span12Mux_v I__1081 (
            .O(N__5873),
            .I(N__5867));
    Sp12to4 I__1080 (
            .O(N__5870),
            .I(N__5864));
    Span12Mux_h I__1079 (
            .O(N__5867),
            .I(N__5861));
    Span12Mux_v I__1078 (
            .O(N__5864),
            .I(N__5858));
    Odrv12 I__1077 (
            .O(N__5861),
            .I(C1_c));
    Odrv12 I__1076 (
            .O(N__5858),
            .I(C1_c));
    InMux I__1075 (
            .O(N__5853),
            .I(N__5849));
    InMux I__1074 (
            .O(N__5852),
            .I(N__5846));
    LocalMux I__1073 (
            .O(N__5849),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1072 (
            .O(N__5846),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__1071 (
            .O(N__5841),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_ ));
    CascadeMux I__1070 (
            .O(N__5838),
            .I(N__5835));
    InMux I__1069 (
            .O(N__5835),
            .I(N__5832));
    LocalMux I__1068 (
            .O(N__5832),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2 ));
    InMux I__1067 (
            .O(N__5829),
            .I(N__5822));
    InMux I__1066 (
            .O(N__5828),
            .I(N__5822));
    InMux I__1065 (
            .O(N__5827),
            .I(N__5819));
    LocalMux I__1064 (
            .O(N__5822),
            .I(N__5816));
    LocalMux I__1063 (
            .O(N__5819),
            .I(N__5813));
    Span4Mux_h I__1062 (
            .O(N__5816),
            .I(N__5810));
    Odrv4 I__1061 (
            .O(N__5813),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3 ));
    Odrv4 I__1060 (
            .O(N__5810),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3 ));
    CascadeMux I__1059 (
            .O(N__5805),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_ ));
    CascadeMux I__1058 (
            .O(N__5802),
            .I(N__5799));
    InMux I__1057 (
            .O(N__5799),
            .I(N__5792));
    InMux I__1056 (
            .O(N__5798),
            .I(N__5786));
    InMux I__1055 (
            .O(N__5797),
            .I(N__5786));
    CascadeMux I__1054 (
            .O(N__5796),
            .I(N__5779));
    InMux I__1053 (
            .O(N__5795),
            .I(N__5775));
    LocalMux I__1052 (
            .O(N__5792),
            .I(N__5772));
    InMux I__1051 (
            .O(N__5791),
            .I(N__5769));
    LocalMux I__1050 (
            .O(N__5786),
            .I(N__5766));
    InMux I__1049 (
            .O(N__5785),
            .I(N__5757));
    InMux I__1048 (
            .O(N__5784),
            .I(N__5757));
    InMux I__1047 (
            .O(N__5783),
            .I(N__5757));
    InMux I__1046 (
            .O(N__5782),
            .I(N__5757));
    InMux I__1045 (
            .O(N__5779),
            .I(N__5752));
    InMux I__1044 (
            .O(N__5778),
            .I(N__5752));
    LocalMux I__1043 (
            .O(N__5775),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1042 (
            .O(N__5772),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1041 (
            .O(N__5769),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1040 (
            .O(N__5766),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1039 (
            .O(N__5757),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1038 (
            .O(N__5752),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1037 (
            .O(N__5739),
            .I(N__5736));
    InMux I__1036 (
            .O(N__5736),
            .I(N__5733));
    LocalMux I__1035 (
            .O(N__5733),
            .I(N__5730));
    Odrv4 I__1034 (
            .O(N__5730),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3 ));
    InMux I__1033 (
            .O(N__5727),
            .I(N__5718));
    InMux I__1032 (
            .O(N__5726),
            .I(N__5718));
    InMux I__1031 (
            .O(N__5725),
            .I(N__5718));
    LocalMux I__1030 (
            .O(N__5718),
            .I(\U712_CHIP_RAM.N_52 ));
    InMux I__1029 (
            .O(N__5715),
            .I(N__5712));
    LocalMux I__1028 (
            .O(N__5712),
            .I(N__5704));
    InMux I__1027 (
            .O(N__5711),
            .I(N__5701));
    InMux I__1026 (
            .O(N__5710),
            .I(N__5696));
    InMux I__1025 (
            .O(N__5709),
            .I(N__5691));
    InMux I__1024 (
            .O(N__5708),
            .I(N__5691));
    InMux I__1023 (
            .O(N__5707),
            .I(N__5688));
    Span4Mux_h I__1022 (
            .O(N__5704),
            .I(N__5683));
    LocalMux I__1021 (
            .O(N__5701),
            .I(N__5683));
    InMux I__1020 (
            .O(N__5700),
            .I(N__5680));
    InMux I__1019 (
            .O(N__5699),
            .I(N__5666));
    LocalMux I__1018 (
            .O(N__5696),
            .I(N__5661));
    LocalMux I__1017 (
            .O(N__5691),
            .I(N__5661));
    LocalMux I__1016 (
            .O(N__5688),
            .I(N__5654));
    Span4Mux_v I__1015 (
            .O(N__5683),
            .I(N__5654));
    LocalMux I__1014 (
            .O(N__5680),
            .I(N__5654));
    InMux I__1013 (
            .O(N__5679),
            .I(N__5647));
    InMux I__1012 (
            .O(N__5678),
            .I(N__5647));
    InMux I__1011 (
            .O(N__5677),
            .I(N__5647));
    InMux I__1010 (
            .O(N__5676),
            .I(N__5638));
    InMux I__1009 (
            .O(N__5675),
            .I(N__5638));
    InMux I__1008 (
            .O(N__5674),
            .I(N__5638));
    InMux I__1007 (
            .O(N__5673),
            .I(N__5638));
    InMux I__1006 (
            .O(N__5672),
            .I(N__5631));
    InMux I__1005 (
            .O(N__5671),
            .I(N__5631));
    InMux I__1004 (
            .O(N__5670),
            .I(N__5631));
    InMux I__1003 (
            .O(N__5669),
            .I(N__5628));
    LocalMux I__1002 (
            .O(N__5666),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1001 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1000 (
            .O(N__5654),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__999 (
            .O(N__5647),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__998 (
            .O(N__5638),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__997 (
            .O(N__5631),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__996 (
            .O(N__5628),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__995 (
            .O(N__5613),
            .I(N__5610));
    InMux I__994 (
            .O(N__5610),
            .I(N__5604));
    InMux I__993 (
            .O(N__5609),
            .I(N__5600));
    InMux I__992 (
            .O(N__5608),
            .I(N__5594));
    InMux I__991 (
            .O(N__5607),
            .I(N__5594));
    LocalMux I__990 (
            .O(N__5604),
            .I(N__5591));
    CascadeMux I__989 (
            .O(N__5603),
            .I(N__5587));
    LocalMux I__988 (
            .O(N__5600),
            .I(N__5583));
    CascadeMux I__987 (
            .O(N__5599),
            .I(N__5579));
    LocalMux I__986 (
            .O(N__5594),
            .I(N__5568));
    Span4Mux_h I__985 (
            .O(N__5591),
            .I(N__5568));
    InMux I__984 (
            .O(N__5590),
            .I(N__5565));
    InMux I__983 (
            .O(N__5587),
            .I(N__5560));
    InMux I__982 (
            .O(N__5586),
            .I(N__5560));
    Span4Mux_h I__981 (
            .O(N__5583),
            .I(N__5557));
    InMux I__980 (
            .O(N__5582),
            .I(N__5548));
    InMux I__979 (
            .O(N__5579),
            .I(N__5548));
    InMux I__978 (
            .O(N__5578),
            .I(N__5548));
    InMux I__977 (
            .O(N__5577),
            .I(N__5548));
    InMux I__976 (
            .O(N__5576),
            .I(N__5543));
    InMux I__975 (
            .O(N__5575),
            .I(N__5543));
    InMux I__974 (
            .O(N__5574),
            .I(N__5540));
    InMux I__973 (
            .O(N__5573),
            .I(N__5537));
    Odrv4 I__972 (
            .O(N__5568),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__971 (
            .O(N__5565),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__970 (
            .O(N__5560),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__969 (
            .O(N__5557),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__968 (
            .O(N__5548),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__967 (
            .O(N__5543),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__966 (
            .O(N__5540),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__965 (
            .O(N__5537),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__964 (
            .O(N__5520),
            .I(N__5515));
    CascadeMux I__963 (
            .O(N__5519),
            .I(N__5511));
    CascadeMux I__962 (
            .O(N__5518),
            .I(N__5506));
    InMux I__961 (
            .O(N__5515),
            .I(N__5498));
    InMux I__960 (
            .O(N__5514),
            .I(N__5495));
    InMux I__959 (
            .O(N__5511),
            .I(N__5488));
    InMux I__958 (
            .O(N__5510),
            .I(N__5488));
    InMux I__957 (
            .O(N__5509),
            .I(N__5488));
    InMux I__956 (
            .O(N__5506),
            .I(N__5485));
    InMux I__955 (
            .O(N__5505),
            .I(N__5480));
    InMux I__954 (
            .O(N__5504),
            .I(N__5480));
    InMux I__953 (
            .O(N__5503),
            .I(N__5473));
    InMux I__952 (
            .O(N__5502),
            .I(N__5473));
    InMux I__951 (
            .O(N__5501),
            .I(N__5473));
    LocalMux I__950 (
            .O(N__5498),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__949 (
            .O(N__5495),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__948 (
            .O(N__5488),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__947 (
            .O(N__5485),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__946 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__945 (
            .O(N__5473),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__944 (
            .O(N__5460),
            .I(N__5456));
    InMux I__943 (
            .O(N__5459),
            .I(N__5453));
    LocalMux I__942 (
            .O(N__5456),
            .I(N__5450));
    LocalMux I__941 (
            .O(N__5453),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv12 I__940 (
            .O(N__5450),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__939 (
            .O(N__5445),
            .I(N__5442));
    LocalMux I__938 (
            .O(N__5442),
            .I(N__5439));
    Odrv12 I__937 (
            .O(N__5439),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__936 (
            .O(N__5436),
            .I(N__5433));
    InMux I__935 (
            .O(N__5433),
            .I(N__5430));
    LocalMux I__934 (
            .O(N__5430),
            .I(N__5426));
    InMux I__933 (
            .O(N__5429),
            .I(N__5423));
    Span4Mux_h I__932 (
            .O(N__5426),
            .I(N__5420));
    LocalMux I__931 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__930 (
            .O(N__5420),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__929 (
            .O(N__5415),
            .I(N__5412));
    LocalMux I__928 (
            .O(N__5412),
            .I(N__5409));
    Odrv12 I__927 (
            .O(N__5409),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__926 (
            .O(N__5406),
            .I(N__5403));
    LocalMux I__925 (
            .O(N__5403),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__924 (
            .O(N__5400),
            .I(N__5397));
    LocalMux I__923 (
            .O(N__5397),
            .I(N__5394));
    Span4Mux_h I__922 (
            .O(N__5394),
            .I(N__5389));
    InMux I__921 (
            .O(N__5393),
            .I(N__5384));
    InMux I__920 (
            .O(N__5392),
            .I(N__5384));
    Odrv4 I__919 (
            .O(N__5389),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__918 (
            .O(N__5384),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    InMux I__917 (
            .O(N__5379),
            .I(N__5376));
    LocalMux I__916 (
            .O(N__5376),
            .I(N__5372));
    InMux I__915 (
            .O(N__5375),
            .I(N__5369));
    Span4Mux_v I__914 (
            .O(N__5372),
            .I(N__5366));
    LocalMux I__913 (
            .O(N__5369),
            .I(N__5363));
    Span4Mux_v I__912 (
            .O(N__5366),
            .I(N__5360));
    Span4Mux_v I__911 (
            .O(N__5363),
            .I(N__5357));
    Sp12to4 I__910 (
            .O(N__5360),
            .I(N__5352));
    Sp12to4 I__909 (
            .O(N__5357),
            .I(N__5352));
    Span12Mux_h I__908 (
            .O(N__5352),
            .I(N__5349));
    Span12Mux_v I__907 (
            .O(N__5349),
            .I(N__5346));
    Odrv12 I__906 (
            .O(N__5346),
            .I(TSn_c));
    CascadeMux I__905 (
            .O(N__5343),
            .I(N__5340));
    InMux I__904 (
            .O(N__5340),
            .I(N__5337));
    LocalMux I__903 (
            .O(N__5337),
            .I(N__5334));
    Span4Mux_v I__902 (
            .O(N__5334),
            .I(N__5331));
    Span4Mux_h I__901 (
            .O(N__5331),
            .I(N__5327));
    IoInMux I__900 (
            .O(N__5330),
            .I(N__5324));
    Sp12to4 I__899 (
            .O(N__5327),
            .I(N__5321));
    LocalMux I__898 (
            .O(N__5324),
            .I(N__5318));
    Span12Mux_v I__897 (
            .O(N__5321),
            .I(N__5315));
    IoSpan4Mux I__896 (
            .O(N__5318),
            .I(N__5312));
    Odrv12 I__895 (
            .O(N__5315),
            .I(RAMENn_c));
    Odrv4 I__894 (
            .O(N__5312),
            .I(RAMENn_c));
    InMux I__893 (
            .O(N__5307),
            .I(N__5303));
    InMux I__892 (
            .O(N__5306),
            .I(N__5297));
    LocalMux I__891 (
            .O(N__5303),
            .I(N__5294));
    InMux I__890 (
            .O(N__5302),
            .I(N__5289));
    InMux I__889 (
            .O(N__5301),
            .I(N__5289));
    InMux I__888 (
            .O(N__5300),
            .I(N__5286));
    LocalMux I__887 (
            .O(N__5297),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__886 (
            .O(N__5294),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__885 (
            .O(N__5289),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__884 (
            .O(N__5286),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__883 (
            .O(N__5277),
            .I(N__5274));
    LocalMux I__882 (
            .O(N__5274),
            .I(N__5270));
    InMux I__881 (
            .O(N__5273),
            .I(N__5267));
    Odrv4 I__880 (
            .O(N__5270),
            .I(\U712_CHIP_RAM.N_492 ));
    LocalMux I__879 (
            .O(N__5267),
            .I(\U712_CHIP_RAM.N_492 ));
    CascadeMux I__878 (
            .O(N__5262),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_ ));
    InMux I__877 (
            .O(N__5259),
            .I(N__5256));
    LocalMux I__876 (
            .O(N__5256),
            .I(N__5252));
    InMux I__875 (
            .O(N__5255),
            .I(N__5249));
    Odrv4 I__874 (
            .O(N__5252),
            .I(\U712_CHIP_RAM.N_331 ));
    LocalMux I__873 (
            .O(N__5249),
            .I(\U712_CHIP_RAM.N_331 ));
    InMux I__872 (
            .O(N__5244),
            .I(N__5237));
    InMux I__871 (
            .O(N__5243),
            .I(N__5237));
    InMux I__870 (
            .O(N__5242),
            .I(N__5234));
    LocalMux I__869 (
            .O(N__5237),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    LocalMux I__868 (
            .O(N__5234),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    InMux I__867 (
            .O(N__5229),
            .I(N__5226));
    LocalMux I__866 (
            .O(N__5226),
            .I(\U712_CHIP_RAM.N_222 ));
    CascadeMux I__865 (
            .O(N__5223),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ));
    InMux I__864 (
            .O(N__5220),
            .I(N__5214));
    InMux I__863 (
            .O(N__5219),
            .I(N__5209));
    InMux I__862 (
            .O(N__5218),
            .I(N__5209));
    InMux I__861 (
            .O(N__5217),
            .I(N__5204));
    LocalMux I__860 (
            .O(N__5214),
            .I(N__5199));
    LocalMux I__859 (
            .O(N__5209),
            .I(N__5199));
    InMux I__858 (
            .O(N__5208),
            .I(N__5194));
    InMux I__857 (
            .O(N__5207),
            .I(N__5194));
    LocalMux I__856 (
            .O(N__5204),
            .I(\U712_CHIP_RAM.N_332 ));
    Odrv4 I__855 (
            .O(N__5199),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__854 (
            .O(N__5194),
            .I(\U712_CHIP_RAM.N_332 ));
    CascadeMux I__853 (
            .O(N__5187),
            .I(N__5182));
    InMux I__852 (
            .O(N__5186),
            .I(N__5175));
    InMux I__851 (
            .O(N__5185),
            .I(N__5172));
    InMux I__850 (
            .O(N__5182),
            .I(N__5169));
    InMux I__849 (
            .O(N__5181),
            .I(N__5166));
    InMux I__848 (
            .O(N__5180),
            .I(N__5163));
    InMux I__847 (
            .O(N__5179),
            .I(N__5158));
    InMux I__846 (
            .O(N__5178),
            .I(N__5158));
    LocalMux I__845 (
            .O(N__5175),
            .I(N__5153));
    LocalMux I__844 (
            .O(N__5172),
            .I(N__5153));
    LocalMux I__843 (
            .O(N__5169),
            .I(\U712_CHIP_RAM.N_346 ));
    LocalMux I__842 (
            .O(N__5166),
            .I(\U712_CHIP_RAM.N_346 ));
    LocalMux I__841 (
            .O(N__5163),
            .I(\U712_CHIP_RAM.N_346 ));
    LocalMux I__840 (
            .O(N__5158),
            .I(\U712_CHIP_RAM.N_346 ));
    Odrv4 I__839 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.N_346 ));
    CascadeMux I__838 (
            .O(N__5142),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_ ));
    InMux I__837 (
            .O(N__5139),
            .I(N__5136));
    LocalMux I__836 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0 ));
    CascadeMux I__835 (
            .O(N__5133),
            .I(N__5127));
    InMux I__834 (
            .O(N__5132),
            .I(N__5124));
    CascadeMux I__833 (
            .O(N__5131),
            .I(N__5120));
    InMux I__832 (
            .O(N__5130),
            .I(N__5116));
    InMux I__831 (
            .O(N__5127),
            .I(N__5113));
    LocalMux I__830 (
            .O(N__5124),
            .I(N__5110));
    InMux I__829 (
            .O(N__5123),
            .I(N__5105));
    InMux I__828 (
            .O(N__5120),
            .I(N__5105));
    InMux I__827 (
            .O(N__5119),
            .I(N__5102));
    LocalMux I__826 (
            .O(N__5116),
            .I(\U712_CHIP_RAM.N_330 ));
    LocalMux I__825 (
            .O(N__5113),
            .I(\U712_CHIP_RAM.N_330 ));
    Odrv4 I__824 (
            .O(N__5110),
            .I(\U712_CHIP_RAM.N_330 ));
    LocalMux I__823 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.N_330 ));
    LocalMux I__822 (
            .O(N__5102),
            .I(\U712_CHIP_RAM.N_330 ));
    InMux I__821 (
            .O(N__5091),
            .I(N__5088));
    LocalMux I__820 (
            .O(N__5088),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0 ));
    InMux I__819 (
            .O(N__5085),
            .I(N__5082));
    LocalMux I__818 (
            .O(N__5082),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0 ));
    CascadeMux I__817 (
            .O(N__5079),
            .I(N__5076));
    InMux I__816 (
            .O(N__5076),
            .I(N__5073));
    LocalMux I__815 (
            .O(N__5073),
            .I(\U712_REG_SM.N_71 ));
    IoInMux I__814 (
            .O(N__5070),
            .I(N__5067));
    LocalMux I__813 (
            .O(N__5067),
            .I(N__5064));
    Odrv12 I__812 (
            .O(N__5064),
            .I(CMA_c_2));
    IoInMux I__811 (
            .O(N__5061),
            .I(N__5058));
    LocalMux I__810 (
            .O(N__5058),
            .I(N__5055));
    Span4Mux_s3_v I__809 (
            .O(N__5055),
            .I(N__5052));
    Span4Mux_v I__808 (
            .O(N__5052),
            .I(N__5049));
    Span4Mux_h I__807 (
            .O(N__5049),
            .I(N__5046));
    Odrv4 I__806 (
            .O(N__5046),
            .I(CONSTANT_ONE_NET));
    InMux I__805 (
            .O(N__5043),
            .I(N__5040));
    LocalMux I__804 (
            .O(N__5040),
            .I(N__5037));
    Span4Mux_v I__803 (
            .O(N__5037),
            .I(N__5034));
    Sp12to4 I__802 (
            .O(N__5034),
            .I(N__5031));
    Span12Mux_h I__801 (
            .O(N__5031),
            .I(N__5028));
    Odrv12 I__800 (
            .O(N__5028),
            .I(A_c_11));
    CascadeMux I__799 (
            .O(N__5025),
            .I(N__5022));
    InMux I__798 (
            .O(N__5022),
            .I(N__5019));
    LocalMux I__797 (
            .O(N__5019),
            .I(N__5016));
    Span4Mux_v I__796 (
            .O(N__5016),
            .I(N__5013));
    Sp12to4 I__795 (
            .O(N__5013),
            .I(N__5010));
    Span12Mux_h I__794 (
            .O(N__5010),
            .I(N__5007));
    Span12Mux_v I__793 (
            .O(N__5007),
            .I(N__5004));
    Odrv12 I__792 (
            .O(N__5004),
            .I(A_c_4));
    InMux I__791 (
            .O(N__5001),
            .I(N__4998));
    LocalMux I__790 (
            .O(N__4998),
            .I(\U712_CHIP_RAM.N_369 ));
    InMux I__789 (
            .O(N__4995),
            .I(N__4992));
    LocalMux I__788 (
            .O(N__4992),
            .I(\U712_CHIP_RAM.N_445 ));
    InMux I__787 (
            .O(N__4989),
            .I(N__4986));
    LocalMux I__786 (
            .O(N__4986),
            .I(N__4983));
    Span4Mux_v I__785 (
            .O(N__4983),
            .I(N__4980));
    Sp12to4 I__784 (
            .O(N__4980),
            .I(N__4977));
    Span12Mux_h I__783 (
            .O(N__4977),
            .I(N__4974));
    Odrv12 I__782 (
            .O(N__4974),
            .I(A_c_12));
    InMux I__781 (
            .O(N__4971),
            .I(N__4968));
    LocalMux I__780 (
            .O(N__4968),
            .I(N__4965));
    Sp12to4 I__779 (
            .O(N__4965),
            .I(N__4962));
    Span12Mux_v I__778 (
            .O(N__4962),
            .I(N__4959));
    Span12Mux_h I__777 (
            .O(N__4959),
            .I(N__4956));
    Odrv12 I__776 (
            .O(N__4956),
            .I(A_c_5));
    SRMux I__775 (
            .O(N__4953),
            .I(N__4950));
    LocalMux I__774 (
            .O(N__4950),
            .I(N__4947));
    Span4Mux_h I__773 (
            .O(N__4947),
            .I(N__4944));
    Span4Mux_h I__772 (
            .O(N__4944),
            .I(N__4941));
    Odrv4 I__771 (
            .O(N__4941),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__770 (
            .O(N__4938),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    InMux I__769 (
            .O(N__4935),
            .I(N__4931));
    InMux I__768 (
            .O(N__4934),
            .I(N__4928));
    LocalMux I__767 (
            .O(N__4931),
            .I(\U712_REG_SM.N_338 ));
    LocalMux I__766 (
            .O(N__4928),
            .I(\U712_REG_SM.N_338 ));
    CascadeMux I__765 (
            .O(N__4923),
            .I(\U712_REG_SM.N_338_cascade_ ));
    CascadeMux I__764 (
            .O(N__4920),
            .I(\U712_REG_SM.N_354_cascade_ ));
    CascadeMux I__763 (
            .O(N__4917),
            .I(N__4914));
    InMux I__762 (
            .O(N__4914),
            .I(N__4911));
    LocalMux I__761 (
            .O(N__4911),
            .I(N__4908));
    Span4Mux_v I__760 (
            .O(N__4908),
            .I(N__4905));
    Sp12to4 I__759 (
            .O(N__4905),
            .I(N__4902));
    Span12Mux_h I__758 (
            .O(N__4902),
            .I(N__4899));
    Span12Mux_v I__757 (
            .O(N__4899),
            .I(N__4896));
    Odrv12 I__756 (
            .O(N__4896),
            .I(REGSPACEn_c));
    CascadeMux I__755 (
            .O(N__4893),
            .I(N__4889));
    InMux I__754 (
            .O(N__4892),
            .I(N__4885));
    InMux I__753 (
            .O(N__4889),
            .I(N__4880));
    InMux I__752 (
            .O(N__4888),
            .I(N__4880));
    LocalMux I__751 (
            .O(N__4885),
            .I(N__4877));
    LocalMux I__750 (
            .O(N__4880),
            .I(N__4874));
    Span4Mux_v I__749 (
            .O(N__4877),
            .I(N__4871));
    Span12Mux_v I__748 (
            .O(N__4874),
            .I(N__4868));
    Sp12to4 I__747 (
            .O(N__4871),
            .I(N__4865));
    Span12Mux_h I__746 (
            .O(N__4868),
            .I(N__4862));
    Span12Mux_h I__745 (
            .O(N__4865),
            .I(N__4859));
    Span12Mux_v I__744 (
            .O(N__4862),
            .I(N__4856));
    Span12Mux_v I__743 (
            .O(N__4859),
            .I(N__4853));
    Odrv12 I__742 (
            .O(N__4856),
            .I(CASUn_c));
    Odrv12 I__741 (
            .O(N__4853),
            .I(CASUn_c));
    CascadeMux I__740 (
            .O(N__4848),
            .I(N__4845));
    InMux I__739 (
            .O(N__4845),
            .I(N__4839));
    InMux I__738 (
            .O(N__4844),
            .I(N__4839));
    LocalMux I__737 (
            .O(N__4839),
            .I(N__4835));
    InMux I__736 (
            .O(N__4838),
            .I(N__4832));
    Span4Mux_v I__735 (
            .O(N__4835),
            .I(N__4829));
    LocalMux I__734 (
            .O(N__4832),
            .I(N__4826));
    Sp12to4 I__733 (
            .O(N__4829),
            .I(N__4823));
    Sp12to4 I__732 (
            .O(N__4826),
            .I(N__4820));
    Span12Mux_h I__731 (
            .O(N__4823),
            .I(N__4817));
    Span12Mux_v I__730 (
            .O(N__4820),
            .I(N__4814));
    Span12Mux_v I__729 (
            .O(N__4817),
            .I(N__4809));
    Span12Mux_h I__728 (
            .O(N__4814),
            .I(N__4809));
    Odrv12 I__727 (
            .O(N__4809),
            .I(CASLn_c));
    InMux I__726 (
            .O(N__4806),
            .I(N__4803));
    LocalMux I__725 (
            .O(N__4803),
            .I(\U712_REG_SM.N_431 ));
    InMux I__724 (
            .O(N__4800),
            .I(N__4796));
    InMux I__723 (
            .O(N__4799),
            .I(N__4793));
    LocalMux I__722 (
            .O(N__4796),
            .I(\U712_REG_SM.N_358 ));
    LocalMux I__721 (
            .O(N__4793),
            .I(\U712_REG_SM.N_358 ));
    InMux I__720 (
            .O(N__4788),
            .I(N__4783));
    InMux I__719 (
            .O(N__4787),
            .I(N__4780));
    InMux I__718 (
            .O(N__4786),
            .I(N__4777));
    LocalMux I__717 (
            .O(N__4783),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__716 (
            .O(N__4780),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__715 (
            .O(N__4777),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__714 (
            .O(N__4770),
            .I(\U712_CHIP_RAM.N_341_cascade_ ));
    InMux I__713 (
            .O(N__4767),
            .I(N__4763));
    InMux I__712 (
            .O(N__4766),
            .I(N__4760));
    LocalMux I__711 (
            .O(N__4763),
            .I(\U712_CHIP_RAM.N_560 ));
    LocalMux I__710 (
            .O(N__4760),
            .I(\U712_CHIP_RAM.N_560 ));
    CascadeMux I__709 (
            .O(N__4755),
            .I(\U712_CHIP_RAM.N_450_cascade_ ));
    CascadeMux I__708 (
            .O(N__4752),
            .I(\U712_CHIP_RAM.N_326_cascade_ ));
    InMux I__707 (
            .O(N__4749),
            .I(N__4743));
    InMux I__706 (
            .O(N__4748),
            .I(N__4743));
    LocalMux I__705 (
            .O(N__4743),
            .I(\U712_CHIP_RAM.N_326 ));
    IoInMux I__704 (
            .O(N__4740),
            .I(N__4737));
    LocalMux I__703 (
            .O(N__4737),
            .I(N__4734));
    Span4Mux_s3_v I__702 (
            .O(N__4734),
            .I(N__4731));
    Span4Mux_h I__701 (
            .O(N__4731),
            .I(N__4724));
    InMux I__700 (
            .O(N__4730),
            .I(N__4719));
    InMux I__699 (
            .O(N__4729),
            .I(N__4719));
    InMux I__698 (
            .O(N__4728),
            .I(N__4714));
    InMux I__697 (
            .O(N__4727),
            .I(N__4714));
    Sp12to4 I__696 (
            .O(N__4724),
            .I(N__4711));
    LocalMux I__695 (
            .O(N__4719),
            .I(N__4708));
    LocalMux I__694 (
            .O(N__4714),
            .I(N__4705));
    Span12Mux_v I__693 (
            .O(N__4711),
            .I(N__4701));
    Span4Mux_v I__692 (
            .O(N__4708),
            .I(N__4696));
    Span4Mux_v I__691 (
            .O(N__4705),
            .I(N__4696));
    InMux I__690 (
            .O(N__4704),
            .I(N__4693));
    Odrv12 I__689 (
            .O(N__4701),
            .I(DBENn_c));
    Odrv4 I__688 (
            .O(N__4696),
            .I(DBENn_c));
    LocalMux I__687 (
            .O(N__4693),
            .I(DBENn_c));
    InMux I__686 (
            .O(N__4686),
            .I(N__4682));
    InMux I__685 (
            .O(N__4685),
            .I(N__4679));
    LocalMux I__684 (
            .O(N__4682),
            .I(\U712_CHIP_RAM.N_450 ));
    LocalMux I__683 (
            .O(N__4679),
            .I(\U712_CHIP_RAM.N_450 ));
    InMux I__682 (
            .O(N__4674),
            .I(N__4670));
    InMux I__681 (
            .O(N__4673),
            .I(N__4667));
    LocalMux I__680 (
            .O(N__4670),
            .I(N__4664));
    LocalMux I__679 (
            .O(N__4667),
            .I(N__4661));
    Span4Mux_v I__678 (
            .O(N__4664),
            .I(N__4658));
    Span4Mux_v I__677 (
            .O(N__4661),
            .I(N__4655));
    Sp12to4 I__676 (
            .O(N__4658),
            .I(N__4650));
    Sp12to4 I__675 (
            .O(N__4655),
            .I(N__4650));
    Span12Mux_h I__674 (
            .O(N__4650),
            .I(N__4647));
    Span12Mux_v I__673 (
            .O(N__4647),
            .I(N__4644));
    Odrv12 I__672 (
            .O(N__4644),
            .I(AWEn_c));
    InMux I__671 (
            .O(N__4641),
            .I(N__4637));
    InMux I__670 (
            .O(N__4640),
            .I(N__4634));
    LocalMux I__669 (
            .O(N__4637),
            .I(N__4627));
    LocalMux I__668 (
            .O(N__4634),
            .I(N__4627));
    InMux I__667 (
            .O(N__4633),
            .I(N__4622));
    InMux I__666 (
            .O(N__4632),
            .I(N__4622));
    Span4Mux_v I__665 (
            .O(N__4627),
            .I(N__4617));
    LocalMux I__664 (
            .O(N__4622),
            .I(N__4617));
    Odrv4 I__663 (
            .O(N__4617),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CEMux I__662 (
            .O(N__4614),
            .I(N__4611));
    LocalMux I__661 (
            .O(N__4611),
            .I(N__4608));
    Odrv4 I__660 (
            .O(N__4608),
            .I(\U712_CHIP_RAM.N_450_0 ));
    CascadeMux I__659 (
            .O(N__4605),
            .I(N__4601));
    InMux I__658 (
            .O(N__4604),
            .I(N__4596));
    InMux I__657 (
            .O(N__4601),
            .I(N__4596));
    LocalMux I__656 (
            .O(N__4596),
            .I(\U712_CHIP_RAM.DMA_CYCLE_7 ));
    InMux I__655 (
            .O(N__4593),
            .I(N__4590));
    LocalMux I__654 (
            .O(N__4590),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0 ));
    CascadeMux I__653 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.N_332_cascade_ ));
    InMux I__652 (
            .O(N__4584),
            .I(N__4578));
    InMux I__651 (
            .O(N__4583),
            .I(N__4575));
    InMux I__650 (
            .O(N__4582),
            .I(N__4570));
    InMux I__649 (
            .O(N__4581),
            .I(N__4570));
    LocalMux I__648 (
            .O(N__4578),
            .I(\U712_CHIP_RAM.N_493 ));
    LocalMux I__647 (
            .O(N__4575),
            .I(\U712_CHIP_RAM.N_493 ));
    LocalMux I__646 (
            .O(N__4570),
            .I(\U712_CHIP_RAM.N_493 ));
    CascadeMux I__645 (
            .O(N__4563),
            .I(N__4560));
    InMux I__644 (
            .O(N__4560),
            .I(N__4556));
    InMux I__643 (
            .O(N__4559),
            .I(N__4551));
    LocalMux I__642 (
            .O(N__4556),
            .I(N__4548));
    InMux I__641 (
            .O(N__4555),
            .I(N__4545));
    InMux I__640 (
            .O(N__4554),
            .I(N__4542));
    LocalMux I__639 (
            .O(N__4551),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    Odrv4 I__638 (
            .O(N__4548),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__637 (
            .O(N__4545),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__636 (
            .O(N__4542),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__635 (
            .O(N__4533),
            .I(N__4528));
    InMux I__634 (
            .O(N__4532),
            .I(N__4525));
    InMux I__633 (
            .O(N__4531),
            .I(N__4522));
    LocalMux I__632 (
            .O(N__4528),
            .I(N__4517));
    LocalMux I__631 (
            .O(N__4525),
            .I(N__4517));
    LocalMux I__630 (
            .O(N__4522),
            .I(\U712_CHIP_RAM.N_351 ));
    Odrv4 I__629 (
            .O(N__4517),
            .I(\U712_CHIP_RAM.N_351 ));
    CascadeMux I__628 (
            .O(N__4512),
            .I(\U712_CHIP_RAM.N_351_cascade_ ));
    InMux I__627 (
            .O(N__4509),
            .I(N__4504));
    InMux I__626 (
            .O(N__4508),
            .I(N__4501));
    InMux I__625 (
            .O(N__4507),
            .I(N__4498));
    LocalMux I__624 (
            .O(N__4504),
            .I(N__4487));
    LocalMux I__623 (
            .O(N__4501),
            .I(N__4487));
    LocalMux I__622 (
            .O(N__4498),
            .I(N__4487));
    InMux I__621 (
            .O(N__4497),
            .I(N__4478));
    InMux I__620 (
            .O(N__4496),
            .I(N__4478));
    InMux I__619 (
            .O(N__4495),
            .I(N__4478));
    InMux I__618 (
            .O(N__4494),
            .I(N__4478));
    Odrv4 I__617 (
            .O(N__4487),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__616 (
            .O(N__4478),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__615 (
            .O(N__4473),
            .I(N__4470));
    LocalMux I__614 (
            .O(N__4470),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1 ));
    InMux I__613 (
            .O(N__4467),
            .I(N__4464));
    LocalMux I__612 (
            .O(N__4464),
            .I(N__4461));
    Odrv4 I__611 (
            .O(N__4461),
            .I(\U712_CHIP_RAM.N_402 ));
    InMux I__610 (
            .O(N__4458),
            .I(N__4455));
    LocalMux I__609 (
            .O(N__4455),
            .I(\U712_CHIP_RAM.N_341 ));
    CascadeMux I__608 (
            .O(N__4452),
            .I(\U712_CHIP_RAM.N_471_cascade_ ));
    CascadeMux I__607 (
            .O(N__4449),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_ ));
    IoInMux I__606 (
            .O(N__4446),
            .I(N__4443));
    LocalMux I__605 (
            .O(N__4443),
            .I(N__4440));
    Span12Mux_s6_h I__604 (
            .O(N__4440),
            .I(N__4437));
    Span12Mux_h I__603 (
            .O(N__4437),
            .I(N__4433));
    InMux I__602 (
            .O(N__4436),
            .I(N__4430));
    Odrv12 I__601 (
            .O(N__4433),
            .I(CLK_EN_c));
    LocalMux I__600 (
            .O(N__4430),
            .I(CLK_EN_c));
    CascadeMux I__599 (
            .O(N__4425),
            .I(\U712_CHIP_RAM.N_447_cascade_ ));
    CascadeMux I__598 (
            .O(N__4422),
            .I(N__4416));
    InMux I__597 (
            .O(N__4421),
            .I(N__4413));
    InMux I__596 (
            .O(N__4420),
            .I(N__4410));
    InMux I__595 (
            .O(N__4419),
            .I(N__4407));
    InMux I__594 (
            .O(N__4416),
            .I(N__4404));
    LocalMux I__593 (
            .O(N__4413),
            .I(N__4401));
    LocalMux I__592 (
            .O(N__4410),
            .I(\U712_CHIP_RAM.N_333 ));
    LocalMux I__591 (
            .O(N__4407),
            .I(\U712_CHIP_RAM.N_333 ));
    LocalMux I__590 (
            .O(N__4404),
            .I(\U712_CHIP_RAM.N_333 ));
    Odrv4 I__589 (
            .O(N__4401),
            .I(\U712_CHIP_RAM.N_333 ));
    InMux I__588 (
            .O(N__4392),
            .I(N__4385));
    InMux I__587 (
            .O(N__4391),
            .I(N__4385));
    InMux I__586 (
            .O(N__4390),
            .I(N__4382));
    LocalMux I__585 (
            .O(N__4385),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__584 (
            .O(N__4382),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__583 (
            .O(N__4377),
            .I(N__4374));
    InMux I__582 (
            .O(N__4374),
            .I(N__4367));
    InMux I__581 (
            .O(N__4373),
            .I(N__4367));
    InMux I__580 (
            .O(N__4372),
            .I(N__4364));
    LocalMux I__579 (
            .O(N__4367),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__578 (
            .O(N__4364),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__577 (
            .O(N__4359),
            .I(N__4355));
    CascadeMux I__576 (
            .O(N__4358),
            .I(N__4351));
    InMux I__575 (
            .O(N__4355),
            .I(N__4346));
    InMux I__574 (
            .O(N__4354),
            .I(N__4346));
    InMux I__573 (
            .O(N__4351),
            .I(N__4343));
    LocalMux I__572 (
            .O(N__4346),
            .I(N__4338));
    LocalMux I__571 (
            .O(N__4343),
            .I(N__4338));
    Odrv4 I__570 (
            .O(N__4338),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__569 (
            .O(N__4335),
            .I(N__4332));
    InMux I__568 (
            .O(N__4332),
            .I(N__4328));
    InMux I__567 (
            .O(N__4331),
            .I(N__4325));
    LocalMux I__566 (
            .O(N__4328),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__565 (
            .O(N__4325),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__564 (
            .O(N__4320),
            .I(\U712_CHIP_RAM.N_330_cascade_ ));
    CascadeMux I__563 (
            .O(N__4317),
            .I(N__4314));
    InMux I__562 (
            .O(N__4314),
            .I(N__4311));
    LocalMux I__561 (
            .O(N__4311),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    InMux I__560 (
            .O(N__4308),
            .I(N__4305));
    LocalMux I__559 (
            .O(N__4305),
            .I(N__4301));
    InMux I__558 (
            .O(N__4304),
            .I(N__4298));
    Span4Mux_h I__557 (
            .O(N__4301),
            .I(N__4295));
    LocalMux I__556 (
            .O(N__4298),
            .I(CPU_TACKm));
    Odrv4 I__555 (
            .O(N__4295),
            .I(CPU_TACKm));
    CascadeMux I__554 (
            .O(N__4290),
            .I(\U712_CHIP_RAM.N_554_cascade_ ));
    InMux I__553 (
            .O(N__4287),
            .I(N__4284));
    LocalMux I__552 (
            .O(N__4284),
            .I(\U712_CHIP_RAM.N_565 ));
    CascadeMux I__551 (
            .O(N__4281),
            .I(\U712_CHIP_RAM.N_565_cascade_ ));
    InMux I__550 (
            .O(N__4278),
            .I(N__4275));
    LocalMux I__549 (
            .O(N__4275),
            .I(\U712_CHIP_RAM.N_563 ));
    CascadeMux I__548 (
            .O(N__4272),
            .I(\U712_CHIP_RAM.N_445_cascade_ ));
    InMux I__547 (
            .O(N__4269),
            .I(N__4266));
    LocalMux I__546 (
            .O(N__4266),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1 ));
    CascadeMux I__545 (
            .O(N__4263),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_ ));
    CascadeMux I__544 (
            .O(N__4260),
            .I(\U712_CHIP_RAM.N_333_cascade_ ));
    InMux I__543 (
            .O(N__4257),
            .I(N__4253));
    InMux I__542 (
            .O(N__4256),
            .I(N__4250));
    LocalMux I__541 (
            .O(N__4253),
            .I(\U712_CHIP_RAM.N_564 ));
    LocalMux I__540 (
            .O(N__4250),
            .I(\U712_CHIP_RAM.N_564 ));
    IoInMux I__539 (
            .O(N__4245),
            .I(N__4242));
    LocalMux I__538 (
            .O(N__4242),
            .I(N__4239));
    Span4Mux_s0_v I__537 (
            .O(N__4239),
            .I(N__4236));
    Span4Mux_h I__536 (
            .O(N__4236),
            .I(N__4233));
    Span4Mux_v I__535 (
            .O(N__4233),
            .I(N__4230));
    Span4Mux_v I__534 (
            .O(N__4230),
            .I(N__4227));
    Sp12to4 I__533 (
            .O(N__4227),
            .I(N__4224));
    Span12Mux_h I__532 (
            .O(N__4224),
            .I(N__4221));
    Odrv12 I__531 (
            .O(N__4221),
            .I(DRDENn_c));
    CascadeMux I__530 (
            .O(N__4218),
            .I(\U712_REG_SM.N_343_cascade_ ));
    CascadeMux I__529 (
            .O(N__4215),
            .I(\U712_REG_SM.N_358_cascade_ ));
    InMux I__528 (
            .O(N__4212),
            .I(N__4209));
    LocalMux I__527 (
            .O(N__4209),
            .I(N__4203));
    InMux I__526 (
            .O(N__4208),
            .I(N__4196));
    InMux I__525 (
            .O(N__4207),
            .I(N__4196));
    InMux I__524 (
            .O(N__4206),
            .I(N__4196));
    Odrv12 I__523 (
            .O(N__4203),
            .I(REG_CYCLEm));
    LocalMux I__522 (
            .O(N__4196),
            .I(REG_CYCLEm));
    CascadeMux I__521 (
            .O(N__4191),
            .I(N__4188));
    InMux I__520 (
            .O(N__4188),
            .I(N__4184));
    InMux I__519 (
            .O(N__4187),
            .I(N__4181));
    LocalMux I__518 (
            .O(N__4184),
            .I(REG_TACK));
    LocalMux I__517 (
            .O(N__4181),
            .I(REG_TACK));
    CascadeMux I__516 (
            .O(N__4176),
            .I(\U712_CHIP_RAM.N_563_cascade_ ));
    CascadeMux I__515 (
            .O(N__4173),
            .I(\U712_CHIP_RAM.N_215_cascade_ ));
    InMux I__514 (
            .O(N__4170),
            .I(N__4167));
    LocalMux I__513 (
            .O(N__4167),
            .I(N__4164));
    Span4Mux_h I__512 (
            .O(N__4164),
            .I(N__4161));
    Sp12to4 I__511 (
            .O(N__4161),
            .I(N__4158));
    Span12Mux_v I__510 (
            .O(N__4158),
            .I(N__4155));
    Odrv12 I__509 (
            .O(N__4155),
            .I(A_c_18));
    CascadeMux I__508 (
            .O(N__4152),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_ ));
    InMux I__507 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__506 (
            .O(N__4146),
            .I(N__4143));
    Sp12to4 I__505 (
            .O(N__4143),
            .I(N__4140));
    Span12Mux_v I__504 (
            .O(N__4140),
            .I(N__4137));
    Span12Mux_h I__503 (
            .O(N__4137),
            .I(N__4134));
    Odrv12 I__502 (
            .O(N__4134),
            .I(A_c_16));
    InMux I__501 (
            .O(N__4131),
            .I(N__4125));
    InMux I__500 (
            .O(N__4130),
            .I(N__4125));
    LocalMux I__499 (
            .O(N__4125),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0 ));
    CascadeMux I__498 (
            .O(N__4122),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_ ));
    InMux I__497 (
            .O(N__4119),
            .I(N__4116));
    LocalMux I__496 (
            .O(N__4116),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6 ));
    InMux I__495 (
            .O(N__4113),
            .I(N__4110));
    LocalMux I__494 (
            .O(N__4110),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ));
    IoInMux I__493 (
            .O(N__4107),
            .I(N__4104));
    LocalMux I__492 (
            .O(N__4104),
            .I(N__4101));
    Span4Mux_s1_v I__491 (
            .O(N__4101),
            .I(N__4098));
    Span4Mux_v I__490 (
            .O(N__4098),
            .I(N__4095));
    Span4Mux_v I__489 (
            .O(N__4095),
            .I(N__4092));
    Span4Mux_v I__488 (
            .O(N__4092),
            .I(N__4087));
    InMux I__487 (
            .O(N__4091),
            .I(N__4084));
    InMux I__486 (
            .O(N__4090),
            .I(N__4081));
    Odrv4 I__485 (
            .O(N__4087),
            .I(DBDIR_c));
    LocalMux I__484 (
            .O(N__4084),
            .I(DBDIR_c));
    LocalMux I__483 (
            .O(N__4081),
            .I(DBDIR_c));
    IoInMux I__482 (
            .O(N__4074),
            .I(N__4071));
    LocalMux I__481 (
            .O(N__4071),
            .I(N__4068));
    Span4Mux_s2_h I__480 (
            .O(N__4068),
            .I(N__4065));
    Span4Mux_v I__479 (
            .O(N__4065),
            .I(N__4062));
    Sp12to4 I__478 (
            .O(N__4062),
            .I(N__4059));
    Span12Mux_s11_h I__477 (
            .O(N__4059),
            .I(N__4056));
    Span12Mux_v I__476 (
            .O(N__4056),
            .I(N__4053));
    Odrv12 I__475 (
            .O(N__4053),
            .I(DRDDIR_i_0));
    InMux I__474 (
            .O(N__4050),
            .I(N__4046));
    InMux I__473 (
            .O(N__4049),
            .I(N__4043));
    LocalMux I__472 (
            .O(N__4046),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ));
    LocalMux I__471 (
            .O(N__4043),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ));
    CascadeMux I__470 (
            .O(N__4038),
            .I(\U712_BYTE_ENABLE.N_459_cascade_ ));
    InMux I__469 (
            .O(N__4035),
            .I(N__4032));
    LocalMux I__468 (
            .O(N__4032),
            .I(\U712_BYTE_ENABLE.N_352 ));
    IoInMux I__467 (
            .O(N__4029),
            .I(N__4026));
    LocalMux I__466 (
            .O(N__4026),
            .I(N__4023));
    Span12Mux_s4_v I__465 (
            .O(N__4023),
            .I(N__4020));
    Odrv12 I__464 (
            .O(N__4020),
            .I(N_47_i));
    CascadeMux I__463 (
            .O(N__4017),
            .I(N__4012));
    InMux I__462 (
            .O(N__4016),
            .I(N__4009));
    InMux I__461 (
            .O(N__4015),
            .I(N__4004));
    InMux I__460 (
            .O(N__4012),
            .I(N__4004));
    LocalMux I__459 (
            .O(N__4009),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__458 (
            .O(N__4004),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__457 (
            .O(N__3999),
            .I(N__3996));
    InMux I__456 (
            .O(N__3996),
            .I(N__3992));
    InMux I__455 (
            .O(N__3995),
            .I(N__3989));
    LocalMux I__454 (
            .O(N__3992),
            .I(N__3984));
    LocalMux I__453 (
            .O(N__3989),
            .I(N__3984));
    Odrv4 I__452 (
            .O(N__3984),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__451 (
            .O(N__3981),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__450 (
            .O(N__3978),
            .I(N__3973));
    InMux I__449 (
            .O(N__3977),
            .I(N__3970));
    InMux I__448 (
            .O(N__3976),
            .I(N__3967));
    LocalMux I__447 (
            .O(N__3973),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__446 (
            .O(N__3970),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__445 (
            .O(N__3967),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__444 (
            .O(N__3960),
            .I(\U712_CYCLE_TERM.N_362_i_0_en_cascade_ ));
    CEMux I__443 (
            .O(N__3957),
            .I(N__3954));
    LocalMux I__442 (
            .O(N__3954),
            .I(N__3951));
    Odrv4 I__441 (
            .O(N__3951),
            .I(\U712_CYCLE_TERM.N_362_i_0_en_0 ));
    IoInMux I__440 (
            .O(N__3948),
            .I(N__3945));
    LocalMux I__439 (
            .O(N__3945),
            .I(N__3942));
    Span12Mux_s10_v I__438 (
            .O(N__3942),
            .I(N__3939));
    Odrv12 I__437 (
            .O(N__3939),
            .I(VBENn_c));
    InMux I__436 (
            .O(N__3936),
            .I(N__3932));
    InMux I__435 (
            .O(N__3935),
            .I(N__3929));
    LocalMux I__434 (
            .O(N__3932),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__433 (
            .O(N__3929),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__432 (
            .O(N__3924),
            .I(N__3920));
    InMux I__431 (
            .O(N__3923),
            .I(N__3917));
    LocalMux I__430 (
            .O(N__3920),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__429 (
            .O(N__3917),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__428 (
            .O(N__3912),
            .I(N__3908));
    InMux I__427 (
            .O(N__3911),
            .I(N__3905));
    InMux I__426 (
            .O(N__3908),
            .I(N__3902));
    LocalMux I__425 (
            .O(N__3905),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__424 (
            .O(N__3902),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__423 (
            .O(N__3897),
            .I(N__3893));
    InMux I__422 (
            .O(N__3896),
            .I(N__3890));
    LocalMux I__421 (
            .O(N__3893),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__420 (
            .O(N__3890),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__419 (
            .O(N__3885),
            .I(N__3881));
    InMux I__418 (
            .O(N__3884),
            .I(N__3878));
    LocalMux I__417 (
            .O(N__3881),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__416 (
            .O(N__3878),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__415 (
            .O(N__3873),
            .I(N__3869));
    InMux I__414 (
            .O(N__3872),
            .I(N__3866));
    LocalMux I__413 (
            .O(N__3869),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__412 (
            .O(N__3866),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__411 (
            .O(N__3861),
            .I(N__3858));
    InMux I__410 (
            .O(N__3858),
            .I(N__3854));
    InMux I__409 (
            .O(N__3857),
            .I(N__3850));
    LocalMux I__408 (
            .O(N__3854),
            .I(N__3847));
    InMux I__407 (
            .O(N__3853),
            .I(N__3844));
    LocalMux I__406 (
            .O(N__3850),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv12 I__405 (
            .O(N__3847),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__404 (
            .O(N__3844),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__403 (
            .O(N__3837),
            .I(N__3834));
    LocalMux I__402 (
            .O(N__3834),
            .I(N__3831));
    IoSpan4Mux I__401 (
            .O(N__3831),
            .I(N__3828));
    Span4Mux_s3_h I__400 (
            .O(N__3828),
            .I(N__3825));
    Span4Mux_h I__399 (
            .O(N__3825),
            .I(N__3822));
    Sp12to4 I__398 (
            .O(N__3822),
            .I(N__3819));
    Span12Mux_v I__397 (
            .O(N__3819),
            .I(N__3815));
    InMux I__396 (
            .O(N__3818),
            .I(N__3812));
    Odrv12 I__395 (
            .O(N__3815),
            .I(TACK_OUTn));
    LocalMux I__394 (
            .O(N__3812),
            .I(TACK_OUTn));
    InMux I__393 (
            .O(N__3807),
            .I(N__3803));
    InMux I__392 (
            .O(N__3806),
            .I(N__3800));
    LocalMux I__391 (
            .O(N__3803),
            .I(N__3797));
    LocalMux I__390 (
            .O(N__3800),
            .I(N__3794));
    Odrv4 I__389 (
            .O(N__3797),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    Odrv4 I__388 (
            .O(N__3794),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__387 (
            .O(N__3789),
            .I(N__3786));
    LocalMux I__386 (
            .O(N__3786),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ));
    InMux I__385 (
            .O(N__3783),
            .I(N__3780));
    LocalMux I__384 (
            .O(N__3780),
            .I(N__3774));
    InMux I__383 (
            .O(N__3779),
            .I(N__3767));
    InMux I__382 (
            .O(N__3778),
            .I(N__3767));
    InMux I__381 (
            .O(N__3777),
            .I(N__3767));
    Span4Mux_h I__380 (
            .O(N__3774),
            .I(N__3762));
    LocalMux I__379 (
            .O(N__3767),
            .I(N__3762));
    Span4Mux_v I__378 (
            .O(N__3762),
            .I(N__3759));
    Span4Mux_h I__377 (
            .O(N__3759),
            .I(N__3756));
    Span4Mux_v I__376 (
            .O(N__3756),
            .I(N__3753));
    Span4Mux_v I__375 (
            .O(N__3753),
            .I(N__3750));
    Odrv4 I__374 (
            .O(N__3750),
            .I(CLK40_OUT_i));
    InMux I__373 (
            .O(N__3747),
            .I(N__3735));
    InMux I__372 (
            .O(N__3746),
            .I(N__3735));
    InMux I__371 (
            .O(N__3745),
            .I(N__3735));
    InMux I__370 (
            .O(N__3744),
            .I(N__3735));
    LocalMux I__369 (
            .O(N__3735),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__368 (
            .O(N__3732),
            .I(N__3729));
    LocalMux I__367 (
            .O(N__3729),
            .I(\U712_BYTE_ENABLE.N_455 ));
    InMux I__366 (
            .O(N__3726),
            .I(N__3720));
    InMux I__365 (
            .O(N__3725),
            .I(N__3720));
    LocalMux I__364 (
            .O(N__3720),
            .I(N__3717));
    Span4Mux_v I__363 (
            .O(N__3717),
            .I(N__3714));
    Sp12to4 I__362 (
            .O(N__3714),
            .I(N__3711));
    Span12Mux_h I__361 (
            .O(N__3711),
            .I(N__3708));
    Span12Mux_v I__360 (
            .O(N__3708),
            .I(N__3705));
    Odrv12 I__359 (
            .O(N__3705),
            .I(SIZ_c_1));
    CascadeMux I__358 (
            .O(N__3702),
            .I(\U712_BYTE_ENABLE.N_352_cascade_ ));
    IoInMux I__357 (
            .O(N__3699),
            .I(N__3696));
    LocalMux I__356 (
            .O(N__3696),
            .I(N__3693));
    IoSpan4Mux I__355 (
            .O(N__3693),
            .I(N__3690));
    Span4Mux_s3_v I__354 (
            .O(N__3690),
            .I(N__3687));
    Sp12to4 I__353 (
            .O(N__3687),
            .I(N__3684));
    Span12Mux_v I__352 (
            .O(N__3684),
            .I(N__3681));
    Span12Mux_h I__351 (
            .O(N__3681),
            .I(N__3678));
    Odrv12 I__350 (
            .O(N__3678),
            .I(N_49_i));
    IoInMux I__349 (
            .O(N__3675),
            .I(N__3672));
    LocalMux I__348 (
            .O(N__3672),
            .I(N__3669));
    Span12Mux_s5_h I__347 (
            .O(N__3669),
            .I(N__3666));
    Odrv12 I__346 (
            .O(N__3666),
            .I(CLK40_OUT_i_i));
    InMux I__345 (
            .O(N__3663),
            .I(N__3657));
    InMux I__344 (
            .O(N__3662),
            .I(N__3657));
    LocalMux I__343 (
            .O(N__3657),
            .I(N__3654));
    Sp12to4 I__342 (
            .O(N__3654),
            .I(N__3651));
    Span12Mux_v I__341 (
            .O(N__3651),
            .I(N__3648));
    Odrv12 I__340 (
            .O(N__3648),
            .I(A_c_1));
    InMux I__339 (
            .O(N__3645),
            .I(N__3642));
    LocalMux I__338 (
            .O(N__3642),
            .I(N__3639));
    Odrv4 I__337 (
            .O(N__3639),
            .I(\U712_BYTE_ENABLE.N_457 ));
    InMux I__336 (
            .O(N__3636),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__335 (
            .O(N__3633),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__334 (
            .O(N__3630),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__333 (
            .O(N__3627),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__332 (
            .O(N__3624),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__331 (
            .O(N__3621),
            .I(N__3618));
    GlobalMux I__330 (
            .O(N__3618),
            .I(N__3615));
    gio2CtrlBuf I__329 (
            .O(N__3615),
            .I(C1_c_g));
    InMux I__328 (
            .O(N__3612),
            .I(N__3609));
    LocalMux I__327 (
            .O(N__3609),
            .I(TACK_EN_i_ess));
    IoInMux I__326 (
            .O(N__3606),
            .I(N__3603));
    LocalMux I__325 (
            .O(N__3603),
            .I(N__3600));
    Span12Mux_s5_h I__324 (
            .O(N__3600),
            .I(N__3597));
    Span12Mux_v I__323 (
            .O(N__3597),
            .I(N__3594));
    Odrv12 I__322 (
            .O(N__3594),
            .I(N_888_i));
    CascadeMux I__321 (
            .O(N__3591),
            .I(\U712_BYTE_ENABLE.N_451_cascade_ ));
    IoInMux I__320 (
            .O(N__3588),
            .I(N__3585));
    LocalMux I__319 (
            .O(N__3585),
            .I(N__3582));
    Span4Mux_s2_h I__318 (
            .O(N__3582),
            .I(N__3579));
    Span4Mux_h I__317 (
            .O(N__3579),
            .I(N__3576));
    Sp12to4 I__316 (
            .O(N__3576),
            .I(N__3573));
    Span12Mux_v I__315 (
            .O(N__3573),
            .I(N__3570));
    Span12Mux_h I__314 (
            .O(N__3570),
            .I(N__3567));
    Odrv12 I__313 (
            .O(N__3567),
            .I(N_48_i));
    IoInMux I__312 (
            .O(N__3564),
            .I(N__3561));
    LocalMux I__311 (
            .O(N__3561),
            .I(N__3558));
    Span4Mux_s2_v I__310 (
            .O(N__3558),
            .I(N__3555));
    Span4Mux_v I__309 (
            .O(N__3555),
            .I(N__3552));
    Odrv4 I__308 (
            .O(N__3552),
            .I(CLK80_OUT_i_i));
    InMux I__307 (
            .O(N__3549),
            .I(bfn_7_7_0_));
    InMux I__306 (
            .O(N__3546),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__305 (
            .O(N__3543),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    IoInMux I__304 (
            .O(N__3540),
            .I(N__3537));
    LocalMux I__303 (
            .O(N__3537),
            .I(N__3534));
    Span4Mux_s0_v I__302 (
            .O(N__3534),
            .I(N__3531));
    Span4Mux_v I__301 (
            .O(N__3531),
            .I(N__3528));
    Sp12to4 I__300 (
            .O(N__3528),
            .I(N__3525));
    Span12Mux_h I__299 (
            .O(N__3525),
            .I(N__3522));
    Span12Mux_v I__298 (
            .O(N__3522),
            .I(N__3519));
    Odrv12 I__297 (
            .O(N__3519),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7437),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5888),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_3.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_3.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9162),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__3897),
            .in2(_gnd_net_),
            .in3(N__3549),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__3924),
            .in2(_gnd_net_),
            .in3(N__3546),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__3936),
            .in2(_gnd_net_),
            .in3(N__3543),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__5459),
            .in2(_gnd_net_),
            .in3(N__3636),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__3911),
            .in2(_gnd_net_),
            .in3(N__3633),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__3873),
            .in2(_gnd_net_),
            .in3(N__3630),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__3885),
            .in2(_gnd_net_),
            .in3(N__3627),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__5429),
            .in2(_gnd_net_),
            .in3(N__3624),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3621),
            .ce(),
            .sr(N__4953));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_8_3 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_8_3  (
            .in0(N__3978),
            .in1(N__7520),
            .in2(_gnd_net_),
            .in3(N__4016),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9157),
            .ce(N__3957),
            .sr(N__8965));
    defparam TACKn_obuft_RNO_LC_7_9_1.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_7_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_7_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3612),
            .lcout(N_888_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_9_4 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_9_4  (
            .in0(N__7374),
            .in1(N__3726),
            .in2(_gnd_net_),
            .in3(N__8155),
            .lcout(\U712_BYTE_ENABLE.N_451 ),
            .ltout(\U712_BYTE_ENABLE.N_451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_9_5 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \U712_BYTE_ENABLE.N_48_i_LC_7_9_5  (
            .in0(N__3645),
            .in1(N__6892),
            .in2(N__3591),
            .in3(N__4049),
            .lcout(N_48_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_o2_LC_7_9_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_o2_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_o2_LC_7_9_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_o2_LC_7_9_6  (
            .in0(N__6893),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3725),
            .lcout(\U712_BYTE_ENABLE.N_352 ),
            .ltout(\U712_BYTE_ENABLE.N_352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_49_i_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_7_9_7 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U712_BYTE_ENABLE.N_49_i_LC_7_9_7  (
            .in0(N__3732),
            .in1(N__7058),
            .in2(N__3702),
            .in3(N__7039),
            .lcout(N_49_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_7_10_1.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_7_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLK40C_obuf_RNO_LC_7_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3783),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_7_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_7_10_2  (
            .in0(N__3662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8156),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_1_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_1_LC_7_10_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_1_LC_7_10_4  (
            .in0(N__3663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8157),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(N__8972));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3857),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9145),
            .ce(),
            .sr(N__8972));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__3853),
            .in2(_gnd_net_),
            .in3(N__3806),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_8_7_3 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_8_7_3  (
            .in0(N__6111),
            .in1(_gnd_net_),
            .in2(N__4893),
            .in3(N__4730),
            .lcout(\U712_BYTE_ENABLE.N_453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_0_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_0_LC_8_7_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_0_LC_8_7_4  (
            .in0(N__4729),
            .in1(N__4888),
            .in2(_gnd_net_),
            .in3(N__6110),
            .lcout(\U712_BYTE_ENABLE.N_457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_7_6 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_7_6  (
            .in0(N__3935),
            .in1(N__3923),
            .in2(N__3912),
            .in3(N__3896),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_7_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__3884),
            .in2(_gnd_net_),
            .in3(N__3872),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_0 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_0  (
            .in0(N__3746),
            .in1(N__3818),
            .in2(N__3861),
            .in3(N__3777),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(N__8951));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_1  (
            .in0(N__3779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3745),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(N__8951));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_3 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_3  (
            .in0(N__3789),
            .in1(N__4015),
            .in2(N__3999),
            .in3(N__3744),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(N__8951));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_4 .LUT_INIT=16'b1010111110001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_4  (
            .in0(N__3747),
            .in1(N__3778),
            .in2(N__4017),
            .in3(N__3977),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9153),
            .ce(),
            .sr(N__8951));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_8_9_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_8_9_0  (
            .in0(N__4728),
            .in1(_gnd_net_),
            .in2(N__4848),
            .in3(N__6109),
            .lcout(\U712_BYTE_ENABLE.N_455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_8_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_8_9_1  (
            .in0(N__6108),
            .in1(N__4844),
            .in2(_gnd_net_),
            .in3(N__4727),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_47_i_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_8_9_2 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_BYTE_ENABLE.N_47_i_LC_8_9_2  (
            .in0(N__7046),
            .in1(N__4050),
            .in2(N__4038),
            .in3(N__4035),
            .lcout(N_47_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__4187),
            .in2(_gnd_net_),
            .in3(N__4308),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_6 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_9_6  (
            .in0(N__7503),
            .in1(N__3995),
            .in2(N__3981),
            .in3(N__3976),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_362_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_9_7  (
            .in0(N__9019),
            .in1(_gnd_net_),
            .in2(N__3960),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_362_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_5_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_5_3  (
            .in0(N__5400),
            .in1(N__7523),
            .in2(N__4563),
            .in3(N__4507),
            .lcout(\U712_CHIP_RAM.N_492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_9_5_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__4212),
            .in2(_gnd_net_),
            .in3(N__8118),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_6  (
            .in0(N__4532),
            .in1(N__5609),
            .in2(N__7527),
            .in3(N__5700),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_a3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_2 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_2  (
            .in0(N__5798),
            .in1(N__9026),
            .in2(N__4359),
            .in3(N__5827),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9136),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_3  (
            .in0(N__7743),
            .in1(N__8115),
            .in2(N__8817),
            .in3(N__8241),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_4  (
            .in0(N__8116),
            .in1(N__4170),
            .in2(N__4152),
            .in3(N__4149),
            .lcout(\U712_CHIP_RAM.N_374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__5797),
            .in2(_gnd_net_),
            .in3(N__4354),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_ac0_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_0  (
            .in0(N__4131),
            .in1(N__9022),
            .in2(N__4377),
            .in3(N__5829),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9146),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_7_3  (
            .in0(N__5828),
            .in1(N__4130),
            .in2(_gnd_net_),
            .in3(N__4373),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_4 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__9023),
            .in2(N__4122),
            .in3(N__4391),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9146),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_6 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_6  (
            .in0(N__4119),
            .in1(N__9024),
            .in2(N__4335),
            .in3(N__4392),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9146),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_7_7 .LUT_INIT=16'b0000000001000001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_7_7  (
            .in0(N__4531),
            .in1(N__5711),
            .in2(N__5613),
            .in3(N__4421),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_8_5  (
            .in0(N__4113),
            .in1(N__4559),
            .in2(_gnd_net_),
            .in3(N__5186),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9149),
            .ce(),
            .sr(N__8943));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_8_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_8_7  (
            .in0(N__4673),
            .in1(N__4090),
            .in2(_gnd_net_),
            .in3(N__4686),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9149),
            .ce(),
            .sr(N__8943));
    defparam \U712_BUFFERS.DRDDIR_i_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_0_LC_9_9_0 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_0_LC_9_9_0  (
            .in0(N__4207),
            .in1(N__7413),
            .in2(N__6097),
            .in3(N__4091),
            .lcout(DRDDIR_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_9_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__4208),
            .in2(_gnd_net_),
            .in3(N__6090),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_9_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_9_5  (
            .in0(N__4934),
            .in1(N__7114),
            .in2(_gnd_net_),
            .in3(N__7149),
            .lcout(\U712_REG_SM.N_343 ),
            .ltout(\U712_REG_SM.N_343_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_9_6 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__5916),
            .in2(N__4218),
            .in3(N__5952),
            .lcout(\U712_REG_SM.N_358 ),
            .ltout(\U712_REG_SM.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_9_7 .LUT_INIT=16'b1011101110001010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_9_7  (
            .in0(N__4787),
            .in1(N__6966),
            .in2(N__4215),
            .in3(N__4206),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9154),
            .ce(),
            .sr(N__8936));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_9_10_0  (
            .in0(N__6476),
            .in1(N__4786),
            .in2(N__6458),
            .in3(N__4800),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9158),
            .ce(),
            .sr(N__8931));
    defparam \U712_REG_SM.REG_TACK_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_9_10_7 .LUT_INIT=16'b1111101101010000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_9_10_7  (
            .in0(N__6965),
            .in1(N__6454),
            .in2(N__4191),
            .in3(N__6475),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9158),
            .ce(),
            .sr(N__8931));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM76F1_1_LC_10_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM76F1_1_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM76F1_1_LC_10_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIM76F1_1_LC_10_4_1  (
            .in0(_gnd_net_),
            .in1(N__5273),
            .in2(_gnd_net_),
            .in3(N__5608),
            .lcout(\U712_CHIP_RAM.N_563 ),
            .ltout(\U712_CHIP_RAM.N_563_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_4_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_4_2  (
            .in0(N__7518),
            .in1(N__4640),
            .in2(N__4176),
            .in3(N__4287),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_4_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(N__5243),
            .in2(N__4173),
            .in3(N__8650),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_4_4 .LUT_INIT=16'b0000100000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_4_4  (
            .in0(N__5607),
            .in1(N__4509),
            .in2(N__4422),
            .in3(N__5699),
            .lcout(\U712_CHIP_RAM.N_565 ),
            .ltout(\U712_CHIP_RAM.N_565_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_10_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_10_4_5 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_10_4_5  (
            .in0(N__5181),
            .in1(N__7519),
            .in2(N__4281),
            .in3(N__4257),
            .lcout(\U712_CHIP_RAM.N_445 ),
            .ltout(\U712_CHIP_RAM.N_445_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .LUT_INIT=16'b1010101100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6  (
            .in0(N__5244),
            .in1(N__4278),
            .in2(N__4272),
            .in3(N__7846),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9123),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_5_0 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_5_0  (
            .in0(N__4533),
            .in1(N__4256),
            .in2(_gnd_net_),
            .in3(N__5178),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_1 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_1  (
            .in0(N__7522),
            .in1(N__4269),
            .in2(N__4263),
            .in3(N__4419),
            .lcout(\U712_CHIP_RAM.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_5_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_10_5_2  (
            .in0(N__5778),
            .in1(N__5501),
            .in2(_gnd_net_),
            .in3(N__5119),
            .lcout(\U712_CHIP_RAM.N_333 ),
            .ltout(\U712_CHIP_RAM.N_333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_5_3 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_5_3  (
            .in0(N__5669),
            .in1(_gnd_net_),
            .in2(N__4260),
            .in3(N__5573),
            .lcout(\U712_CHIP_RAM.N_346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_10_5_4 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_10_5_4  (
            .in0(N__4581),
            .in1(N__5502),
            .in2(N__5796),
            .in3(N__4508),
            .lcout(\U712_CHIP_RAM.N_564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_5  (
            .in0(N__5503),
            .in1(N__5218),
            .in2(N__5802),
            .in3(N__4582),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_6 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_6  (
            .in0(N__5219),
            .in1(_gnd_net_),
            .in2(N__4452),
            .in3(N__5179),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_7 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_10_5_7  (
            .in0(N__4436),
            .in1(N__4641),
            .in2(N__4449),
            .in3(N__5707),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9127),
            .ce(),
            .sr(N__8966));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_6_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_6_0  (
            .in0(N__8117),
            .in1(N__4632),
            .in2(N__5520),
            .in3(N__4583),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_6_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_6_1  (
            .in0(N__4633),
            .in1(N__5672),
            .in2(N__4425),
            .in3(N__4420),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_6_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_6_2  (
            .in0(N__4390),
            .in1(N__4372),
            .in2(N__4358),
            .in3(N__4331),
            .lcout(\U712_CHIP_RAM.N_330 ),
            .ltout(\U712_CHIP_RAM.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_10_6_3 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__5574),
            .in2(N__4320),
            .in3(N__5670),
            .lcout(\U712_CHIP_RAM.N_493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_10_6_4 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_10_6_4  (
            .in0(N__5130),
            .in1(N__4593),
            .in2(N__4317),
            .in3(N__4304),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9132),
            .ce(),
            .sr(N__8952));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU9AV6_0_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU9AV6_0_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU9AV6_0_LC_10_6_5 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIU9AV6_0_LC_10_6_5  (
            .in0(N__4766),
            .in1(N__5255),
            .in2(N__5133),
            .in3(N__5671),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_6_6 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_6_6  (
            .in0(N__9025),
            .in1(N__4467),
            .in2(N__4290),
            .in3(N__5180),
            .lcout(\U712_CHIP_RAM.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_0  (
            .in0(N__5784),
            .in1(N__5710),
            .in2(N__5603),
            .in3(N__5217),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_7_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_7_1  (
            .in0(N__4494),
            .in1(N__5393),
            .in2(_gnd_net_),
            .in3(N__4554),
            .lcout(\U712_CHIP_RAM.N_332 ),
            .ltout(\U712_CHIP_RAM.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_10_7_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_10_7_2  (
            .in0(N__5783),
            .in1(N__5576),
            .in2(N__4587),
            .in3(N__5510),
            .lcout(\U712_CHIP_RAM.N_560 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_3 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_3  (
            .in0(N__4497),
            .in1(N__4584),
            .in2(N__5519),
            .in3(N__5785),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9137),
            .ce(),
            .sr(N__8944));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_4 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_4  (
            .in0(N__5392),
            .in1(N__4555),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(\U712_CHIP_RAM.N_351 ),
            .ltout(\U712_CHIP_RAM.N_351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_2_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_2_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_2_LC_10_7_5 .LUT_INIT=16'b0010011000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_2_LC_10_7_5  (
            .in0(N__5509),
            .in1(N__5586),
            .in2(N__4512),
            .in3(N__4473),
            .lcout(\U712_CHIP_RAM.N_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP0891_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP0891_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP0891_LC_10_7_6 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP0891_LC_10_7_6  (
            .in0(N__5782),
            .in1(N__5575),
            .in2(_gnd_net_),
            .in3(N__4495),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__5207),
            .in2(_gnd_net_),
            .in3(N__4458),
            .lcout(\U712_CHIP_RAM.N_402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_1  (
            .in0(N__5300),
            .in1(N__5937),
            .in2(N__6050),
            .in3(N__5902),
            .lcout(\U712_CHIP_RAM.N_341 ),
            .ltout(\U712_CHIP_RAM.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI7Q5U5_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__5208),
            .in2(N__4770),
            .in3(N__5185),
            .lcout(\U712_CHIP_RAM.N_450 ),
            .ltout(\U712_CHIP_RAM.N_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_10_8_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_10_8_3  (
            .in0(N__4767),
            .in1(N__5708),
            .in2(N__4755),
            .in3(N__5132),
            .lcout(\U712_CHIP_RAM.N_326 ),
            .ltout(\U712_CHIP_RAM.N_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_4 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_4  (
            .in0(N__5709),
            .in1(N__8076),
            .in2(N__4752),
            .in3(N__6037),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9147),
            .ce(),
            .sr(N__8937));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_10_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_10_8_5  (
            .in0(N__4749),
            .in1(N__6084),
            .in2(_gnd_net_),
            .in3(N__4604),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9147),
            .ce(),
            .sr(N__8937));
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_6 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_8_6  (
            .in0(N__7752),
            .in1(N__4704),
            .in2(N__4605),
            .in3(N__4748),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9147),
            .ce(),
            .sr(N__8937));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_8_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_8_7  (
            .in0(N__9018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4685),
            .lcout(\U712_CHIP_RAM.N_450_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_9_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_9_0  (
            .in0(N__4674),
            .in1(N__5307),
            .in2(N__7424),
            .in3(N__6053),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9150),
            .ce(N__4614),
            .sr(N__8932));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_10_9_1  (
            .in0(N__6052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5715),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_9_3  (
            .in0(N__7146),
            .in1(N__4935),
            .in2(_gnd_net_),
            .in3(N__7115),
            .lcout(\U712_REG_SM.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_9_4  (
            .in0(N__6435),
            .in1(N__6766),
            .in2(N__6402),
            .in3(N__6722),
            .lcout(\U712_REG_SM.N_338 ),
            .ltout(\U712_REG_SM.N_338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_9_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_10_9_5  (
            .in0(N__7147),
            .in1(N__5989),
            .in2(N__4923),
            .in3(N__7116),
            .lcout(\U712_REG_SM.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_10_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__6767),
            .in2(_gnd_net_),
            .in3(N__6721),
            .lcout(\U712_REG_SM.N_354 ),
            .ltout(\U712_REG_SM.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_10_9_7 .LUT_INIT=16'b0101010100000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_10_9_7  (
            .in0(N__6808),
            .in1(N__6983),
            .in2(N__4920),
            .in3(N__6270),
            .lcout(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_10_1 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_10_10_1  (
            .in0(N__5375),
            .in1(N__6260),
            .in2(N__4917),
            .in3(N__6225),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8928));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_10_10_2  (
            .in0(N__4892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4838),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8928));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6149),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8928));
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_REG_SM.DS_EN_LC_10_10_4  (
            .in0(N__7559),
            .in1(N__4806),
            .in2(N__5079),
            .in3(N__6132),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8928));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_10_6 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_10_10_6  (
            .in0(N__4788),
            .in1(N__6009),
            .in2(N__5997),
            .in3(N__4799),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9155),
            .ce(),
            .sr(N__8928));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_11_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_10_11_0  (
            .in0(N__7420),
            .in1(N__6391),
            .in2(_gnd_net_),
            .in3(N__6733),
            .lcout(\U712_REG_SM.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_2_0  (
            .in0(N__5001),
            .in1(N__8577),
            .in2(_gnd_net_),
            .in3(N__8654),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9116),
            .ce(N__8475),
            .sr(N__8978));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_3_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_3_2 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_3_2  (
            .in0(N__8539),
            .in1(N__8788),
            .in2(_gnd_net_),
            .in3(N__8614),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_7 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_7  (
            .in0(N__5043),
            .in1(N__6279),
            .in2(N__5025),
            .in3(N__8153),
            .lcout(\U712_CHIP_RAM.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_4_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_4_1  (
            .in0(N__8538),
            .in1(N__5242),
            .in2(_gnd_net_),
            .in3(N__4995),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_3  (
            .in0(N__8161),
            .in1(N__4989),
            .in2(N__5739),
            .in3(N__4971),
            .lcout(\U712_CHIP_RAM.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_4_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_4_6  (
            .in0(N__8536),
            .in1(N__8613),
            .in2(N__8769),
            .in3(N__7838),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_4_7 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_4_7  (
            .in0(N__8537),
            .in1(N__8733),
            .in2(N__4938),
            .in3(N__7839),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_11_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_11_5_0  (
            .in0(N__5123),
            .in1(N__5791),
            .in2(N__5838),
            .in3(N__5139),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICDSCD_0_LC_11_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICDSCD_0_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICDSCD_0_LC_11_5_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNICDSCD_0_LC_11_5_1  (
            .in0(N__5091),
            .in1(N__5277),
            .in2(N__5262),
            .in3(N__5259),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_5_2 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__5229),
            .in2(N__5223),
            .in3(N__8768),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_5_3 .LUT_INIT=16'b1111000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_5_3  (
            .in0(N__5220),
            .in1(N__5085),
            .in2(N__5187),
            .in3(N__5679),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_5_4 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_5_4  (
            .in0(N__9021),
            .in1(_gnd_net_),
            .in2(N__5142),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9124),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_5_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_5_5  (
            .in0(N__5590),
            .in1(N__5677),
            .in2(_gnd_net_),
            .in3(N__5514),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_11_5_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_11_5_6  (
            .in0(N__5678),
            .in1(_gnd_net_),
            .in2(N__5131),
            .in3(N__7521),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_6_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_6_0  (
            .in0(N__5912),
            .in1(N__5948),
            .in2(N__6051),
            .in3(N__5302),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_0_i_a3_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7TES1_LC_11_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7TES1_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7TES1_LC_11_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI7TES1_LC_11_6_1  (
            .in0(N__5578),
            .in1(N__5674),
            .in2(N__5518),
            .in3(N__6038),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRB433_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRB433_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIRB433_LC_11_6_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIRB433_LC_11_6_2  (
            .in0(N__5911),
            .in1(N__5947),
            .in2(N__5841),
            .in3(N__5301),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_11_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_11_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_11_6_3  (
            .in0(N__5577),
            .in1(N__5673),
            .in2(_gnd_net_),
            .in3(N__5504),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_4 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__5795),
            .in2(N__5805),
            .in3(N__5727),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_6_5 .LUT_INIT=16'b0000111100110101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_6_5  (
            .in0(N__6573),
            .in1(N__6660),
            .in2(N__8789),
            .in3(N__8104),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_6_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_6_6  (
            .in0(N__5675),
            .in1(N__5582),
            .in2(_gnd_net_),
            .in3(N__5725),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_6_7  (
            .in0(N__5726),
            .in1(N__5676),
            .in2(N__5599),
            .in3(N__5505),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9128),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_7_0 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_7_0  (
            .in0(N__5460),
            .in1(N__5445),
            .in2(N__5436),
            .in3(N__5415),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9133),
            .ce(),
            .sr(N__8938));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_11_7_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_11_7_1  (
            .in0(N__8074),
            .in1(N__5406),
            .in2(_gnd_net_),
            .in3(N__6086),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9133),
            .ce(),
            .sr(N__8938));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_7_4 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_7_4  (
            .in0(N__5379),
            .in1(N__8075),
            .in2(N__5343),
            .in3(N__5306),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9133),
            .ce(),
            .sr(N__8938));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_7_6  (
            .in0(N__6168),
            .in1(N__6153),
            .in2(N__6054),
            .in3(N__6085),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9133),
            .ce(),
            .sr(N__8938));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_8_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_11_8_0  (
            .in0(N__5993),
            .in1(N__6861),
            .in2(_gnd_net_),
            .in3(N__6008),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9138),
            .ce(),
            .sr(N__8933));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_11_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5973),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9138),
            .ce(),
            .sr(N__8933));
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6732),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9138),
            .ce(),
            .sr(N__8933));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_11_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_11_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5946),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9138),
            .ce(),
            .sr(N__8933));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5889),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9138),
            .ce(),
            .sr(N__8933));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_9_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_11_9_0  (
            .in0(N__6860),
            .in1(N__5853),
            .in2(N__6240),
            .in3(N__6259),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8929));
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_11_9_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_11_9_1  (
            .in0(N__7142),
            .in1(N__5852),
            .in2(_gnd_net_),
            .in3(N__7100),
            .lcout(\U712_REG_SM.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6398),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8929));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_11_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__7099),
            .in2(_gnd_net_),
            .in3(N__7141),
            .lcout(\U712_REG_SM.N_347 ),
            .ltout(\U712_REG_SM.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_11_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_11_9_5  (
            .in0(N__6925),
            .in1(N__6768),
            .in2(N__6273),
            .in3(N__6720),
            .lcout(\U712_REG_SM.N_559 ),
            .ltout(\U712_REG_SM.N_559_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_9_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_9_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_9_6  (
            .in0(N__6235),
            .in1(N__6258),
            .in2(N__6264),
            .in3(N__6809),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8929));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_11_9_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_11_9_7  (
            .in0(N__6224),
            .in1(N__6261),
            .in2(N__6870),
            .in3(N__6236),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9148),
            .ce(),
            .sr(N__8929));
    defparam \U712_REG_SM.REGENn_1_ess_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_LC_11_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_ess_LC_11_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_LC_11_10_0  (
            .in0(N__6779),
            .in1(N__6926),
            .in2(N__6743),
            .in3(N__6691),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9151),
            .ce(N__6120),
            .sr(N__8923));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_10_1 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_10_1  (
            .in0(N__9016),
            .in1(N__6164),
            .in2(_gnd_net_),
            .in3(N__6148),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_11_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_RNO_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__9017),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(\U712_REG_SM.N_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_11_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__6387),
            .in2(_gnd_net_),
            .in3(N__6428),
            .lcout(\U712_REG_SM.N_348 ),
            .ltout(\U712_REG_SM.N_348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_11_11_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__7001),
            .in2(N__6114),
            .in3(N__6692),
            .lcout(\U712_REG_SM.N_364 ),
            .ltout(\U712_REG_SM.N_364_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_11_4 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_11_4  (
            .in0(N__6483),
            .in1(N__6952),
            .in2(N__6462),
            .in3(N__6459),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9156),
            .ce(),
            .sr(N__8922));
    defparam \U712_REG_SM.C1_SYNC_2_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_11_11_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_11_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_11_11_5  (
            .in0(N__6780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9156),
            .ce(),
            .sr(N__8922));
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_11_11_6  (
            .in0(N__6417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9156),
            .ce(),
            .sr(N__8922));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_3_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_3_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_3_2  (
            .in0(N__8676),
            .in1(N__6366),
            .in2(_gnd_net_),
            .in3(N__8559),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9115),
            .ce(N__8464),
            .sr(N__8964));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3  (
            .in0(N__8558),
            .in1(N__8677),
            .in2(N__8813),
            .in3(N__6285),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9115),
            .ce(N__8464),
            .sr(N__8964));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_3 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_3  (
            .in0(N__8159),
            .in1(N__6648),
            .in2(N__6495),
            .in3(N__8758),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_4  (
            .in0(N__6327),
            .in1(N__6306),
            .in2(N__6288),
            .in3(N__8160),
            .lcout(\U712_CHIP_RAM.N_368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_6 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_6  (
            .in0(N__6540),
            .in1(N__8158),
            .in2(N__8790),
            .in3(N__6654),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_4_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_4_7  (
            .in0(N__6666),
            .in1(N__9020),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_5_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__6567),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9119),
            .ce(N__8193),
            .sr(N__8942));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6527),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9119),
            .ce(N__8193),
            .sr(N__8942));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7983),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9119),
            .ce(N__8193),
            .sr(N__8942));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_12_6_2  (
            .in0(N__9221),
            .in1(N__7281),
            .in2(N__6642),
            .in3(N__8154),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8467),
            .sr(N__8935));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_12_6_7  (
            .in0(N__6603),
            .in1(N__8576),
            .in2(_gnd_net_),
            .in3(N__8671),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9122),
            .ce(N__8467),
            .sr(N__8935));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_1  (
            .in0(N__8423),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9126),
            .ce(N__7923),
            .sr(N__8930));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6566),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9126),
            .ce(N__7923),
            .sr(N__8930));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_7_6  (
            .in0(N__6531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9126),
            .ce(N__7923),
            .sr(N__8930));
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_12_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7148),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9131),
            .ce(),
            .sr(N__8927));
    defparam \U712_BYTE_ENABLE.N_50_i_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_50_i_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_50_i_LC_12_9_5 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \U712_BYTE_ENABLE.N_50_i_LC_12_9_5  (
            .in0(N__6909),
            .in1(N__7083),
            .in2(N__7071),
            .in3(N__7047),
            .lcout(N_50_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_12_9_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_12_9_7  (
            .in0(N__7002),
            .in1(N__6984),
            .in2(_gnd_net_),
            .in3(N__6810),
            .lcout(\U712_REG_SM.N_395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_10_3 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_12_10_3  (
            .in0(N__6672),
            .in1(N__6972),
            .in2(N__6930),
            .in3(N__6951),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9141),
            .ce(),
            .sr(N__8921));
    defparam \U712_REG_SM.LDS_OUT_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_12_10_5 .LUT_INIT=16'b1100110010101111;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_12_10_5  (
            .in0(N__6907),
            .in1(N__6836),
            .in2(N__7340),
            .in3(N__6862),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9141),
            .ce(),
            .sr(N__8921));
    defparam \U712_REG_SM.UDS_OUT_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_12_10_7 .LUT_INIT=16'b1100110001011111;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_12_10_7  (
            .in0(N__6908),
            .in1(N__7583),
            .in2(N__7341),
            .in3(N__6863),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9141),
            .ce(),
            .sr(N__8921));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_12_11_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_12_11_2  (
            .in0(N__6837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7571),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_12_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_12_11_3  (
            .in0(N__6807),
            .in1(N__6778),
            .in2(N__6744),
            .in3(N__6693),
            .lcout(\U712_REG_SM.N_433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_12_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_12_0  (
            .in0(N__7587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7572),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_12_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_12_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7473),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_2_0_a3_0_a3_0_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_2_0_a3_0_a3_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_2_0_a3_0_a3_0_LC_12_12_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U712_REG_SM.LDS_OUT_2_0_a3_0_a3_0_LC_12_12_3  (
            .in0(N__7425),
            .in1(N__7373),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_a3_0_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_3_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_3_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_3_2  (
            .in0(N__8578),
            .in1(N__8679),
            .in2(N__8820),
            .in3(N__7853),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9117),
            .ce(N__8466),
            .sr(N__8973));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_3_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_3_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_3_5  (
            .in0(N__8678),
            .in1(N__7653),
            .in2(_gnd_net_),
            .in3(N__8579),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9117),
            .ce(N__8466),
            .sr(N__8973));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_3_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_3_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_3_7 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_3_7  (
            .in0(N__7280),
            .in1(N__7263),
            .in2(N__8358),
            .in3(N__8162),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9117),
            .ce(N__8466),
            .sr(N__8973));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_1 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_1  (
            .in0(N__7224),
            .in1(N__7155),
            .in2(N__7203),
            .in3(N__8144),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_5_2 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(N__8580),
            .in2(N__7176),
            .in3(N__8672),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9125),
            .ce(N__8465),
            .sr(N__8953));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_6_6 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_6_6  (
            .in0(N__7950),
            .in1(N__8142),
            .in2(N__8818),
            .in3(N__8202),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_8_0  (
            .in0(N__8231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9139),
            .ce(N__7924),
            .sr(N__8934));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_8_5  (
            .in0(N__8381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9139),
            .ce(N__7924),
            .sr(N__8934));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_4_2 .LUT_INIT=16'b1110001100100011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_4_2  (
            .in0(N__7731),
            .in1(N__7611),
            .in2(N__8163),
            .in3(N__7716),
            .lcout(\U712_CHIP_RAM.N_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_4_5 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_4_5  (
            .in0(N__7695),
            .in1(N__8152),
            .in2(N__7677),
            .in3(N__7599),
            .lcout(\U712_CHIP_RAM.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_4_7 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_4_7  (
            .in0(N__7647),
            .in1(N__8151),
            .in2(N__7629),
            .in3(N__7989),
            .lcout(\U712_CHIP_RAM.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_5_1 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_5_1  (
            .in0(N__8130),
            .in1(N__7605),
            .in2(N__8800),
            .in3(N__8310),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_5_2  (
            .in0(N__8304),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9129),
            .ce(N__7935),
            .sr(N__8967));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_5_3 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_5_3  (
            .in0(N__8391),
            .in1(N__7593),
            .in2(N__8802),
            .in3(N__8143),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8339),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9129),
            .ce(N__7935),
            .sr(N__8967));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_5_5 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_14_5_5  (
            .in0(N__8131),
            .in1(N__7944),
            .in2(N__8801),
            .in3(N__8280),
            .lcout(\U712_CHIP_RAM.CMA_5_3_i_m2_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7976),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9134),
            .ce(N__7931),
            .sr(N__8954));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_14_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_14_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_14_6_4  (
            .in0(N__8274),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9134),
            .ce(N__7931),
            .sr(N__8954));
    defparam \U712_CHIP_RAM.CASn_LC_15_1_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_15_1_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_15_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8812),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(),
            .sr(N__8982));
    defparam \U712_CHIP_RAM.WEn_LC_15_1_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_15_1_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_15_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_15_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8673),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9118),
            .ce(),
            .sr(N__8982));
    defparam \U712_CHIP_RAM.CRCSn_LC_15_2_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_2_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_15_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7857),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9121),
            .ce(),
            .sr(N__8981));
    defparam \U712_CHIP_RAM.RASn_LC_15_2_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_15_2_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_15_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8583),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9121),
            .ce(),
            .sr(N__8981));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_4_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_15_4_2  (
            .in0(N__7779),
            .in1(_gnd_net_),
            .in2(N__8675),
            .in3(N__8581),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9130),
            .ce(N__8474),
            .sr(N__8979));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_15_4_6 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_15_4_6  (
            .in0(N__8826),
            .in1(N__8819),
            .in2(N__8674),
            .in3(N__8582),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9130),
            .ce(N__8474),
            .sr(N__8979));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_5_1  (
            .in0(N__8424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(N__8186),
            .sr(N__8974));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8385),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(N__8186),
            .sr(N__8974));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8343),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(N__8186),
            .sr(N__8974));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8303),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9135),
            .ce(N__8186),
            .sr(N__8974));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8270),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9140),
            .ce(N__8185),
            .sr(N__8968));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_6_4  (
            .in0(N__8232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9140),
            .ce(N__8185),
            .sr(N__8968));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_6_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_6_3  (
            .in0(N__9027),
            .in1(N__8169),
            .in2(_gnd_net_),
            .in3(N__9173),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_6_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9174),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9152),
            .ce(),
            .sr(N__8980));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_6_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_17_6_6  (
            .in0(N__9222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9189),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9152),
            .ce(),
            .sr(N__8980));
endmodule // U712_TOP

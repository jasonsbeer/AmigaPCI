-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 6 2024 09:04:20

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    CLK40B : out std_logic;
    TAn : out std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TBIn : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : in std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__7741\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \RnW_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \U111_CYCLE_SM.TS_EN10_cascade_\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_r_1\ : std_logic;
signal \INVU111_CYCLE_SM.A_OUTC_net\ : std_logic;
signal \CLK40\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_4\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \TAn_0_i\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \INVU111_CYCLE_SM.TA_EN_nessC_net\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\ : std_logic;
signal \TACKn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANS_0\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \U111_CYCLE_SM.FLIP\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \TACKn_wire\ <= TACKn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    CLK40A <= \CLK40A_wire\;
    TBIn <= \TBIn_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    TAn <= \TAn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__2876\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__7741\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__7741\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7725\,
            DIN => \N__7724\,
            DOUT => \N__7723\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7725\,
            PADOUT => \N__7724\,
            PADIN => \N__7723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4892\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__5651\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7716\,
            DIN => \N__7715\,
            DOUT => \N__7714\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7716\,
            PADOUT => \N__7715\,
            PADIN => \N__7714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2463\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__5984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7707\,
            DIN => \N__7706\,
            DOUT => \N__7705\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7707\,
            PADOUT => \N__7706\,
            PADIN => \N__7705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2471\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__5501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7698\,
            DIN => \N__7697\,
            DOUT => \N__7696\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7698\,
            PADOUT => \N__7697\,
            PADIN => \N__7696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TACKn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7689\,
            DIN => \N__7688\,
            DOUT => \N__7687\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7689\,
            PADOUT => \N__7688\,
            PADIN => \N__7687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4951\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__4103\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7680\,
            DIN => \N__7679\,
            DOUT => \N__7678\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7680\,
            PADOUT => \N__7679\,
            PADIN => \N__7678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7671\,
            DIN => \N__7670\,
            DOUT => \N__7669\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7671\,
            PADOUT => \N__7670\,
            PADIN => \N__7669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4995\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__2897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7662\,
            DIN => \N__7661\,
            DOUT => \N__7660\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7662\,
            PADOUT => \N__7661\,
            PADIN => \N__7660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2462\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__3290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7653\,
            DIN => \N__7652\,
            DOUT => \N__7651\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7653\,
            PADOUT => \N__7652\,
            PADIN => \N__7651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2450\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__3329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7644\,
            DIN => \N__7643\,
            DOUT => \N__7642\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7644\,
            PADOUT => \N__7643\,
            PADIN => \N__7642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4946\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__6437\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7635\,
            DIN => \N__7634\,
            DOUT => \N__7633\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7635\,
            PADOUT => \N__7634\,
            PADIN => \N__7633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7626\,
            DIN => \N__7625\,
            DOUT => \N__7624\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7626\,
            PADOUT => \N__7625\,
            PADIN => \N__7624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2310\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__6071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7617\,
            DIN => \N__7616\,
            DOUT => \N__7615\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7617\,
            PADOUT => \N__7616\,
            PADIN => \N__7615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4996\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__3143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7608\,
            DIN => \N__7607\,
            DOUT => \N__7606\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7608\,
            PADOUT => \N__7607\,
            PADIN => \N__7606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2470\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3065\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7599\,
            DIN => \N__7598\,
            DOUT => \N__7597\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7599\,
            PADOUT => \N__7598\,
            PADIN => \N__7597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2362\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__2963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7590\,
            DIN => \N__7589\,
            DOUT => \N__7588\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7590\,
            PADOUT => \N__7589\,
            PADIN => \N__7588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7581\,
            DIN => \N__7580\,
            DOUT => \N__7579\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7581\,
            PADOUT => \N__7580\,
            PADIN => \N__7579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4807\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__3809\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7572\,
            DIN => \N__7571\,
            DOUT => \N__7570\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7572\,
            PADOUT => \N__7571\,
            PADIN => \N__7570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4947\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__4163\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7563\,
            DIN => \N__7562\,
            DOUT => \N__7561\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7563\,
            PADOUT => \N__7562\,
            PADIN => \N__7561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3471\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7554\,
            DIN => \N__7553\,
            DOUT => \N__7552\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7554\,
            PADOUT => \N__7553\,
            PADIN => \N__7552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2363\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__3593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7545\,
            DIN => \N__7544\,
            DOUT => \N__7543\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7545\,
            PADOUT => \N__7544\,
            PADIN => \N__7543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4869\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6236\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7536\,
            DIN => \N__7535\,
            DOUT => \N__7534\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7536\,
            PADOUT => \N__7535\,
            PADIN => \N__7534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2407\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__2774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7527\,
            DIN => \N__7526\,
            DOUT => \N__7525\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7527\,
            PADOUT => \N__7526\,
            PADIN => \N__7525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7518\,
            DIN => \N__7517\,
            DOUT => \N__7516\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7518\,
            PADOUT => \N__7517\,
            PADIN => \N__7516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2435\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__2825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7509\,
            DIN => \N__7508\,
            DOUT => \N__7507\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7509\,
            PADOUT => \N__7508\,
            PADIN => \N__7507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4890\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__4580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7500\,
            DIN => \N__7499\,
            DOUT => \N__7498\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7500\,
            PADOUT => \N__7499\,
            PADIN => \N__7498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3491\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7491\,
            DIN => \N__7490\,
            DOUT => \N__7489\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7491\,
            PADOUT => \N__7490\,
            PADIN => \N__7489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4926\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__4076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7482\,
            DIN => \N__7481\,
            DOUT => \N__7480\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7482\,
            PADOUT => \N__7481\,
            PADIN => \N__7480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7473\,
            DIN => \N__7472\,
            DOUT => \N__7471\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7473\,
            PADOUT => \N__7472\,
            PADIN => \N__7471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5015\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__2549\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7464\,
            DIN => \N__7463\,
            DOUT => \N__7462\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7464\,
            PADOUT => \N__7463\,
            PADIN => \N__7462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2434\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__3050\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7455\,
            DIN => \N__7454\,
            DOUT => \N__7453\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7455\,
            PADOUT => \N__7454\,
            PADIN => \N__7453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2409\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__3176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7446\,
            DIN => \N__7445\,
            DOUT => \N__7444\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7446\,
            PADOUT => \N__7445\,
            PADIN => \N__7444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7437\,
            DIN => \N__7436\,
            DOUT => \N__7435\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7437\,
            PADOUT => \N__7436\,
            PADIN => \N__7435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2411\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__5564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7428\,
            DIN => \N__7427\,
            DOUT => \N__7426\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7428\,
            PADOUT => \N__7427\,
            PADIN => \N__7426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4990\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__4517\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7419\,
            DIN => \N__7418\,
            DOUT => \N__7417\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7419\,
            PADOUT => \N__7418\,
            PADIN => \N__7417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7410\,
            DIN => \N__7409\,
            DOUT => \N__7408\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7410\,
            PADOUT => \N__7409\,
            PADIN => \N__7408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4788\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__3410\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7401\,
            DIN => \N__7400\,
            DOUT => \N__7399\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7401\,
            PADOUT => \N__7400\,
            PADIN => \N__7399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4948\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__4313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7392\,
            DIN => \N__7391\,
            DOUT => \N__7390\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7392\,
            PADOUT => \N__7391\,
            PADIN => \N__7390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7383\,
            DIN => \N__7382\,
            DOUT => \N__7381\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7383\,
            PADOUT => \N__7382\,
            PADIN => \N__7381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5014\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__2738\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7374\,
            DIN => \N__7373\,
            DOUT => \N__7372\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7374\,
            PADOUT => \N__7373\,
            PADIN => \N__7372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2473\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__3394\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7365\,
            DIN => \N__7364\,
            DOUT => \N__7363\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7365\,
            PADOUT => \N__7364\,
            PADIN => \N__7363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2408\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__6584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7356\,
            DIN => \N__7355\,
            DOUT => \N__7354\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7356\,
            PADOUT => \N__7355\,
            PADIN => \N__7354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4893\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__5585\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7347\,
            DIN => \N__7346\,
            DOUT => \N__7345\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7347\,
            PADOUT => \N__7346\,
            PADIN => \N__7345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2472\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__6008\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7338\,
            DIN => \N__7337\,
            DOUT => \N__7336\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7338\,
            PADOUT => \N__7337\,
            PADIN => \N__7336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2247\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__5897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7329\,
            DIN => \N__7328\,
            DOUT => \N__7327\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7329\,
            PADOUT => \N__7328\,
            PADIN => \N__7327\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4966\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3443\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7320\,
            DIN => \N__7319\,
            DOUT => \N__7318\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7320\,
            PADOUT => \N__7319\,
            PADIN => \N__7318\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4997\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__2699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7311\,
            DIN => \N__7310\,
            DOUT => \N__7309\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7311\,
            PADOUT => \N__7310\,
            PADIN => \N__7309\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2436\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3119\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7302\,
            DIN => \N__7301\,
            DOUT => \N__7300\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7302\,
            PADOUT => \N__7301\,
            PADIN => \N__7300\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2410\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__2582\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7293\,
            DIN => \N__7292\,
            DOUT => \N__7291\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7293\,
            PADOUT => \N__7292\,
            PADIN => \N__7291\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2412\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__5921\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7284\,
            DIN => \N__7283\,
            DOUT => \N__7282\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7284\,
            PADOUT => \N__7283\,
            PADIN => \N__7282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4949\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__4238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7275\,
            DIN => \N__7274\,
            DOUT => \N__7273\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7275\,
            PADOUT => \N__7274\,
            PADIN => \N__7273\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3539\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7266\,
            DIN => \N__7265\,
            DOUT => \N__7264\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7266\,
            PADOUT => \N__7265\,
            PADIN => \N__7264\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4830\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__5378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7257\,
            DIN => \N__7256\,
            DOUT => \N__7255\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7257\,
            PADOUT => \N__7256\,
            PADIN => \N__7255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4999\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__3671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7248\,
            DIN => \N__7247\,
            DOUT => \N__7246\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7248\,
            PADOUT => \N__7247\,
            PADIN => \N__7246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7239\,
            DIN => \N__7238\,
            DOUT => \N__7237\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7239\,
            PADOUT => \N__7238\,
            PADIN => \N__7237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2474\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__3650\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7230\,
            DIN => \N__7229\,
            DOUT => \N__7228\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7230\,
            PADOUT => \N__7229\,
            PADIN => \N__7228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2452\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__3251\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7221\,
            DIN => \N__7220\,
            DOUT => \N__7219\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7221\,
            PADOUT => \N__7220\,
            PADIN => \N__7219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2406\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__3743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7212\,
            DIN => \N__7211\,
            DOUT => \N__7210\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7212\,
            PADOUT => \N__7211\,
            PADIN => \N__7210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7203\,
            DIN => \N__7202\,
            DOUT => \N__7201\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7203\,
            PADOUT => \N__7202\,
            PADIN => \N__7201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2414\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__2642\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7194\,
            DIN => \N__7193\,
            DOUT => \N__7192\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7194\,
            PADOUT => \N__7193\,
            PADIN => \N__7192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7185\,
            DIN => \N__7184\,
            DOUT => \N__7183\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7185\,
            PADOUT => \N__7184\,
            PADIN => \N__7183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4832\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3851\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7176\,
            DIN => \N__7175\,
            DOUT => \N__7174\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7176\,
            PADOUT => \N__7175\,
            PADIN => \N__7174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4789\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__5390\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7167\,
            DIN => \N__7166\,
            DOUT => \N__7165\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7167\,
            PADOUT => \N__7166\,
            PADIN => \N__7165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7158\,
            DIN => \N__7157\,
            DOUT => \N__7156\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7158\,
            PADOUT => \N__7157\,
            PADIN => \N__7156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7149\,
            DIN => \N__7148\,
            DOUT => \N__7147\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7149\,
            PADOUT => \N__7148\,
            PADIN => \N__7147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4998\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__5462\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7140\,
            DIN => \N__7139\,
            DOUT => \N__7138\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7140\,
            PADOUT => \N__7139\,
            PADIN => \N__7138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2437\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__6923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7131\,
            DIN => \N__7130\,
            DOUT => \N__7129\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7131\,
            PADOUT => \N__7130\,
            PADIN => \N__7129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2361\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__6161\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7122\,
            DIN => \N__7121\,
            DOUT => \N__7120\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7122\,
            PADOUT => \N__7121\,
            PADIN => \N__7120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4989\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__4388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7113\,
            DIN => \N__7112\,
            DOUT => \N__7111\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7113\,
            PADOUT => \N__7112\,
            PADIN => \N__7111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2360\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__3781\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7104\,
            DIN => \N__7103\,
            DOUT => \N__7102\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7104\,
            PADOUT => \N__7103\,
            PADIN => \N__7102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7095\,
            DIN => \N__7094\,
            DOUT => \N__7093\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7095\,
            PADOUT => \N__7094\,
            PADIN => \N__7093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5023\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__2198\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7086\,
            DIN => \N__7085\,
            DOUT => \N__7084\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7086\,
            PADOUT => \N__7085\,
            PADIN => \N__7084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4965\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__5429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7077\,
            DIN => \N__7076\,
            DOUT => \N__7075\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7077\,
            PADOUT => \N__7076\,
            PADIN => \N__7075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7068\,
            DIN => \N__7067\,
            DOUT => \N__7066\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7068\,
            PADOUT => \N__7067\,
            PADIN => \N__7066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2451\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__2984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7059\,
            DIN => \N__7058\,
            DOUT => \N__7057\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7059\,
            PADOUT => \N__7058\,
            PADIN => \N__7057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2413\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__3212\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7050\,
            DIN => \N__7049\,
            DOUT => \N__7048\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7050\,
            PADOUT => \N__7049\,
            PADIN => \N__7048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7041\,
            DIN => \N__7040\,
            DOUT => \N__7039\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7041\,
            PADOUT => \N__7040\,
            PADIN => \N__7039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2489\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7032\,
            DIN => \N__7031\,
            DOUT => \N__7030\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7032\,
            PADOUT => \N__7031\,
            PADIN => \N__7030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4879\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__2663\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7023\,
            DIN => \N__7022\,
            DOUT => \N__7021\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7023\,
            PADOUT => \N__7022\,
            PADIN => \N__7021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4891\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__4451\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7014\,
            DIN => \N__7013\,
            DOUT => \N__7012\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7014\,
            PADOUT => \N__7013\,
            PADIN => \N__7012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7005\,
            DIN => \N__7004\,
            DOUT => \N__7003\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7005\,
            PADOUT => \N__7004\,
            PADIN => \N__7003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2449\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__5840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6996\,
            DIN => \N__6995\,
            DOUT => \N__6994\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6996\,
            PADOUT => \N__6995\,
            PADIN => \N__6994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3490\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6987\,
            DIN => \N__6986\,
            DOUT => \N__6985\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6987\,
            PADOUT => \N__6986\,
            PADIN => \N__6985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4831\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__5408\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6978\,
            DIN => \N__6977\,
            DOUT => \N__6976\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6978\,
            PADOUT => \N__6977\,
            PADIN => \N__6976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2309\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__6218\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6969\,
            DIN => \N__6968\,
            DOUT => \N__6967\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6969\,
            PADOUT => \N__6968\,
            PADIN => \N__6967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2297\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__3887\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6960\,
            DIN => \N__6959\,
            DOUT => \N__6958\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6960\,
            PADOUT => \N__6959\,
            PADIN => \N__6958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4950\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__6515\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6951\,
            DIN => \N__6950\,
            DOUT => \N__6949\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6951\,
            PADOUT => \N__6950\,
            PADIN => \N__6949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6942\,
            DIN => \N__6941\,
            DOUT => \N__6940\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6942\,
            PADOUT => \N__6941\,
            PADIN => \N__6940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5024\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__3704\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1771\ : IoInMux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1769\ : IoSpan4Mux
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1768\ : Span4Mux_s3_h
    port map (
            O => \N__6914\,
            I => \N__6910\
        );

    \I__1767\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1766\ : Sp12to4
    port map (
            O => \N__6910\,
            I => \N__6904\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__6907\,
            I => \N__6901\
        );

    \I__1764\ : Span12Mux_v
    port map (
            O => \N__6904\,
            I => \N__6898\
        );

    \I__1763\ : Span12Mux_v
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__1762\ : Span12Mux_h
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1761\ : Span12Mux_v
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1760\ : Span12Mux_h
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1759\ : Span12Mux_h
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__6886\,
            I => \D_LL_040_in_5\
        );

    \I__1757\ : Odrv12
    port map (
            O => \N__6883\,
            I => \D_LL_040_in_5\
        );

    \I__1756\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6874\
        );

    \I__1755\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6871\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__6874\,
            I => \N__6862\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6862\
        );

    \I__1752\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6859\
        );

    \I__1751\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6856\
        );

    \I__1750\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6853\
        );

    \I__1749\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6850\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__6862\,
            I => \N__6841\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__6859\,
            I => \N__6841\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6841\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6834\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__6850\,
            I => \N__6834\
        );

    \I__1743\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6829\
        );

    \I__1742\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6819\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__6841\,
            I => \N__6810\
        );

    \I__1740\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6807\
        );

    \I__1739\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6804\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6801\
        );

    \I__1737\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6798\
        );

    \I__1736\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6794\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__6829\,
            I => \N__6791\
        );

    \I__1734\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6788\
        );

    \I__1733\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6785\
        );

    \I__1732\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6782\
        );

    \I__1731\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6779\
        );

    \I__1730\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6776\
        );

    \I__1729\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6773\
        );

    \I__1728\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6766\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__6819\,
            I => \N__6763\
        );

    \I__1726\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6760\
        );

    \I__1725\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6757\
        );

    \I__1724\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6754\
        );

    \I__1723\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6751\
        );

    \I__1722\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6746\
        );

    \I__1721\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6743\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__6810\,
            I => \N__6736\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6736\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6736\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__6801\,
            I => \N__6731\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6731\
        );

    \I__1715\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6728\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6725\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__6791\,
            I => \N__6712\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6712\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6712\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__6782\,
            I => \N__6712\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6712\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__6776\,
            I => \N__6712\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__6773\,
            I => \N__6709\
        );

    \I__1706\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6706\
        );

    \I__1705\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6703\
        );

    \I__1704\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6700\
        );

    \I__1703\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6697\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__6766\,
            I => \N__6694\
        );

    \I__1701\ : Sp12to4
    port map (
            O => \N__6763\,
            I => \N__6689\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__6760\,
            I => \N__6689\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__6757\,
            I => \N__6684\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6684\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__6751\,
            I => \N__6681\
        );

    \I__1696\ : InMux
    port map (
            O => \N__6750\,
            I => \N__6678\
        );

    \I__1695\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6675\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__6746\,
            I => \N__6670\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6670\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__6736\,
            I => \N__6663\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__6731\,
            I => \N__6663\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6663\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__6725\,
            I => \N__6658\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__6712\,
            I => \N__6658\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__6709\,
            I => \N__6653\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__6706\,
            I => \N__6653\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N__6648\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__6700\,
            I => \N__6648\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__6697\,
            I => \N__6645\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__6694\,
            I => \N__6642\
        );

    \I__1681\ : Span12Mux_v
    port map (
            O => \N__6689\,
            I => \N__6637\
        );

    \I__1680\ : Span12Mux_s10_v
    port map (
            O => \N__6684\,
            I => \N__6637\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__6681\,
            I => \N__6634\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__6678\,
            I => \N__6629\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6629\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__6670\,
            I => \N__6624\
        );

    \I__1675\ : Span4Mux_v
    port map (
            O => \N__6663\,
            I => \N__6624\
        );

    \I__1674\ : Span4Mux_h
    port map (
            O => \N__6658\,
            I => \N__6615\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__6653\,
            I => \N__6615\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__6648\,
            I => \N__6615\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__6645\,
            I => \N__6615\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__6642\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__6637\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__6634\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1667\ : Odrv12
    port map (
            O => \N__6629\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__6624\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__6615\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1664\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1662\ : Span4Mux_v
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1661\ : Sp12to4
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1660\ : Span12Mux_h
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1659\ : Odrv12
    port map (
            O => \N__6587\,
            I => \D_UM_040_in_5\
        );

    \I__1658\ : IoInMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1656\ : Span4Mux_s2_v
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__1654\ : Sp12to4
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__1653\ : Span12Mux_h
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1652\ : Odrv12
    port map (
            O => \N__6566\,
            I => \un1_D_UM_040_5\
        );

    \I__1651\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6557\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__6557\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1648\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6548\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__6548\,
            I => \N__6544\
        );

    \I__1645\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__6544\,
            I => \N__6535\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__1642\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6532\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__6535\,
            I => \N__6527\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__6532\,
            I => \N__6527\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1638\ : Sp12to4
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1637\ : Span12Mux_h
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__6518\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1635\ : IoInMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1633\ : Span4Mux_s3_v
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__6506\,
            I => \N__6503\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__6497\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1628\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__6488\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__6479\,
            I => \N__6475\
        );

    \I__1622\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__6475\,
            I => \N__6466\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__1619\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6463\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__6466\,
            I => \N__6460\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__6460\,
            I => \N__6454\
        );

    \I__1615\ : Span12Mux_h
    port map (
            O => \N__6457\,
            I => \N__6451\
        );

    \I__1614\ : Sp12to4
    port map (
            O => \N__6454\,
            I => \N__6448\
        );

    \I__1613\ : Span12Mux_h
    port map (
            O => \N__6451\,
            I => \N__6445\
        );

    \I__1612\ : Span12Mux_h
    port map (
            O => \N__6448\,
            I => \N__6442\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__6445\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__6442\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1609\ : IoInMux
    port map (
            O => \N__6437\,
            I => \N__6434\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6431\
        );

    \I__1607\ : Span12Mux_s7_v
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__1606\ : Span12Mux_h
    port map (
            O => \N__6428\,
            I => \N__6425\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__6425\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1604\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__6416\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1601\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__6404\,
            I => \N__6399\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6396\
        );

    \I__1596\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6393\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__6399\,
            I => \N__6390\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6387\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__6393\,
            I => \N__6384\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__6390\,
            I => \N__6377\
        );

    \I__1591\ : Span12Mux_h
    port map (
            O => \N__6387\,
            I => \N__6377\
        );

    \I__1590\ : Span12Mux_s9_v
    port map (
            O => \N__6384\,
            I => \N__6377\
        );

    \I__1589\ : Span12Mux_h
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__6374\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6365\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6365\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__6362\,
            I => \N__6358\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6352\
        );

    \I__1582\ : Sp12to4
    port map (
            O => \N__6358\,
            I => \N__6344\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6335\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6332\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6329\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6352\,
            I => \N__6326\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6321\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6321\
        );

    \I__1575\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6316\
        );

    \I__1574\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6316\
        );

    \I__1573\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6313\
        );

    \I__1572\ : Span12Mux_h
    port map (
            O => \N__6344\,
            I => \N__6308\
        );

    \I__1571\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6305\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6296\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6296\
        );

    \I__1568\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6296\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6296\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6293\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6335\,
            I => \N__6286\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6332\,
            I => \N__6286\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__6329\,
            I => \N__6286\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__6326\,
            I => \N__6277\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6277\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6277\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6277\
        );

    \I__1558\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6272\
        );

    \I__1557\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6272\
        );

    \I__1556\ : Span12Mux_v
    port map (
            O => \N__6308\,
            I => \N__6263\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__6305\,
            I => \N__6263\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6263\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6260\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__6286\,
            I => \N__6255\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__6277\,
            I => \N__6255\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__6272\,
            I => \N__6252\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6247\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6247\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__6263\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__6255\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__6252\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6247\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1542\ : IoInMux
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1540\ : Span4Mux_s3_v
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1539\ : Sp12to4
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__1538\ : Span12Mux_h
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1537\ : Odrv12
    port map (
            O => \N__6221\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1536\ : IoInMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6211\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6208\
        );

    \I__1533\ : IoSpan4Mux
    port map (
            O => \N__6211\,
            I => \N__6205\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6202\
        );

    \I__1531\ : Span4Mux_s2_h
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__1529\ : Sp12to4
    port map (
            O => \N__6199\,
            I => \N__6193\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__6196\,
            I => \N__6190\
        );

    \I__1527\ : Span12Mux_h
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__6190\,
            I => \N__6184\
        );

    \I__1525\ : Span12Mux_h
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__1524\ : Span12Mux_v
    port map (
            O => \N__6184\,
            I => \N__6178\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__6181\,
            I => \D_LL_040_in_0\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__6178\,
            I => \D_LL_040_in_0\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__6164\,
            I => \D_UM_040_in_0\
        );

    \I__1517\ : IoInMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1515\ : IoSpan4Mux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__1514\ : Sp12to4
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__1513\ : Span12Mux_h
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1512\ : Odrv12
    port map (
            O => \N__6146\,
            I => \un1_D_UM_040_0\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6136\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6133\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__1505\ : Span4Mux_v
    port map (
            O => \N__6127\,
            I => \N__6121\
        );

    \I__1504\ : Sp12to4
    port map (
            O => \N__6124\,
            I => \N__6116\
        );

    \I__1503\ : Sp12to4
    port map (
            O => \N__6121\,
            I => \N__6116\
        );

    \I__1502\ : Span12Mux_h
    port map (
            O => \N__6116\,
            I => \N__6113\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__6113\,
            I => \SIZ_c_0\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6106\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6103\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6106\,
            I => \N__6100\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6103\,
            I => \N__6097\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__6100\,
            I => \N__6092\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__6097\,
            I => \N__6092\
        );

    \I__1494\ : Sp12to4
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1493\ : Span12Mux_h
    port map (
            O => \N__6089\,
            I => \N__6086\
        );

    \I__1492\ : Odrv12
    port map (
            O => \N__6086\,
            I => \SIZ_c_1\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6080\,
            I => \N__6077\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__6077\,
            I => \N__6074\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__6074\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1487\ : IoInMux
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6065\
        );

    \I__1485\ : IoSpan4Mux
    port map (
            O => \N__6065\,
            I => \N__6061\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__1483\ : IoSpan4Mux
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__1481\ : Span4Mux_s2_h
    port map (
            O => \N__6055\,
            I => \N__6049\
        );

    \I__1480\ : Span4Mux_v
    port map (
            O => \N__6052\,
            I => \N__6046\
        );

    \I__1479\ : Sp12to4
    port map (
            O => \N__6049\,
            I => \N__6043\
        );

    \I__1478\ : Sp12to4
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__1477\ : Span12Mux_h
    port map (
            O => \N__6043\,
            I => \N__6037\
        );

    \I__1476\ : Span12Mux_h
    port map (
            O => \N__6040\,
            I => \N__6034\
        );

    \I__1475\ : Span12Mux_h
    port map (
            O => \N__6037\,
            I => \N__6031\
        );

    \I__1474\ : Span12Mux_v
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__1473\ : Odrv12
    port map (
            O => \N__6031\,
            I => \D_LM_040_in_3\
        );

    \I__1472\ : Odrv12
    port map (
            O => \N__6028\,
            I => \D_LM_040_in_3\
        );

    \I__1471\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__1469\ : Span12Mux_v
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1468\ : Span12Mux_h
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__6011\,
            I => \D_UU_040_in_3\
        );

    \I__1466\ : IoInMux
    port map (
            O => \N__6008\,
            I => \N__6005\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6005\,
            I => \N__6002\
        );

    \I__1464\ : Span4Mux_s3_v
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__1463\ : Span4Mux_h
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__1460\ : Span4Mux_h
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__5987\,
            I => \un1_D_UU_040_3\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1456\ : Span4Mux_s3_h
    port map (
            O => \N__5978\,
            I => \N__5974\
        );

    \I__1455\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5971\
        );

    \I__1454\ : Sp12to4
    port map (
            O => \N__5974\,
            I => \N__5968\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__1452\ : Span12Mux_v
    port map (
            O => \N__5968\,
            I => \N__5962\
        );

    \I__1451\ : Span12Mux_v
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__1450\ : Span12Mux_h
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__1449\ : Span12Mux_v
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__1448\ : Span12Mux_h
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__1447\ : Span12Mux_h
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__5950\,
            I => \D_LL_040_in_1\
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__5947\,
            I => \D_LL_040_in_1\
        );

    \I__1444\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__1441\ : Sp12to4
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__1440\ : Span12Mux_h
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__1439\ : Span12Mux_v
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__5924\,
            I => \D_UM_040_in_1\
        );

    \I__1437\ : IoInMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__1435\ : Span4Mux_s3_h
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__1432\ : Span4Mux_h
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__5900\,
            I => \un1_D_UM_040_1\
        );

    \I__1429\ : IoInMux
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1427\ : Span4Mux_s3_h
    port map (
            O => \N__5891\,
            I => \N__5887\
        );

    \I__1426\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5884\
        );

    \I__1425\ : Sp12to4
    port map (
            O => \N__5887\,
            I => \N__5881\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__5884\,
            I => \N__5878\
        );

    \I__1423\ : Span12Mux_v
    port map (
            O => \N__5881\,
            I => \N__5875\
        );

    \I__1422\ : Span12Mux_v
    port map (
            O => \N__5878\,
            I => \N__5872\
        );

    \I__1421\ : Span12Mux_h
    port map (
            O => \N__5875\,
            I => \N__5869\
        );

    \I__1420\ : Span12Mux_v
    port map (
            O => \N__5872\,
            I => \N__5866\
        );

    \I__1419\ : Span12Mux_h
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__1418\ : Span12Mux_h
    port map (
            O => \N__5866\,
            I => \N__5860\
        );

    \I__1417\ : Odrv12
    port map (
            O => \N__5863\,
            I => \D_LM_040_in_1\
        );

    \I__1416\ : Odrv12
    port map (
            O => \N__5860\,
            I => \D_LM_040_in_1\
        );

    \I__1415\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__1413\ : Span12Mux_v
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__1412\ : Span12Mux_h
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__1411\ : Odrv12
    port map (
            O => \N__5843\,
            I => \D_UU_040_in_1\
        );

    \I__1410\ : IoInMux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__1408\ : IoSpan4Mux
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__1407\ : Span4Mux_s2_h
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__1406\ : Sp12to4
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__1405\ : Span12Mux_h
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__5822\,
            I => \un1_D_UU_040_1\
        );

    \I__1403\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__5813\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1400\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__1398\ : Sp12to4
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1397\ : Span12Mux_v
    port map (
            O => \N__5801\,
            I => \N__5797\
        );

    \I__1396\ : IoInMux
    port map (
            O => \N__5800\,
            I => \N__5794\
        );

    \I__1395\ : Span12Mux_h
    port map (
            O => \N__5797\,
            I => \N__5791\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5788\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__5791\,
            I => \A_AMIGA_c_1\
        );

    \I__1392\ : Odrv12
    port map (
            O => \N__5788\,
            I => \A_AMIGA_c_1\
        );

    \I__1391\ : CEMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__5780\,
            I => \N__5775\
        );

    \I__1389\ : CEMux
    port map (
            O => \N__5779\,
            I => \N__5772\
        );

    \I__1388\ : CEMux
    port map (
            O => \N__5778\,
            I => \N__5769\
        );

    \I__1387\ : Span4Mux_v
    port map (
            O => \N__5775\,
            I => \N__5766\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__5772\,
            I => \N__5763\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5760\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__5766\,
            I => \N__5757\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__5763\,
            I => \N__5752\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__5760\,
            I => \N__5752\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__5757\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__5752\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1379\ : SRMux
    port map (
            O => \N__5747\,
            I => \N__5744\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5739\
        );

    \I__1377\ : SRMux
    port map (
            O => \N__5743\,
            I => \N__5736\
        );

    \I__1376\ : SRMux
    port map (
            O => \N__5742\,
            I => \N__5733\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__5739\,
            I => \N__5730\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__5736\,
            I => \N__5727\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5724\
        );

    \I__1372\ : Span4Mux_h
    port map (
            O => \N__5730\,
            I => \N__5720\
        );

    \I__1371\ : Span4Mux_h
    port map (
            O => \N__5727\,
            I => \N__5715\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__5724\,
            I => \N__5715\
        );

    \I__1369\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5712\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__5720\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__5715\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5712\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5698\
        );

    \I__1363\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5691\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5695\,
            I => \N__5688\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5685\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__5691\,
            I => \N__5682\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__5688\,
            I => \N__5677\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__5685\,
            I => \N__5677\
        );

    \I__1356\ : Sp12to4
    port map (
            O => \N__5682\,
            I => \N__5674\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__1354\ : Span12Mux_h
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__1352\ : Span12Mux_v
    port map (
            O => \N__5668\,
            I => \N__5660\
        );

    \I__1351\ : Span12Mux_h
    port map (
            O => \N__5665\,
            I => \N__5660\
        );

    \I__1350\ : Odrv12
    port map (
            O => \N__5660\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1349\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__5654\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1347\ : IoInMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1345\ : Span4Mux_s2_h
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__1344\ : Sp12to4
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__1343\ : Span12Mux_s9_v
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1342\ : Span12Mux_h
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__5633\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5627\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1338\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__5618\,
            I => \N__5614\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5611\
        );

    \I__1334\ : Span4Mux_v
    port map (
            O => \N__5614\,
            I => \N__5605\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5602\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__5605\,
            I => \N__5597\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__5602\,
            I => \N__5597\
        );

    \I__1329\ : Span4Mux_v
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1328\ : Sp12to4
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__1327\ : Span12Mux_h
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__5588\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1325\ : IoInMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1323\ : IoSpan4Mux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__1322\ : IoSpan4Mux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1321\ : Span4Mux_s3_h
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__1320\ : Sp12to4
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__1319\ : Odrv12
    port map (
            O => \N__5567\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1318\ : IoInMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1316\ : IoSpan4Mux
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1315\ : IoSpan4Mux
    port map (
            O => \N__5555\,
            I => \N__5551\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__1313\ : Span4Mux_s2_h
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__1311\ : Sp12to4
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__1309\ : Span12Mux_h
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__1308\ : Span12Mux_v
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__1306\ : Span12Mux_h
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__5527\,
            I => \D_LM_040_in_5\
        );

    \I__1304\ : Odrv12
    port map (
            O => \N__5524\,
            I => \D_LM_040_in_5\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__1301\ : Sp12to4
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__1300\ : Span12Mux_v
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__1299\ : Span12Mux_h
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__5504\,
            I => \D_UU_040_in_5\
        );

    \I__1297\ : IoInMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__1295\ : Span4Mux_s3_h
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__1293\ : Sp12to4
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__1292\ : Span12Mux_h
    port map (
            O => \N__5486\,
            I => \N__5483\
        );

    \I__1291\ : Odrv12
    port map (
            O => \N__5483\,
            I => \un1_D_UU_040_5\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1287\ : Sp12to4
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__1286\ : Span12Mux_h
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__5465\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__1282\ : IoSpan4Mux
    port map (
            O => \N__5456\,
            I => \N__5453\
        );

    \I__1281\ : Span4Mux_s0_h
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__1280\ : Sp12to4
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__1279\ : Span12Mux_h
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__5444\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__1275\ : Span12Mux_h
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__5432\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__1273\ : IoInMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__1271\ : IoSpan4Mux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__1270\ : Span4Mux_s0_h
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__1269\ : Sp12to4
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__1268\ : Span12Mux_h
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__5411\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__1266\ : IoInMux
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__1264\ : IoSpan4Mux
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__1263\ : Span4Mux_s3_h
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__5393\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1260\ : IoInMux
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__1258\ : Span12Mux_s7_h
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__1257\ : Odrv12
    port map (
            O => \N__5381\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1256\ : IoInMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__1254\ : Span4Mux_s3_h
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__1252\ : Sp12to4
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__1251\ : Odrv12
    port map (
            O => \N__5363\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5352\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5349\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5346\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__5352\,
            I => \N__5343\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5338\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5338\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__5343\,
            I => \N__5333\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__5338\,
            I => \N__5333\
        );

    \I__1241\ : Sp12to4
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__1240\ : Span12Mux_h
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__1239\ : Span12Mux_v
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__1238\ : Odrv12
    port map (
            O => \N__5324\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__5315\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5303\,
            I => \N__5299\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5296\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5299\,
            I => \N__5292\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5296\,
            I => \N__5289\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5286\
        );

    \I__1226\ : Sp12to4
    port map (
            O => \N__5292\,
            I => \N__5281\
        );

    \I__1225\ : Span12Mux_v
    port map (
            O => \N__5289\,
            I => \N__5281\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5278\
        );

    \I__1223\ : Span12Mux_h
    port map (
            O => \N__5281\,
            I => \N__5275\
        );

    \I__1222\ : Span12Mux_h
    port map (
            O => \N__5278\,
            I => \N__5272\
        );

    \I__1221\ : Odrv12
    port map (
            O => \N__5275\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__5272\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5264\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5254\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__1214\ : Span4Mux_h
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5245\
        );

    \I__1212\ : Sp12to4
    port map (
            O => \N__5248\,
            I => \N__5241\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__5245\,
            I => \N__5238\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5235\
        );

    \I__1209\ : Span12Mux_v
    port map (
            O => \N__5241\,
            I => \N__5232\
        );

    \I__1208\ : Sp12to4
    port map (
            O => \N__5238\,
            I => \N__5227\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5235\,
            I => \N__5227\
        );

    \I__1206\ : Span12Mux_h
    port map (
            O => \N__5232\,
            I => \N__5224\
        );

    \I__1205\ : Span12Mux_h
    port map (
            O => \N__5227\,
            I => \N__5221\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__5224\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__5221\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1202\ : IoInMux
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__1200\ : Sp12to4
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__1199\ : Span12Mux_v
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__5204\,
            I => \TAn_0_i\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1195\ : CEMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5186\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\
        );

    \I__1191\ : SRMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5180\,
            I => \N__5176\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5173\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__5176\,
            I => \N__5170\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5173\,
            I => \RESETn_c_i\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__5170\,
            I => \RESETn_c_i\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5154\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5154\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5154\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5151\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \N__5148\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5143\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5143\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5140\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__5143\,
            I => \N__5137\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__1175\ : Sp12to4
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__1173\ : Span12Mux_h
    port map (
            O => \N__5131\,
            I => \N__5125\
        );

    \I__1172\ : Sp12to4
    port map (
            O => \N__5128\,
            I => \N__5122\
        );

    \I__1171\ : Span12Mux_v
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__1170\ : Span12Mux_v
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__1169\ : Odrv12
    port map (
            O => \N__5119\,
            I => \TACKn_c\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__5116\,
            I => \TACKn_c\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__5111\,
            I => \N__5107\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5096\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5093\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5090\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5081\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5081\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5081\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5081\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5074\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5074\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5074\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5096\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5090\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5074\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5054\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5051\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5046\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5046\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5039\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5039\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5039\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5046\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5027\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5027\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__1138\ : IoInMux
    port map (
            O => \N__5024\,
            I => \N__5019\
        );

    \I__1137\ : IoInMux
    port map (
            O => \N__5023\,
            I => \N__5016\
        );

    \I__1136\ : IoInMux
    port map (
            O => \N__5022\,
            I => \N__5011\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5006\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5016\,
            I => \N__5006\
        );

    \I__1133\ : IoInMux
    port map (
            O => \N__5015\,
            I => \N__5003\
        );

    \I__1132\ : IoInMux
    port map (
            O => \N__5014\,
            I => \N__5000\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__4992\
        );

    \I__1130\ : IoSpan4Mux
    port map (
            O => \N__5006\,
            I => \N__4982\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__4982\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5000\,
            I => \N__4982\
        );

    \I__1127\ : IoInMux
    port map (
            O => \N__4999\,
            I => \N__4979\
        );

    \I__1126\ : IoInMux
    port map (
            O => \N__4998\,
            I => \N__4976\
        );

    \I__1125\ : IoInMux
    port map (
            O => \N__4997\,
            I => \N__4973\
        );

    \I__1124\ : IoInMux
    port map (
            O => \N__4996\,
            I => \N__4970\
        );

    \I__1123\ : IoInMux
    port map (
            O => \N__4995\,
            I => \N__4967\
        );

    \I__1122\ : Span4Mux_s3_v
    port map (
            O => \N__4992\,
            I => \N__4962\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4959\
        );

    \I__1120\ : IoInMux
    port map (
            O => \N__4990\,
            I => \N__4955\
        );

    \I__1119\ : IoInMux
    port map (
            O => \N__4989\,
            I => \N__4952\
        );

    \I__1118\ : IoSpan4Mux
    port map (
            O => \N__4982\,
            I => \N__4933\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4933\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__4976\,
            I => \N__4933\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4933\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__4970\,
            I => \N__4933\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4933\
        );

    \I__1112\ : IoInMux
    port map (
            O => \N__4966\,
            I => \N__4930\
        );

    \I__1111\ : IoInMux
    port map (
            O => \N__4965\,
            I => \N__4927\
        );

    \I__1110\ : Span4Mux_h
    port map (
            O => \N__4962\,
            I => \N__4923\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4920\
        );

    \I__1108\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4917\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4912\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4912\
        );

    \I__1105\ : IoInMux
    port map (
            O => \N__4951\,
            I => \N__4909\
        );

    \I__1104\ : IoInMux
    port map (
            O => \N__4950\,
            I => \N__4906\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__4949\,
            I => \N__4903\
        );

    \I__1102\ : IoInMux
    port map (
            O => \N__4948\,
            I => \N__4900\
        );

    \I__1101\ : IoInMux
    port map (
            O => \N__4947\,
            I => \N__4897\
        );

    \I__1100\ : IoInMux
    port map (
            O => \N__4946\,
            I => \N__4894\
        );

    \I__1099\ : IoSpan4Mux
    port map (
            O => \N__4933\,
            I => \N__4883\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__4930\,
            I => \N__4883\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__4927\,
            I => \N__4883\
        );

    \I__1096\ : IoInMux
    port map (
            O => \N__4926\,
            I => \N__4880\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__4923\,
            I => \N__4876\
        );

    \I__1094\ : Span4Mux_v
    port map (
            O => \N__4920\,
            I => \N__4873\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4870\
        );

    \I__1092\ : IoSpan4Mux
    port map (
            O => \N__4912\,
            I => \N__4854\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4854\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4906\,
            I => \N__4854\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4854\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4854\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4854\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__4894\,
            I => \N__4854\
        );

    \I__1085\ : IoInMux
    port map (
            O => \N__4893\,
            I => \N__4851\
        );

    \I__1084\ : IoInMux
    port map (
            O => \N__4892\,
            I => \N__4848\
        );

    \I__1083\ : IoInMux
    port map (
            O => \N__4891\,
            I => \N__4845\
        );

    \I__1082\ : IoInMux
    port map (
            O => \N__4890\,
            I => \N__4842\
        );

    \I__1081\ : IoSpan4Mux
    port map (
            O => \N__4883\,
            I => \N__4839\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4836\
        );

    \I__1079\ : IoInMux
    port map (
            O => \N__4879\,
            I => \N__4833\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__4876\,
            I => \N__4825\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__4873\,
            I => \N__4825\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__4870\,
            I => \N__4822\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__4869\,
            I => \N__4819\
        );

    \I__1074\ : IoSpan4Mux
    port map (
            O => \N__4854\,
            I => \N__4808\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__4851\,
            I => \N__4808\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4848\,
            I => \N__4808\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4808\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4842\,
            I => \N__4808\
        );

    \I__1069\ : IoSpan4Mux
    port map (
            O => \N__4839\,
            I => \N__4802\
        );

    \I__1068\ : IoSpan4Mux
    port map (
            O => \N__4836\,
            I => \N__4802\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__4833\,
            I => \N__4799\
        );

    \I__1066\ : IoInMux
    port map (
            O => \N__4832\,
            I => \N__4796\
        );

    \I__1065\ : IoInMux
    port map (
            O => \N__4831\,
            I => \N__4793\
        );

    \I__1064\ : IoInMux
    port map (
            O => \N__4830\,
            I => \N__4790\
        );

    \I__1063\ : Sp12to4
    port map (
            O => \N__4825\,
            I => \N__4785\
        );

    \I__1062\ : Sp12to4
    port map (
            O => \N__4822\,
            I => \N__4782\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4779\
        );

    \I__1060\ : IoSpan4Mux
    port map (
            O => \N__4808\,
            I => \N__4776\
        );

    \I__1059\ : IoInMux
    port map (
            O => \N__4807\,
            I => \N__4773\
        );

    \I__1058\ : IoSpan4Mux
    port map (
            O => \N__4802\,
            I => \N__4762\
        );

    \I__1057\ : IoSpan4Mux
    port map (
            O => \N__4799\,
            I => \N__4762\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4762\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4762\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4790\,
            I => \N__4762\
        );

    \I__1053\ : IoInMux
    port map (
            O => \N__4789\,
            I => \N__4759\
        );

    \I__1052\ : IoInMux
    port map (
            O => \N__4788\,
            I => \N__4756\
        );

    \I__1051\ : Span12Mux_h
    port map (
            O => \N__4785\,
            I => \N__4753\
        );

    \I__1050\ : Span12Mux_h
    port map (
            O => \N__4782\,
            I => \N__4748\
        );

    \I__1049\ : Span12Mux_s11_v
    port map (
            O => \N__4779\,
            I => \N__4748\
        );

    \I__1048\ : IoSpan4Mux
    port map (
            O => \N__4776\,
            I => \N__4743\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4773\,
            I => \N__4743\
        );

    \I__1046\ : IoSpan4Mux
    port map (
            O => \N__4762\,
            I => \N__4738\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4759\,
            I => \N__4738\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4756\,
            I => \N__4735\
        );

    \I__1043\ : Odrv12
    port map (
            O => \N__4753\,
            I => \RnW_c\
        );

    \I__1042\ : Odrv12
    port map (
            O => \N__4748\,
            I => \RnW_c\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__4743\,
            I => \RnW_c\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__4738\,
            I => \RnW_c\
        );

    \I__1039\ : Odrv12
    port map (
            O => \N__4735\,
            I => \RnW_c\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__4724\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \N__4712\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__4719\,
            I => \N__4706\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4698\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4698\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4698\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4695\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4692\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4687\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4687\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__4705\,
            I => \N__4684\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4698\,
            I => \N__4680\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4695\,
            I => \N__4677\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4692\,
            I => \N__4672\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4687\,
            I => \N__4672\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4669\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4666\
        );

    \I__1020\ : Span4Mux_v
    port map (
            O => \N__4680\,
            I => \N__4661\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__4677\,
            I => \N__4661\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__4672\,
            I => \N__4654\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4654\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4666\,
            I => \N__4654\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__4661\,
            I => \N__4651\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__4654\,
            I => \N__4648\
        );

    \I__1013\ : Sp12to4
    port map (
            O => \N__4651\,
            I => \N__4645\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__4648\,
            I => \N__4642\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__4645\,
            I => \N__4637\
        );

    \I__1010\ : Sp12to4
    port map (
            O => \N__4642\,
            I => \N__4637\
        );

    \I__1009\ : Span12Mux_v
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__4634\,
            I => \RESETn_c\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4628\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4622\,
            I => \N__4617\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4614\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4611\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__4617\,
            I => \N__4608\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4603\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4611\,
            I => \N__4603\
        );

    \I__998\ : Sp12to4
    port map (
            O => \N__4608\,
            I => \N__4600\
        );

    \I__997\ : Span4Mux_v
    port map (
            O => \N__4603\,
            I => \N__4597\
        );

    \I__996\ : Span12Mux_h
    port map (
            O => \N__4600\,
            I => \N__4594\
        );

    \I__995\ : Sp12to4
    port map (
            O => \N__4597\,
            I => \N__4591\
        );

    \I__994\ : Span12Mux_v
    port map (
            O => \N__4594\,
            I => \N__4588\
        );

    \I__993\ : Span12Mux_h
    port map (
            O => \N__4591\,
            I => \N__4585\
        );

    \I__992\ : Odrv12
    port map (
            O => \N__4588\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__4585\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__990\ : IoInMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__988\ : Span4Mux_s3_h
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__987\ : Span4Mux_h
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__986\ : Sp12to4
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__985\ : Span12Mux_s9_v
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__4562\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__983\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4556\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__981\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4550\,
            I => \N__4545\
        );

    \I__979\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4542\
        );

    \I__978\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4539\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__4545\,
            I => \N__4536\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4542\,
            I => \N__4531\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4539\,
            I => \N__4531\
        );

    \I__974\ : Span4Mux_v
    port map (
            O => \N__4536\,
            I => \N__4526\
        );

    \I__973\ : Span4Mux_v
    port map (
            O => \N__4531\,
            I => \N__4526\
        );

    \I__972\ : Sp12to4
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__971\ : Span12Mux_h
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__4520\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__969\ : IoInMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__967\ : IoSpan4Mux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__966\ : Span4Mux_s1_v
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__965\ : Sp12to4
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__964\ : Span12Mux_s8_v
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__963\ : Odrv12
    port map (
            O => \N__4499\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__962\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4493\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__960\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4487\,
            I => \N__4482\
        );

    \I__958\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4479\
        );

    \I__957\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4476\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__4482\,
            I => \N__4473\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4479\,
            I => \N__4468\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4476\,
            I => \N__4468\
        );

    \I__953\ : Sp12to4
    port map (
            O => \N__4473\,
            I => \N__4465\
        );

    \I__952\ : Span12Mux_v
    port map (
            O => \N__4468\,
            I => \N__4462\
        );

    \I__951\ : Span12Mux_v
    port map (
            O => \N__4465\,
            I => \N__4459\
        );

    \I__950\ : Span12Mux_h
    port map (
            O => \N__4462\,
            I => \N__4456\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__4459\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__948\ : Odrv12
    port map (
            O => \N__4456\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__947\ : IoInMux
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__945\ : Span4Mux_s3_h
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__944\ : Span4Mux_v
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__943\ : Sp12to4
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__942\ : Span12Mux_h
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__941\ : Odrv12
    port map (
            O => \N__4433\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__940\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__4424\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__937\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4416\
        );

    \I__936\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4413\
        );

    \I__935\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4410\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4407\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4402\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4402\
        );

    \I__931\ : Span4Mux_v
    port map (
            O => \N__4407\,
            I => \N__4397\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__4402\,
            I => \N__4397\
        );

    \I__929\ : Sp12to4
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__928\ : Span12Mux_h
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__927\ : Odrv12
    port map (
            O => \N__4391\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__926\ : IoInMux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__924\ : Span4Mux_s3_v
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__923\ : Span4Mux_h
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__4370\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__919\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__4361\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__916\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4354\
        );

    \I__915\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4351\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4354\,
            I => \N__4348\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4351\,
            I => \N__4345\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__4348\,
            I => \N__4342\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__910\ : Sp12to4
    port map (
            O => \N__4342\,
            I => \N__4335\
        );

    \I__909\ : Span4Mux_h
    port map (
            O => \N__4339\,
            I => \N__4332\
        );

    \I__908\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4329\
        );

    \I__907\ : Span12Mux_h
    port map (
            O => \N__4335\,
            I => \N__4326\
        );

    \I__906\ : Sp12to4
    port map (
            O => \N__4332\,
            I => \N__4321\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4329\,
            I => \N__4321\
        );

    \I__904\ : Span12Mux_v
    port map (
            O => \N__4326\,
            I => \N__4316\
        );

    \I__903\ : Span12Mux_h
    port map (
            O => \N__4321\,
            I => \N__4316\
        );

    \I__902\ : Odrv12
    port map (
            O => \N__4316\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__901\ : IoInMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__899\ : IoSpan4Mux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__898\ : Span4Mux_s3_v
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__896\ : Sp12to4
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__4295\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__894\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__4286\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__891\ : InMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4275\
        );

    \I__889\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4272\
        );

    \I__888\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4269\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__4275\,
            I => \N__4266\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4272\,
            I => \N__4261\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4269\,
            I => \N__4261\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__4266\,
            I => \N__4258\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__4261\,
            I => \N__4255\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__4255\,
            I => \N__4249\
        );

    \I__880\ : Sp12to4
    port map (
            O => \N__4252\,
            I => \N__4244\
        );

    \I__879\ : Sp12to4
    port map (
            O => \N__4249\,
            I => \N__4244\
        );

    \I__878\ : Span12Mux_h
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__4241\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__876\ : IoInMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__874\ : Span12Mux_s7_v
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__873\ : Span12Mux_h
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__872\ : Odrv12
    port map (
            O => \N__4226\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__871\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4216\
        );

    \I__869\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4213\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__4216\,
            I => \N__4209\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4206\
        );

    \I__866\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4203\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__4209\,
            I => \N__4200\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__4206\,
            I => \N__4197\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4203\,
            I => \N__4194\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__4200\,
            I => \N__4191\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__4197\,
            I => \N__4186\
        );

    \I__860\ : Span4Mux_v
    port map (
            O => \N__4194\,
            I => \N__4186\
        );

    \I__859\ : Span12Mux_h
    port map (
            O => \N__4191\,
            I => \N__4183\
        );

    \I__858\ : Sp12to4
    port map (
            O => \N__4186\,
            I => \N__4180\
        );

    \I__857\ : Span12Mux_v
    port map (
            O => \N__4183\,
            I => \N__4175\
        );

    \I__856\ : Span12Mux_h
    port map (
            O => \N__4180\,
            I => \N__4175\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__4175\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__854\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__4166\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__851\ : IoInMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__849\ : Span4Mux_s3_v
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__848\ : Span4Mux_h
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__846\ : Sp12to4
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__4145\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__844\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__4136\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__841\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4129\
        );

    \I__840\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4129\,
            I => \N__4122\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4119\
        );

    \I__837\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4116\
        );

    \I__836\ : Sp12to4
    port map (
            O => \N__4122\,
            I => \N__4109\
        );

    \I__835\ : Span12Mux_s9_v
    port map (
            O => \N__4119\,
            I => \N__4109\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4109\
        );

    \I__833\ : Span12Mux_h
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__832\ : Odrv12
    port map (
            O => \N__4106\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__831\ : IoInMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__829\ : Span12Mux_s6_v
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__828\ : Span12Mux_h
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__4091\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__826\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__824\ : Span12Mux_h
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__4079\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__822\ : IoInMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__820\ : IoSpan4Mux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__819\ : Span4Mux_s2_h
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__818\ : Sp12to4
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__817\ : Span12Mux_h
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__4058\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__815\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4051\
        );

    \I__814\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4048\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4051\,
            I => \N__4045\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4048\,
            I => \N__4041\
        );

    \I__811\ : Glb2LocalMux
    port map (
            O => \N__4045\,
            I => \N__4034\
        );

    \I__810\ : ClkMux
    port map (
            O => \N__4044\,
            I => \N__4034\
        );

    \I__809\ : Glb2LocalMux
    port map (
            O => \N__4041\,
            I => \N__4034\
        );

    \I__808\ : GlobalMux
    port map (
            O => \N__4034\,
            I => \CLK40\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__806\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__804\ : Span4Mux_h
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__4013\,
            I => \TS_CPUn_c\
        );

    \I__800\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4007\,
            I => \U111_CYCLE_SM.TS_EN_4\
        );

    \I__798\ : InMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__794\ : Span12Mux_h
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__793\ : Span12Mux_v
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__3986\,
            I => \PORTSIZE_c\
        );

    \I__791\ : IoInMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__789\ : Span4Mux_s2_v
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__788\ : Span4Mux_h
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__787\ : Sp12to4
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__786\ : Span12Mux_s9_v
    port map (
            O => \N__3968\,
            I => \N__3964\
        );

    \I__785\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3961\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__3964\,
            I => \TSn_c\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3961\,
            I => \TSn_c\
        );

    \I__782\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__780\ : Span4Mux_v
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__778\ : Span12Mux_h
    port map (
            O => \N__3944\,
            I => \N__3940\
        );

    \I__777\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3937\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__3940\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__3932\,
            I => \U111_CYCLE_SM.TS_EN10_cascade_\
        );

    \I__773\ : InMux
    port map (
            O => \N__3929\,
            I => \N__3925\
        );

    \I__772\ : InMux
    port map (
            O => \N__3928\,
            I => \N__3922\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3925\,
            I => \N__3919\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3922\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__3919\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__3914\,
            I => \N__3910\
        );

    \I__767\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3905\
        );

    \I__766\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3905\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3905\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__764\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3899\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__3896\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\
        );

    \I__761\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3890\,
            I => \U111_CYCLE_SM.LW_CYCLE_r_1\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3884\,
            I => \N__3881\
        );

    \I__757\ : IoSpan4Mux
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__756\ : Sp12to4
    port map (
            O => \N__3878\,
            I => \N__3875\
        );

    \I__755\ : Span12Mux_s6_v
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__3872\,
            I => \un1_D_UU_040_4\
        );

    \I__753\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__750\ : Sp12to4
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__749\ : Span12Mux_h
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__748\ : Odrv12
    port map (
            O => \N__3854\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__745\ : IoSpan4Mux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__744\ : IoSpan4Mux
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__743\ : Span4Mux_s2_h
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__742\ : Sp12to4
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__741\ : Span12Mux_s11_h
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__740\ : Odrv12
    port map (
            O => \N__3830\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__739\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3824\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__3821\,
            I => \N__3818\
        );

    \I__736\ : Sp12to4
    port map (
            O => \N__3818\,
            I => \N__3815\
        );

    \I__735\ : Span12Mux_h
    port map (
            O => \N__3815\,
            I => \N__3812\
        );

    \I__734\ : Odrv12
    port map (
            O => \N__3812\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__733\ : IoInMux
    port map (
            O => \N__3809\,
            I => \N__3806\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3806\,
            I => \N__3803\
        );

    \I__731\ : Span12Mux_s9_h
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__3800\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__729\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3794\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__727\ : Span12Mux_v
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__726\ : Span12Mux_h
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__3785\,
            I => \D_UU_040_in_2\
        );

    \I__724\ : InMux
    port map (
            O => \N__3782\,
            I => \N__3778\
        );

    \I__723\ : IoInMux
    port map (
            O => \N__3781\,
            I => \N__3775\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__3772\,
            I => \N__3766\
        );

    \I__719\ : Span12Mux_s5_h
    port map (
            O => \N__3769\,
            I => \N__3763\
        );

    \I__718\ : Sp12to4
    port map (
            O => \N__3766\,
            I => \N__3760\
        );

    \I__717\ : Span12Mux_v
    port map (
            O => \N__3763\,
            I => \N__3757\
        );

    \I__716\ : Span12Mux_v
    port map (
            O => \N__3760\,
            I => \N__3754\
        );

    \I__715\ : Span12Mux_h
    port map (
            O => \N__3757\,
            I => \N__3749\
        );

    \I__714\ : Span12Mux_v
    port map (
            O => \N__3754\,
            I => \N__3749\
        );

    \I__713\ : Span12Mux_h
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__712\ : Odrv12
    port map (
            O => \N__3746\,
            I => \D_LM_040_in_2\
        );

    \I__711\ : IoInMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__709\ : IoSpan4Mux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__708\ : IoSpan4Mux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__707\ : Span4Mux_s2_v
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__3725\,
            I => \un1_D_UU_040_2\
        );

    \I__704\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__701\ : Sp12to4
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__700\ : Span12Mux_h
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__3707\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__698\ : IoInMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__696\ : Span12Mux_s4_h
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__695\ : Span12Mux_h
    port map (
            O => \N__3695\,
            I => \N__3692\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__3692\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__693\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__689\ : Span12Mux_h
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__3674\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__687\ : IoInMux
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__685\ : IoSpan4Mux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__684\ : IoSpan4Mux
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__683\ : Span4Mux_s3_h
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__682\ : Sp12to4
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__681\ : Odrv12
    port map (
            O => \N__3653\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__680\ : IoInMux
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3647\,
            I => \N__3643\
        );

    \I__678\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3640\
        );

    \I__677\ : IoSpan4Mux
    port map (
            O => \N__3643\,
            I => \N__3637\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3640\,
            I => \N__3634\
        );

    \I__675\ : Span4Mux_s2_h
    port map (
            O => \N__3637\,
            I => \N__3631\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__3634\,
            I => \N__3628\
        );

    \I__673\ : Sp12to4
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__672\ : Sp12to4
    port map (
            O => \N__3628\,
            I => \N__3622\
        );

    \I__671\ : Span12Mux_h
    port map (
            O => \N__3625\,
            I => \N__3619\
        );

    \I__670\ : Span12Mux_h
    port map (
            O => \N__3622\,
            I => \N__3616\
        );

    \I__669\ : Span12Mux_h
    port map (
            O => \N__3619\,
            I => \N__3613\
        );

    \I__668\ : Span12Mux_v
    port map (
            O => \N__3616\,
            I => \N__3610\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__3613\,
            I => \D_LL_040_in_2\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__3610\,
            I => \D_LL_040_in_2\
        );

    \I__665\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__663\ : Span12Mux_h
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__3596\,
            I => \D_UM_040_in_2\
        );

    \I__661\ : IoInMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__659\ : Span4Mux_s2_h
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__657\ : Sp12to4
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__655\ : Odrv12
    port map (
            O => \N__3575\,
            I => \un1_D_UM_040_2\
        );

    \I__654\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__652\ : Glb2LocalMux
    port map (
            O => \N__3566\,
            I => \N__3542\
        );

    \I__651\ : ClkMux
    port map (
            O => \N__3565\,
            I => \N__3542\
        );

    \I__650\ : ClkMux
    port map (
            O => \N__3564\,
            I => \N__3542\
        );

    \I__649\ : ClkMux
    port map (
            O => \N__3563\,
            I => \N__3542\
        );

    \I__648\ : ClkMux
    port map (
            O => \N__3562\,
            I => \N__3542\
        );

    \I__647\ : ClkMux
    port map (
            O => \N__3561\,
            I => \N__3542\
        );

    \I__646\ : ClkMux
    port map (
            O => \N__3560\,
            I => \N__3542\
        );

    \I__645\ : ClkMux
    port map (
            O => \N__3559\,
            I => \N__3542\
        );

    \I__644\ : GlobalMux
    port map (
            O => \N__3542\,
            I => \CLK80\
        );

    \I__643\ : IoInMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3536\,
            I => \N__3533\
        );

    \I__641\ : IoSpan4Mux
    port map (
            O => \N__3533\,
            I => \N__3529\
        );

    \I__640\ : IoInMux
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__639\ : IoSpan4Mux
    port map (
            O => \N__3529\,
            I => \N__3521\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3526\,
            I => \N__3521\
        );

    \I__637\ : Span4Mux_s2_v
    port map (
            O => \N__3521\,
            I => \N__3517\
        );

    \I__636\ : IoInMux
    port map (
            O => \N__3520\,
            I => \N__3514\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__3517\,
            I => \N__3511\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3514\,
            I => \N__3508\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__3511\,
            I => \N__3505\
        );

    \I__632\ : Span12Mux_s4_h
    port map (
            O => \N__3508\,
            I => \N__3502\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__3505\,
            I => \N__3499\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__3502\,
            I => \N__3496\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__3499\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3496\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__627\ : IoInMux
    port map (
            O => \N__3491\,
            I => \N__3487\
        );

    \I__626\ : IoInMux
    port map (
            O => \N__3490\,
            I => \N__3484\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3481\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3478\
        );

    \I__623\ : Span4Mux_s3_h
    port map (
            O => \N__3481\,
            I => \N__3475\
        );

    \I__622\ : Span4Mux_s3_h
    port map (
            O => \N__3478\,
            I => \N__3472\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__3475\,
            I => \N__3468\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__3472\,
            I => \N__3465\
        );

    \I__619\ : IoInMux
    port map (
            O => \N__3471\,
            I => \N__3462\
        );

    \I__618\ : Sp12to4
    port map (
            O => \N__3468\,
            I => \N__3459\
        );

    \I__617\ : Span12Mux_v
    port map (
            O => \N__3465\,
            I => \N__3456\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3462\,
            I => \N__3453\
        );

    \I__615\ : Span12Mux_h
    port map (
            O => \N__3459\,
            I => \N__3446\
        );

    \I__614\ : Span12Mux_h
    port map (
            O => \N__3456\,
            I => \N__3446\
        );

    \I__613\ : Span12Mux_s11_v
    port map (
            O => \N__3453\,
            I => \N__3446\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__3446\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__611\ : IoInMux
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__609\ : Span12Mux_s10_h
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__608\ : Span12Mux_v
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__3431\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__606\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__603\ : Sp12to4
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__602\ : Span12Mux_h
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__3413\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__600\ : IoInMux
    port map (
            O => \N__3410\,
            I => \N__3407\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3407\,
            I => \N__3404\
        );

    \I__598\ : Span12Mux_s7_h
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__597\ : Span12Mux_h
    port map (
            O => \N__3401\,
            I => \N__3398\
        );

    \I__596\ : Odrv12
    port map (
            O => \N__3398\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__595\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3391\
        );

    \I__594\ : IoInMux
    port map (
            O => \N__3394\,
            I => \N__3388\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3391\,
            I => \N__3385\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3388\,
            I => \N__3382\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__3385\,
            I => \N__3379\
        );

    \I__590\ : Span4Mux_s3_h
    port map (
            O => \N__3382\,
            I => \N__3376\
        );

    \I__589\ : Sp12to4
    port map (
            O => \N__3379\,
            I => \N__3373\
        );

    \I__588\ : Sp12to4
    port map (
            O => \N__3376\,
            I => \N__3370\
        );

    \I__587\ : Span12Mux_h
    port map (
            O => \N__3373\,
            I => \N__3367\
        );

    \I__586\ : Span12Mux_v
    port map (
            O => \N__3370\,
            I => \N__3364\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__3367\,
            I => \N__3361\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__3364\,
            I => \N__3358\
        );

    \I__583\ : Span12Mux_v
    port map (
            O => \N__3361\,
            I => \N__3355\
        );

    \I__582\ : Span12Mux_h
    port map (
            O => \N__3358\,
            I => \N__3352\
        );

    \I__581\ : Odrv12
    port map (
            O => \N__3355\,
            I => \D_LL_040_in_3\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__3352\,
            I => \D_LL_040_in_3\
        );

    \I__579\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3344\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3344\,
            I => \N__3341\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__3341\,
            I => \N__3338\
        );

    \I__576\ : Span12Mux_v
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__3335\,
            I => \N__3332\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__3332\,
            I => \D_UM_040_in_3\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__571\ : IoSpan4Mux
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__570\ : Sp12to4
    port map (
            O => \N__3320\,
            I => \N__3317\
        );

    \I__569\ : Span12Mux_s6_h
    port map (
            O => \N__3317\,
            I => \N__3314\
        );

    \I__568\ : Odrv12
    port map (
            O => \N__3314\,
            I => \un1_D_UM_040_3\
        );

    \I__567\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__564\ : Span4Mux_h
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__563\ : Sp12to4
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__562\ : Span12Mux_h
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__3293\,
            I => \D_UM_040_in_4\
        );

    \I__560\ : IoInMux
    port map (
            O => \N__3290\,
            I => \N__3286\
        );

    \I__559\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3283\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3286\,
            I => \N__3280\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3283\,
            I => \N__3277\
        );

    \I__556\ : Span4Mux_s2_h
    port map (
            O => \N__3280\,
            I => \N__3274\
        );

    \I__555\ : Sp12to4
    port map (
            O => \N__3277\,
            I => \N__3271\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__3274\,
            I => \N__3268\
        );

    \I__553\ : Span12Mux_v
    port map (
            O => \N__3271\,
            I => \N__3265\
        );

    \I__552\ : Sp12to4
    port map (
            O => \N__3268\,
            I => \N__3262\
        );

    \I__551\ : Span12Mux_v
    port map (
            O => \N__3265\,
            I => \N__3257\
        );

    \I__550\ : Span12Mux_h
    port map (
            O => \N__3262\,
            I => \N__3257\
        );

    \I__549\ : Span12Mux_h
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__548\ : Odrv12
    port map (
            O => \N__3254\,
            I => \D_LL_040_in_4\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__545\ : IoSpan4Mux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__544\ : Sp12to4
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__543\ : Span12Mux_h
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__3236\,
            I => \un1_D_UM_040_4\
        );

    \I__541\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__536\ : Span12Mux_h
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__535\ : Odrv12
    port map (
            O => \N__3215\,
            I => \D_UU_040_in_7\
        );

    \I__534\ : IoInMux
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__532\ : IoSpan4Mux
    port map (
            O => \N__3206\,
            I => \N__3202\
        );

    \I__531\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3199\
        );

    \I__530\ : Span4Mux_s2_h
    port map (
            O => \N__3202\,
            I => \N__3196\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__3196\,
            I => \N__3190\
        );

    \I__527\ : Sp12to4
    port map (
            O => \N__3193\,
            I => \N__3187\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__3190\,
            I => \N__3182\
        );

    \I__525\ : Span12Mux_s9_v
    port map (
            O => \N__3187\,
            I => \N__3182\
        );

    \I__524\ : Span12Mux_h
    port map (
            O => \N__3182\,
            I => \N__3179\
        );

    \I__523\ : Odrv12
    port map (
            O => \N__3179\,
            I => \D_LM_040_in_7\
        );

    \I__522\ : IoInMux
    port map (
            O => \N__3176\,
            I => \N__3173\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__520\ : IoSpan4Mux
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__519\ : Sp12to4
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__518\ : Span12Mux_s6_v
    port map (
            O => \N__3164\,
            I => \N__3161\
        );

    \I__517\ : Odrv12
    port map (
            O => \N__3161\,
            I => \un1_D_UU_040_7\
        );

    \I__516\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__514\ : Span12Mux_v
    port map (
            O => \N__3152\,
            I => \N__3149\
        );

    \I__513\ : Span12Mux_h
    port map (
            O => \N__3149\,
            I => \N__3146\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__3146\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__511\ : IoInMux
    port map (
            O => \N__3143\,
            I => \N__3140\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3140\,
            I => \N__3137\
        );

    \I__509\ : Span4Mux_s3_h
    port map (
            O => \N__3137\,
            I => \N__3134\
        );

    \I__508\ : Span4Mux_v
    port map (
            O => \N__3134\,
            I => \N__3131\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3131\,
            I => \N__3128\
        );

    \I__506\ : Sp12to4
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__505\ : Span12Mux_s11_h
    port map (
            O => \N__3125\,
            I => \N__3122\
        );

    \I__504\ : Odrv12
    port map (
            O => \N__3122\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__503\ : IoInMux
    port map (
            O => \N__3119\,
            I => \N__3116\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__501\ : IoSpan4Mux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__500\ : IoSpan4Mux
    port map (
            O => \N__3110\,
            I => \N__3106\
        );

    \I__499\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3103\
        );

    \I__498\ : Span4Mux_s2_h
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__496\ : Sp12to4
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__495\ : Span12Mux_v
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__494\ : Span12Mux_h
    port map (
            O => \N__3094\,
            I => \N__3086\
        );

    \I__493\ : Span12Mux_v
    port map (
            O => \N__3091\,
            I => \N__3086\
        );

    \I__492\ : Span12Mux_h
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__3083\,
            I => \D_LL_040_in_6\
        );

    \I__490\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__488\ : Span12Mux_v
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__487\ : Span12Mux_h
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__3068\,
            I => \D_UM_040_in_6\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__483\ : Span12Mux_s10_h
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__482\ : Span12Mux_v
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__481\ : Odrv12
    port map (
            O => \N__3053\,
            I => \un1_D_UM_040_6\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3043\
        );

    \I__478\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3040\
        );

    \I__477\ : IoSpan4Mux
    port map (
            O => \N__3043\,
            I => \N__3037\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3040\,
            I => \N__3034\
        );

    \I__475\ : Span4Mux_s3_h
    port map (
            O => \N__3037\,
            I => \N__3031\
        );

    \I__474\ : Span4Mux_h
    port map (
            O => \N__3034\,
            I => \N__3028\
        );

    \I__473\ : Sp12to4
    port map (
            O => \N__3031\,
            I => \N__3025\
        );

    \I__472\ : Sp12to4
    port map (
            O => \N__3028\,
            I => \N__3022\
        );

    \I__471\ : Span12Mux_v
    port map (
            O => \N__3025\,
            I => \N__3019\
        );

    \I__470\ : Span12Mux_v
    port map (
            O => \N__3022\,
            I => \N__3016\
        );

    \I__469\ : Span12Mux_h
    port map (
            O => \N__3019\,
            I => \N__3011\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__3016\,
            I => \N__3011\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__3008\,
            I => \D_LL_040_in_7\
        );

    \I__465\ : InMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__461\ : Sp12to4
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__460\ : Span12Mux_h
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__459\ : Odrv12
    port map (
            O => \N__2987\,
            I => \D_UM_040_in_7\
        );

    \I__458\ : IoInMux
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__456\ : Span4Mux_s1_h
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__455\ : Span4Mux_h
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__454\ : Span4Mux_h
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__453\ : Span4Mux_h
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__2966\,
            I => \un1_D_UM_040_7\
        );

    \I__451\ : IoInMux
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__449\ : Span4Mux_s1_h
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__448\ : Sp12to4
    port map (
            O => \N__2954\,
            I => \N__2950\
        );

    \I__447\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2947\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__2950\,
            I => \N__2944\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__444\ : Span12Mux_h
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__443\ : Span12Mux_h
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__442\ : Span12Mux_h
    port map (
            O => \N__2938\,
            I => \N__2930\
        );

    \I__441\ : Span12Mux_v
    port map (
            O => \N__2935\,
            I => \N__2930\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__2930\,
            I => \D_LM_040_in_4\
        );

    \I__439\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__436\ : Span12Mux_h
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__2915\,
            I => \D_UU_040_in_4\
        );

    \I__434\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__432\ : Span4Mux_v
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__431\ : Sp12to4
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__2900\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__429\ : IoInMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__427\ : Span4Mux_s1_h
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__426\ : Sp12to4
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__425\ : Span12Mux_v
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__424\ : Span12Mux_h
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__2879\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__422\ : IoInMux
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2873\,
            I => \N__2870\
        );

    \I__420\ : IoSpan4Mux
    port map (
            O => \N__2870\,
            I => \N__2866\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__2869\,
            I => \N__2863\
        );

    \I__418\ : IoSpan4Mux
    port map (
            O => \N__2866\,
            I => \N__2860\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2863\,
            I => \N__2857\
        );

    \I__416\ : IoSpan4Mux
    port map (
            O => \N__2860\,
            I => \N__2852\
        );

    \I__415\ : IoSpan4Mux
    port map (
            O => \N__2857\,
            I => \N__2852\
        );

    \I__414\ : Span4Mux_s3_v
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__413\ : Odrv4
    port map (
            O => \N__2849\,
            I => \CONSTANT_ONE_NET\
        );

    \I__412\ : InMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__410\ : Span4Mux_v
    port map (
            O => \N__2840\,
            I => \N__2837\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__408\ : Sp12to4
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__407\ : Span12Mux_h
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__406\ : Odrv12
    port map (
            O => \N__2828\,
            I => \D_UU_040_in_0\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__2825\,
            I => \N__2821\
        );

    \I__404\ : InMux
    port map (
            O => \N__2824\,
            I => \N__2818\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2821\,
            I => \N__2815\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2818\,
            I => \N__2812\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__2815\,
            I => \N__2809\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__2812\,
            I => \N__2806\
        );

    \I__399\ : IoSpan4Mux
    port map (
            O => \N__2809\,
            I => \N__2803\
        );

    \I__398\ : Sp12to4
    port map (
            O => \N__2806\,
            I => \N__2800\
        );

    \I__397\ : Span4Mux_s2_h
    port map (
            O => \N__2803\,
            I => \N__2797\
        );

    \I__396\ : Span12Mux_h
    port map (
            O => \N__2800\,
            I => \N__2794\
        );

    \I__395\ : Sp12to4
    port map (
            O => \N__2797\,
            I => \N__2791\
        );

    \I__394\ : Span12Mux_v
    port map (
            O => \N__2794\,
            I => \N__2788\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__2791\,
            I => \N__2785\
        );

    \I__392\ : Span12Mux_v
    port map (
            O => \N__2788\,
            I => \N__2782\
        );

    \I__391\ : Span12Mux_h
    port map (
            O => \N__2785\,
            I => \N__2779\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__2782\,
            I => \D_LM_040_in_0\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__2779\,
            I => \D_LM_040_in_0\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2771\,
            I => \N__2768\
        );

    \I__386\ : IoSpan4Mux
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__385\ : Span4Mux_s2_v
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__384\ : Span4Mux_v
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2759\,
            I => \un1_D_UU_040_0\
        );

    \I__382\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2753\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__380\ : Span4Mux_v
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__379\ : Sp12to4
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__378\ : Span12Mux_h
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__2741\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2735\,
            I => \N__2732\
        );

    \I__374\ : Span4Mux_s3_h
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__373\ : Sp12to4
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__372\ : Span12Mux_s8_v
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__371\ : Span12Mux_h
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__2720\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__369\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__366\ : Sp12to4
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__365\ : Span12Mux_h
    port map (
            O => \N__2705\,
            I => \N__2702\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__2702\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__363\ : IoInMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__361\ : Span4Mux_s3_h
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__359\ : Span4Mux_v
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__358\ : Sp12to4
    port map (
            O => \N__2684\,
            I => \N__2681\
        );

    \I__357\ : Span12Mux_h
    port map (
            O => \N__2681\,
            I => \N__2678\
        );

    \I__356\ : Odrv12
    port map (
            O => \N__2678\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__355\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2672\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2672\,
            I => \N__2669\
        );

    \I__353\ : Span12Mux_v
    port map (
            O => \N__2669\,
            I => \N__2666\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__2666\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__351\ : IoInMux
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__349\ : Span4Mux_s1_h
    port map (
            O => \N__2657\,
            I => \N__2654\
        );

    \I__348\ : Sp12to4
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__347\ : Span12Mux_v
    port map (
            O => \N__2651\,
            I => \N__2648\
        );

    \I__346\ : Span12Mux_h
    port map (
            O => \N__2648\,
            I => \N__2645\
        );

    \I__345\ : Odrv12
    port map (
            O => \N__2645\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__2642\,
            I => \N__2639\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2639\,
            I => \N__2635\
        );

    \I__342\ : InMux
    port map (
            O => \N__2638\,
            I => \N__2632\
        );

    \I__341\ : Span4Mux_s2_h
    port map (
            O => \N__2635\,
            I => \N__2629\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2632\,
            I => \N__2626\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__2629\,
            I => \N__2623\
        );

    \I__338\ : Span4Mux_v
    port map (
            O => \N__2626\,
            I => \N__2620\
        );

    \I__337\ : Sp12to4
    port map (
            O => \N__2623\,
            I => \N__2617\
        );

    \I__336\ : Span4Mux_v
    port map (
            O => \N__2620\,
            I => \N__2614\
        );

    \I__335\ : Span12Mux_h
    port map (
            O => \N__2617\,
            I => \N__2609\
        );

    \I__334\ : Sp12to4
    port map (
            O => \N__2614\,
            I => \N__2609\
        );

    \I__333\ : Span12Mux_h
    port map (
            O => \N__2609\,
            I => \N__2606\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__2606\,
            I => \D_LM_040_in_6\
        );

    \I__331\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2600\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2600\,
            I => \N__2597\
        );

    \I__329\ : Span4Mux_v
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__328\ : Span4Mux_h
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__327\ : Sp12to4
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__326\ : Span12Mux_h
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__325\ : Odrv12
    port map (
            O => \N__2585\,
            I => \D_UU_040_in_6\
        );

    \I__324\ : IoInMux
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__322\ : IoSpan4Mux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__321\ : IoSpan4Mux
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__320\ : Span4Mux_s3_v
    port map (
            O => \N__2570\,
            I => \N__2567\
        );

    \I__319\ : Odrv4
    port map (
            O => \N__2567\,
            I => \un1_D_UU_040_6\
        );

    \I__318\ : InMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__316\ : Span4Mux_v
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__315\ : Sp12to4
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__314\ : Odrv12
    port map (
            O => \N__2552\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__313\ : IoInMux
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__311\ : Span4Mux_s0_h
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__310\ : Sp12to4
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__309\ : Span12Mux_s8_v
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__308\ : Span12Mux_h
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__307\ : Odrv12
    port map (
            O => \N__2531\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__306\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__304\ : Span12Mux_h
    port map (
            O => \N__2522\,
            I => \N__2519\
        );

    \I__303\ : Odrv12
    port map (
            O => \N__2519\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__302\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2513\,
            I => \N__2510\
        );

    \I__300\ : Span12Mux_h
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__299\ : Odrv12
    port map (
            O => \N__2507\,
            I => \A_040_c_1\
        );

    \I__298\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2501\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2501\,
            I => \N__2498\
        );

    \I__296\ : Span4Mux_h
    port map (
            O => \N__2498\,
            I => \N__2495\
        );

    \I__295\ : Span4Mux_v
    port map (
            O => \N__2495\,
            I => \N__2492\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2492\,
            I => \A_040_c_0\
        );

    \I__293\ : IoInMux
    port map (
            O => \N__2489\,
            I => \N__2486\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2486\,
            I => \N__2483\
        );

    \I__291\ : Span4Mux_s2_v
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__290\ : Span4Mux_v
    port map (
            O => \N__2480\,
            I => \N__2477\
        );

    \I__289\ : Odrv4
    port map (
            O => \N__2477\,
            I => \A_AMIGA_c_0\
        );

    \I__288\ : IoInMux
    port map (
            O => \N__2474\,
            I => \N__2467\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2473\,
            I => \N__2464\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2472\,
            I => \N__2459\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2471\,
            I => \N__2456\
        );

    \I__284\ : IoInMux
    port map (
            O => \N__2470\,
            I => \N__2453\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2467\,
            I => \N__2444\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2464\,
            I => \N__2444\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__2463\,
            I => \N__2441\
        );

    \I__280\ : IoInMux
    port map (
            O => \N__2462\,
            I => \N__2438\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2459\,
            I => \N__2427\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2456\,
            I => \N__2427\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2453\,
            I => \N__2427\
        );

    \I__276\ : IoInMux
    port map (
            O => \N__2452\,
            I => \N__2424\
        );

    \I__275\ : IoInMux
    port map (
            O => \N__2451\,
            I => \N__2421\
        );

    \I__274\ : IoInMux
    port map (
            O => \N__2450\,
            I => \N__2418\
        );

    \I__273\ : IoInMux
    port map (
            O => \N__2449\,
            I => \N__2415\
        );

    \I__272\ : IoSpan4Mux
    port map (
            O => \N__2444\,
            I => \N__2399\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2441\,
            I => \N__2399\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2438\,
            I => \N__2399\
        );

    \I__269\ : IoInMux
    port map (
            O => \N__2437\,
            I => \N__2396\
        );

    \I__268\ : IoInMux
    port map (
            O => \N__2436\,
            I => \N__2393\
        );

    \I__267\ : IoInMux
    port map (
            O => \N__2435\,
            I => \N__2390\
        );

    \I__266\ : IoInMux
    port map (
            O => \N__2434\,
            I => \N__2387\
        );

    \I__265\ : IoSpan4Mux
    port map (
            O => \N__2427\,
            I => \N__2376\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2424\,
            I => \N__2376\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2421\,
            I => \N__2376\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2418\,
            I => \N__2376\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2415\,
            I => \N__2376\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__2414\,
            I => \N__2373\
        );

    \I__259\ : IoInMux
    port map (
            O => \N__2413\,
            I => \N__2370\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2412\,
            I => \N__2367\
        );

    \I__257\ : IoInMux
    port map (
            O => \N__2411\,
            I => \N__2364\
        );

    \I__256\ : IoInMux
    port map (
            O => \N__2410\,
            I => \N__2357\
        );

    \I__255\ : IoInMux
    port map (
            O => \N__2409\,
            I => \N__2354\
        );

    \I__254\ : IoInMux
    port map (
            O => \N__2408\,
            I => \N__2351\
        );

    \I__253\ : IoInMux
    port map (
            O => \N__2407\,
            I => \N__2348\
        );

    \I__252\ : IoInMux
    port map (
            O => \N__2406\,
            I => \N__2345\
        );

    \I__251\ : IoSpan4Mux
    port map (
            O => \N__2399\,
            I => \N__2334\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2396\,
            I => \N__2334\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2393\,
            I => \N__2334\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2390\,
            I => \N__2334\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2387\,
            I => \N__2334\
        );

    \I__246\ : IoSpan4Mux
    port map (
            O => \N__2376\,
            I => \N__2323\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2373\,
            I => \N__2323\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2370\,
            I => \N__2323\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2367\,
            I => \N__2323\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2364\,
            I => \N__2323\
        );

    \I__241\ : IoInMux
    port map (
            O => \N__2363\,
            I => \N__2320\
        );

    \I__240\ : IoInMux
    port map (
            O => \N__2362\,
            I => \N__2317\
        );

    \I__239\ : IoInMux
    port map (
            O => \N__2361\,
            I => \N__2314\
        );

    \I__238\ : IoInMux
    port map (
            O => \N__2360\,
            I => \N__2311\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2357\,
            I => \N__2298\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2354\,
            I => \N__2298\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2351\,
            I => \N__2298\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2348\,
            I => \N__2298\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2345\,
            I => \N__2298\
        );

    \I__232\ : IoSpan4Mux
    port map (
            O => \N__2334\,
            I => \N__2294\
        );

    \I__231\ : IoSpan4Mux
    port map (
            O => \N__2323\,
            I => \N__2283\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2320\,
            I => \N__2283\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2317\,
            I => \N__2283\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2314\,
            I => \N__2283\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2311\,
            I => \N__2283\
        );

    \I__226\ : IoInMux
    port map (
            O => \N__2310\,
            I => \N__2280\
        );

    \I__225\ : IoInMux
    port map (
            O => \N__2309\,
            I => \N__2277\
        );

    \I__224\ : IoSpan4Mux
    port map (
            O => \N__2298\,
            I => \N__2274\
        );

    \I__223\ : IoInMux
    port map (
            O => \N__2297\,
            I => \N__2271\
        );

    \I__222\ : IoSpan4Mux
    port map (
            O => \N__2294\,
            I => \N__2266\
        );

    \I__221\ : IoSpan4Mux
    port map (
            O => \N__2283\,
            I => \N__2266\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2263\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2277\,
            I => \N__2260\
        );

    \I__218\ : Span4Mux_s3_v
    port map (
            O => \N__2274\,
            I => \N__2257\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2271\,
            I => \N__2254\
        );

    \I__216\ : Span4Mux_s1_h
    port map (
            O => \N__2266\,
            I => \N__2251\
        );

    \I__215\ : Span4Mux_s1_h
    port map (
            O => \N__2263\,
            I => \N__2248\
        );

    \I__214\ : Span12Mux_s6_h
    port map (
            O => \N__2260\,
            I => \N__2244\
        );

    \I__213\ : Sp12to4
    port map (
            O => \N__2257\,
            I => \N__2239\
        );

    \I__212\ : Span12Mux_s4_v
    port map (
            O => \N__2254\,
            I => \N__2239\
        );

    \I__211\ : Span4Mux_h
    port map (
            O => \N__2251\,
            I => \N__2234\
        );

    \I__210\ : Span4Mux_h
    port map (
            O => \N__2248\,
            I => \N__2234\
        );

    \I__209\ : IoInMux
    port map (
            O => \N__2247\,
            I => \N__2231\
        );

    \I__208\ : Span12Mux_v
    port map (
            O => \N__2244\,
            I => \N__2226\
        );

    \I__207\ : Span12Mux_v
    port map (
            O => \N__2239\,
            I => \N__2226\
        );

    \I__206\ : Span4Mux_h
    port map (
            O => \N__2234\,
            I => \N__2223\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2231\,
            I => \N__2220\
        );

    \I__204\ : Odrv12
    port map (
            O => \N__2226\,
            I => \RnW_c_i_0\
        );

    \I__203\ : Odrv4
    port map (
            O => \N__2223\,
            I => \RnW_c_i_0\
        );

    \I__202\ : Odrv12
    port map (
            O => \N__2220\,
            I => \RnW_c_i_0\
        );

    \I__201\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2210\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2210\,
            I => \N__2207\
        );

    \I__199\ : Span4Mux_v
    port map (
            O => \N__2207\,
            I => \N__2204\
        );

    \I__198\ : Sp12to4
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__197\ : Odrv12
    port map (
            O => \N__2201\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__196\ : IoInMux
    port map (
            O => \N__2198\,
            I => \N__2195\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__2195\,
            I => \N__2192\
        );

    \I__194\ : IoSpan4Mux
    port map (
            O => \N__2192\,
            I => \N__2189\
        );

    \I__193\ : Sp12to4
    port map (
            O => \N__2189\,
            I => \N__2186\
        );

    \I__192\ : Span12Mux_s7_v
    port map (
            O => \N__2186\,
            I => \N__2183\
        );

    \I__191\ : Span12Mux_h
    port map (
            O => \N__2183\,
            I => \N__2180\
        );

    \I__190\ : Odrv12
    port map (
            O => \N__2180\,
            I => \un1_D_LL_AMIGA_3\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            I => \N__3562\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            I => \N__3565\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_1C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            I => \N__3561\
        );

    \INVU111_CYCLE_SM.TA_EN_nessC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            I => \N__3564\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            I => \N__3559\
        );

    \INVU111_CYCLE_SM.A_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.A_OUTC_net\,
            I => \N__3560\
        );

    \INVU111_CYCLE_SM.LW_CYCLE_STARTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            I => \N__3563\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__4044\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__2516\,
            in2 => \_gnd_net_\,
            in3 => \N__3956\,
            lcout => \A_AMIGA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6371\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RnW_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBVV92_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__6878\,
            in2 => \_gnd_net_\,
            in3 => \N__2213\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJ70A2_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2912\,
            in1 => \N__6870\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOVRM1_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2846\,
            in1 => \N__6849\,
            in2 => \_gnd_net_\,
            in3 => \N__2824\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7RV92_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2756\,
            in1 => \N__6877\,
            in2 => \_gnd_net_\,
            in3 => \N__4625\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIF30A2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4358\,
            in1 => \N__6869\,
            in2 => \_gnd_net_\,
            in3 => \N__2717\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIM8L62_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4553\,
            in1 => \N__6832\,
            in2 => \_gnd_net_\,
            in3 => \N__2675\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI4CSM1_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2638\,
            in1 => \N__6828\,
            in2 => \_gnd_net_\,
            in3 => \N__2603\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNID10A2_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2564\,
            in1 => \N__6848\,
            in2 => \_gnd_net_\,
            in3 => \N__4223\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNII4L62_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4421\,
            in1 => \N__6840\,
            in2 => \_gnd_net_\,
            in3 => \N__2528\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQCL62_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6824\,
            in1 => \N__4125\,
            in2 => \_gnd_net_\,
            in3 => \N__3428\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILGQ22_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3395\,
            in1 => \N__6825\,
            in2 => \_gnd_net_\,
            in3 => \N__3347\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINIQ22_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6826\,
            in1 => \N__3311\,
            in2 => \_gnd_net_\,
            in3 => \N__3289\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI6ESM1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3233\,
            in1 => \N__6827\,
            in2 => \_gnd_net_\,
            in3 => \N__3205\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIE0L62_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6413\,
            in1 => \N__6818\,
            in2 => \_gnd_net_\,
            in3 => \N__3158\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRMQ22_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3109\,
            in1 => \N__6839\,
            in2 => \_gnd_net_\,
            in3 => \N__3080\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITOQ22_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3046\,
            in1 => \N__6816\,
            in2 => \_gnd_net_\,
            in3 => \N__3005\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI08SM1_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2953\,
            in1 => \N__6817\,
            in2 => \_gnd_net_\,
            in3 => \N__2927\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOAL62_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6797\,
            in1 => \N__4283\,
            in2 => \_gnd_net_\,
            in3 => \N__3869\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISEL62_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3827\,
            in1 => \N__6813\,
            in2 => \_gnd_net_\,
            in3 => \N__6540\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIS3SM1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3797\,
            in1 => \N__3782\,
            in2 => \_gnd_net_\,
            in3 => \N__6814\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5PV92_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__6868\,
            in2 => \_gnd_net_\,
            in3 => \N__5261\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9TV92_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3689\,
            in1 => \N__6867\,
            in2 => \_gnd_net_\,
            in3 => \N__5312\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJEQ22_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3646\,
            in1 => \N__6833\,
            in2 => \_gnd_net_\,
            in3 => \N__3605\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3572\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4055\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4683\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3929\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6083\,
            in1 => \N__4004\,
            in2 => \N__4705\,
            in3 => \N__3967\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__5105\,
            in1 => \N__3943\,
            in2 => \N__4719\,
            in3 => \N__3902\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000100010"
        )
    port map (
            in0 => \N__3913\,
            in1 => \N__5061\,
            in2 => \N__5161\,
            in3 => \N__5103\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.TS_EN10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__4710\,
            in1 => \N__4010\,
            in2 => \N__3932\,
            in3 => \N__3928\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__6270\,
            in1 => \N__5060\,
            in2 => \N__3914\,
            in3 => \N__5102\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\,
            ltout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNO_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3896\,
            in3 => \N__5179\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__6271\,
            in1 => \N__3893\,
            in2 => \N__5111\,
            in3 => \N__4709\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__4054\,
            in1 => \N__5063\,
            in2 => \N__4031\,
            in3 => \N__5106\,
            lcout => \U111_CYCLE_SM.TS_EN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4420\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4486\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4279\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4549\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4219\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4620\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4133\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__5778\,
            sr => \N__5742\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4559\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \N__6312\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__4496\,
            in2 => \_gnd_net_\,
            in3 => \N__4485\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6341\,
            in1 => \N__4430\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6340\,
            in1 => \N__4367\,
            in2 => \_gnd_net_\,
            in3 => \N__4338\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6342\,
            in1 => \N__4292\,
            in2 => \_gnd_net_\,
            in3 => \N__4278\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4212\,
            in1 => \N__4172\,
            in2 => \_gnd_net_\,
            in3 => \N__6339\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4142\,
            in1 => \N__4132\,
            in2 => \_gnd_net_\,
            in3 => \N__6343\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIK6L62_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4088\,
            in1 => \N__6815\,
            in2 => \_gnd_net_\,
            in3 => \N__6485\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5201\,
            in2 => \_gnd_net_\,
            in3 => \N__5162\,
            lcout => \TAn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4711\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5110\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            ce => \N__5195\,
            sr => \N__5183\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5030\,
            in2 => \_gnd_net_\,
            in3 => \N__5723\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000001000000"
        )
    port map (
            in0 => \N__5164\,
            in1 => \N__5059\,
            in2 => \N__4721\,
            in3 => \N__5101\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__5163\,
            in1 => \N__5058\,
            in2 => \N__4720\,
            in3 => \N__5100\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5165\,
            in1 => \N__5099\,
            in2 => \_gnd_net_\,
            in3 => \N__5057\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__4958\,
            in1 => \_gnd_net_\,
            in2 => \N__4724\,
            in3 => \N__4718\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6338\,
            in1 => \N__4631\,
            in2 => \_gnd_net_\,
            in3 => \N__4621\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI2ASM1_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5554\,
            in1 => \N__6772\,
            in2 => \_gnd_net_\,
            in3 => \N__5519\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIH50A2_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5480\,
            in1 => \N__5360\,
            in2 => \_gnd_net_\,
            in3 => \N__6750\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIG2L62_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6749\,
            in1 => \N__5624\,
            in2 => \_gnd_net_\,
            in3 => \N__5441\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6357\,
            in1 => \N__5819\,
            in2 => \_gnd_net_\,
            in3 => \N__5244\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5356\,
            in1 => \N__5321\,
            in2 => \_gnd_net_\,
            in3 => \N__6356\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6355\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__5295\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5783\,
            sr => \N__5747\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5302\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5783\,
            sr => \N__5747\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5257\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5783\,
            sr => \N__5747\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIHM0E1_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000000000"
        )
    port map (
            in0 => \N__6347\,
            in1 => \N__6110\,
            in2 => \N__6143\,
            in3 => \N__5810\,
            lcout => \U111_CYCLE_SM.FLIP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6403\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5779\,
            sr => \N__5743\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5779\,
            sr => \N__5743\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5701\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5779\,
            sr => \N__5743\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5779\,
            sr => \N__5743\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5779\,
            sr => \N__5743\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5694\,
            in1 => \N__5657\,
            in2 => \_gnd_net_\,
            in3 => \N__6348\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6349\,
            in1 => \N__5630\,
            in2 => \_gnd_net_\,
            in3 => \N__5610\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6351\,
            in1 => \N__6563\,
            in2 => \_gnd_net_\,
            in3 => \N__6547\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6494\,
            in1 => \N__6478\,
            in2 => \_gnd_net_\,
            in3 => \N__6350\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6422\,
            in1 => \N__6402\,
            in2 => \_gnd_net_\,
            in3 => \N__6361\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIFAQ22_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6214\,
            in1 => \N__6822\,
            in2 => \_gnd_net_\,
            in3 => \N__6173\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6109\,
            lcout => \U111_CYCLE_SM.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU5SM1_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6823\,
            in1 => \N__6064\,
            in2 => \_gnd_net_\,
            in3 => \N__6023\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIHCQ22_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5977\,
            in1 => \N__6769\,
            in2 => \_gnd_net_\,
            in3 => \N__5942\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQ1SM1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5890\,
            in1 => \N__6770\,
            in2 => \_gnd_net_\,
            in3 => \N__5855\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPKQ22_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6913\,
            in1 => \N__6771\,
            in2 => \_gnd_net_\,
            in3 => \N__6602\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 13 2025 21:12:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    PRnW : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    BLSn : out std_logic;
    TCIn : out std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_iso_i\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_STATE_3C_net\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.N_592_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_482_cascade_\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_483\ : std_logic;
signal \U712_CHIP_RAM.N_335_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_507_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_477\ : std_logic;
signal \U712_CHIP_RAM.N_477_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.N_406_cascade_\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_OUTC_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_478\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER19_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_349_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_349\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.N_509\ : std_logic;
signal \U712_CHIP_RAM.N_509_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_504\ : std_logic;
signal \U712_CHIP_RAM.N_583_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_591\ : std_logic;
signal \U712_CHIP_RAM.N_402_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_375_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_375_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_402\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_426\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_586\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \U712_CHIP_RAM.N_586_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_419_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_332_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_510_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.N_343_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_334\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_366_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_335\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_1_cascade_\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \DRDDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_503_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_420\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_590\ : std_logic;
signal \U712_CHIP_RAM.N_476\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_248_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_358_i_cascade_\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_STATE_1C_net\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM.N_352_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.N_429\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_493\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.N_383\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_343\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_514_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_350\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_501\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_481_cascade_\ : std_logic;
signal \U712_REG_SM.N_428_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_500\ : std_logic;
signal \U712_CHIP_RAM.N_503\ : std_logic;
signal \U712_CHIP_RAM.N_500_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_514\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_337\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_332\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.N_248_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \C3_c\ : std_logic;
signal \BLSn_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_345_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_396\ : std_logic;
signal \U712_REG_SM.N_435_cascade_\ : std_logic;
signal \U712_REG_SM.N_352\ : std_logic;
signal \U712_REG_SM.N_357\ : std_logic;
signal \U712_REG_SM.N_353\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_450\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_510\ : std_logic;
signal \U712_CHIP_RAM.N_461\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \PRnW_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_351_cascade_\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_448_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.N_365\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_4\ : std_logic;
signal \U712_REG_SM.N_588\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_8\ : std_logic;
signal \U712_REG_SM.N_395_cascade_\ : std_logic;
signal \U712_REG_SM.N_439_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_5_iv_0_0\ : std_logic;
signal \U712_REG_SM.N_395\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_131\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_7\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_196_i\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_492\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_351\ : std_logic;
signal \U712_REG_SM.N_435\ : std_logic;
signal \U712_REG_SM.N_345\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_131_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \N_412_i\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_BYTE_ENABLE.N_467\ : std_logic;
signal \U712_BYTE_ENABLE.N_455_cascade_\ : std_logic;
signal \N_38_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_455\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_\ : std_logic;
signal \N_209_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_331_i\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \N_205\ : std_logic;
signal \N_411_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_213\ : std_logic;
signal \U712_BYTE_ENABLE.N_464\ : std_logic;
signal \N_40_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_452\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \N_208_i\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_456\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \PRnW_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \BLSn_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    PRnW <= \PRnW_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    BLSn <= \BLSn_wire\;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    TCIn <= \TCIn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4521\,
            RESETB => \N__8409\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12850\,
            DIN => \N__12849\,
            DOUT => \N__12848\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12850\,
            PADOUT => \N__12849\,
            PADIN => \N__12848\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12841\,
            DIN => \N__12840\,
            DOUT => \N__12839\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12841\,
            PADOUT => \N__12840\,
            PADIN => \N__12839\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12832\,
            DIN => \N__12831\,
            DOUT => \N__12830\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12832\,
            PADOUT => \N__12831\,
            PADIN => \N__12830\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7635\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12823\,
            DIN => \N__12822\,
            DOUT => \N__12821\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12823\,
            PADOUT => \N__12822\,
            PADIN => \N__12821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12814\,
            DIN => \N__12813\,
            DOUT => \N__12812\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12814\,
            PADOUT => \N__12813\,
            PADIN => \N__12812\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12805\,
            DIN => \N__12804\,
            DOUT => \N__12803\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12805\,
            PADOUT => \N__12804\,
            PADIN => \N__12803\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12796\,
            DIN => \N__12795\,
            DOUT => \N__12794\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12796\,
            PADOUT => \N__12795\,
            PADIN => \N__12794\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12787\,
            DIN => \N__12786\,
            DOUT => \N__12785\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12787\,
            PADOUT => \N__12786\,
            PADIN => \N__12785\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12778\,
            DIN => \N__12777\,
            DOUT => \N__12776\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12778\,
            PADOUT => \N__12777\,
            PADIN => \N__12776\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12769\,
            DIN => \N__12768\,
            DOUT => \N__12767\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12769\,
            PADOUT => \N__12768\,
            PADIN => \N__12767\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12760\,
            DIN => \N__12759\,
            DOUT => \N__12758\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12760\,
            PADOUT => \N__12759\,
            PADIN => \N__12758\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12751\,
            DIN => \N__12750\,
            DOUT => \N__12749\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12751\,
            PADOUT => \N__12750\,
            PADIN => \N__12749\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6084\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12742\,
            DIN => \N__12741\,
            DOUT => \N__12740\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12742\,
            PADOUT => \N__12741\,
            PADIN => \N__12740\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11058\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12733\,
            DIN => \N__12732\,
            DOUT => \N__12731\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12733\,
            PADOUT => \N__12732\,
            PADIN => \N__12731\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12724\,
            DIN => \N__12723\,
            DOUT => \N__12722\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12724\,
            PADOUT => \N__12723\,
            PADIN => \N__12722\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8114\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12715\,
            DIN => \N__12714\,
            DOUT => \N__12713\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12715\,
            PADOUT => \N__12714\,
            PADIN => \N__12713\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12706\,
            DIN => \N__12705\,
            DOUT => \N__12704\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12706\,
            PADOUT => \N__12705\,
            PADIN => \N__12704\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12697\,
            DIN => \N__12696\,
            DOUT => \N__12695\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12697\,
            PADOUT => \N__12696\,
            PADIN => \N__12695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12688\,
            DIN => \N__12687\,
            DOUT => \N__12686\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12688\,
            PADOUT => \N__12687\,
            PADIN => \N__12686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12679\,
            DIN => \N__12678\,
            DOUT => \N__12677\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12679\,
            PADOUT => \N__12678\,
            PADIN => \N__12677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12670\,
            DIN => \N__12669\,
            DOUT => \N__12668\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12670\,
            PADOUT => \N__12669\,
            PADIN => \N__12668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5079\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12661\,
            DIN => \N__12660\,
            DOUT => \N__12659\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12661\,
            PADOUT => \N__12660\,
            PADIN => \N__12659\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12652\,
            DIN => \N__12651\,
            DOUT => \N__12650\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12652\,
            PADOUT => \N__12651\,
            PADIN => \N__12650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12643\,
            DIN => \N__12642\,
            DOUT => \N__12641\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12643\,
            PADOUT => \N__12642\,
            PADIN => \N__12641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12634\,
            DIN => \N__12633\,
            DOUT => \N__12632\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12634\,
            PADOUT => \N__12633\,
            PADIN => \N__12632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12625\,
            DIN => \N__12624\,
            DOUT => \N__12623\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12625\,
            PADOUT => \N__12624\,
            PADIN => \N__12623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5775\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12616\,
            DIN => \N__12615\,
            DOUT => \N__12614\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12616\,
            PADOUT => \N__12615\,
            PADIN => \N__12614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12607\,
            DIN => \N__12606\,
            DOUT => \N__12605\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12607\,
            PADOUT => \N__12606\,
            PADIN => \N__12605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12598\,
            DIN => \N__12597\,
            DOUT => \N__12596\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12598\,
            PADOUT => \N__12597\,
            PADIN => \N__12596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12589\,
            DIN => \N__12588\,
            DOUT => \N__12587\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12589\,
            PADOUT => \N__12588\,
            PADIN => \N__12587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12580\,
            DIN => \N__12579\,
            DOUT => \N__12578\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12580\,
            PADOUT => \N__12579\,
            PADIN => \N__12578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12571\,
            DIN => \N__12570\,
            DOUT => \N__12569\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12571\,
            PADOUT => \N__12570\,
            PADIN => \N__12569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5265\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12562\,
            DIN => \N__12561\,
            DOUT => \N__12560\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12562\,
            PADOUT => \N__12561\,
            PADIN => \N__12560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12553\,
            DIN => \N__12552\,
            DOUT => \N__12551\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12553\,
            PADOUT => \N__12552\,
            PADIN => \N__12551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12544\,
            DIN => \N__12543\,
            DOUT => \N__12542\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12544\,
            PADOUT => \N__12543\,
            PADIN => \N__12542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12535\,
            DIN => \N__12534\,
            DOUT => \N__12533\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12535\,
            PADOUT => \N__12534\,
            PADIN => \N__12533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12526\,
            DIN => \N__12525\,
            DOUT => \N__12524\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12526\,
            PADOUT => \N__12525\,
            PADIN => \N__12524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12517\,
            DIN => \N__12516\,
            DOUT => \N__12515\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12517\,
            PADOUT => \N__12516\,
            PADIN => \N__12515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7572\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12508\,
            DIN => \N__12507\,
            DOUT => \N__12506\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12508\,
            PADOUT => \N__12507\,
            PADIN => \N__12506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12499\,
            DIN => \N__12498\,
            DOUT => \N__12497\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12499\,
            PADOUT => \N__12498\,
            PADIN => \N__12497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12490\,
            DIN => \N__12489\,
            DOUT => \N__12488\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12490\,
            PADOUT => \N__12489\,
            PADIN => \N__12488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9375\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12481\,
            DIN => \N__12480\,
            DOUT => \N__12479\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12481\,
            PADOUT => \N__12480\,
            PADIN => \N__12479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12472\,
            DIN => \N__12471\,
            DOUT => \N__12470\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12472\,
            PADOUT => \N__12471\,
            PADIN => \N__12470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12463\,
            DIN => \N__12462\,
            DOUT => \N__12461\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12463\,
            PADOUT => \N__12462\,
            PADIN => \N__12461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12454\,
            DIN => \N__12453\,
            DOUT => \N__12452\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12454\,
            PADOUT => \N__12453\,
            PADIN => \N__12452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6132\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12445\,
            DIN => \N__12444\,
            DOUT => \N__12443\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12445\,
            PADOUT => \N__12444\,
            PADIN => \N__12443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12436\,
            DIN => \N__12435\,
            DOUT => \N__12434\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12436\,
            PADOUT => \N__12435\,
            PADIN => \N__12434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11382\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12427\,
            DIN => \N__12426\,
            DOUT => \N__12425\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12427\,
            PADOUT => \N__12426\,
            PADIN => \N__12425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12418\,
            DIN => \N__12417\,
            DOUT => \N__12416\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12418\,
            PADOUT => \N__12417\,
            PADIN => \N__12416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5325\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12409\,
            DIN => \N__12408\,
            DOUT => \N__12407\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12409\,
            PADOUT => \N__12408\,
            PADIN => \N__12407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11943\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12400\,
            DIN => \N__12399\,
            DOUT => \N__12398\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12400\,
            PADOUT => \N__12399\,
            PADIN => \N__12398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12391\,
            DIN => \N__12390\,
            DOUT => \N__12389\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12391\,
            PADOUT => \N__12390\,
            PADIN => \N__12389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12382\,
            DIN => \N__12381\,
            DOUT => \N__12380\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12382\,
            PADOUT => \N__12381\,
            PADIN => \N__12380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4770\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12373\,
            DIN => \N__12372\,
            DOUT => \N__12371\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12373\,
            PADOUT => \N__12372\,
            PADIN => \N__12371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12364\,
            DIN => \N__12363\,
            DOUT => \N__12362\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12364\,
            PADOUT => \N__12363\,
            PADIN => \N__12362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12355\,
            DIN => \N__12354\,
            DOUT => \N__12353\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12355\,
            PADOUT => \N__12354\,
            PADIN => \N__12353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5058\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12346\,
            DIN => \N__12345\,
            DOUT => \N__12344\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12346\,
            PADOUT => \N__12345\,
            PADIN => \N__12344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12337\,
            DIN => \N__12336\,
            DOUT => \N__12335\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12337\,
            PADOUT => \N__12336\,
            PADIN => \N__12335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12328\,
            DIN => \N__12327\,
            DOUT => \N__12326\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12328\,
            PADOUT => \N__12327\,
            PADIN => \N__12326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11298\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12319\,
            DIN => \N__12318\,
            DOUT => \N__12317\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12319\,
            PADOUT => \N__12318\,
            PADIN => \N__12317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5770\,
            DIN0 => OPEN,
            DOUT0 => \N__4665\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12310\,
            DIN => \N__12309\,
            DOUT => \N__12308\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12310\,
            PADOUT => \N__12309\,
            PADIN => \N__12308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12301\,
            DIN => \N__12300\,
            DOUT => \N__12299\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12301\,
            PADOUT => \N__12300\,
            PADIN => \N__12299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12292\,
            DIN => \N__12291\,
            DOUT => \N__12290\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12292\,
            PADOUT => \N__12291\,
            PADIN => \N__12290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12283\,
            DIN => \N__12282\,
            DOUT => \N__12281\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12283\,
            PADOUT => \N__12282\,
            PADIN => \N__12281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5991\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12274\,
            DIN => \N__12273\,
            DOUT => \N__12272\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12274\,
            PADOUT => \N__12273\,
            PADIN => \N__12272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12265\,
            DIN => \N__12264\,
            DOUT => \N__12263\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12265\,
            PADOUT => \N__12264\,
            PADIN => \N__12263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12256\,
            DIN => \N__12255\,
            DOUT => \N__12254\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12256\,
            PADOUT => \N__12255\,
            PADIN => \N__12254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12247\,
            DIN => \N__12246\,
            DOUT => \N__12245\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12247\,
            PADOUT => \N__12246\,
            PADIN => \N__12245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12238\,
            DIN => \N__12237\,
            DOUT => \N__12236\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12238\,
            PADOUT => \N__12237\,
            PADIN => \N__12236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12229\,
            DIN => \N__12228\,
            DOUT => \N__12227\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12229\,
            PADOUT => \N__12228\,
            PADIN => \N__12227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5040\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12220\,
            DIN => \N__12219\,
            DOUT => \N__12218\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12220\,
            PADOUT => \N__12219\,
            PADIN => \N__12218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12211\,
            DIN => \N__12210\,
            DOUT => \N__12209\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12211\,
            PADOUT => \N__12210\,
            PADIN => \N__12209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12202\,
            DIN => \N__12201\,
            DOUT => \N__12200\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12202\,
            PADOUT => \N__12201\,
            PADIN => \N__12200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4929\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12193\,
            DIN => \N__12192\,
            DOUT => \N__12191\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12193\,
            PADOUT => \N__12192\,
            PADIN => \N__12191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12184\,
            DIN => \N__12183\,
            DOUT => \N__12182\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12184\,
            PADOUT => \N__12183\,
            PADIN => \N__12182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12175\,
            DIN => \N__12174\,
            DOUT => \N__12173\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12175\,
            PADOUT => \N__12174\,
            PADIN => \N__12173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6117\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12166\,
            DIN => \N__12165\,
            DOUT => \N__12164\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12166\,
            PADOUT => \N__12165\,
            PADIN => \N__12164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12157\,
            DIN => \N__12156\,
            DOUT => \N__12155\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12157\,
            PADOUT => \N__12156\,
            PADIN => \N__12155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12148\,
            DIN => \N__12147\,
            DOUT => \N__12146\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12148\,
            PADOUT => \N__12147\,
            PADIN => \N__12146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7680\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12139\,
            DIN => \N__12138\,
            DOUT => \N__12137\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12139\,
            PADOUT => \N__12138\,
            PADIN => \N__12137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5895\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12130\,
            DIN => \N__12129\,
            DOUT => \N__12128\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12130\,
            PADOUT => \N__12129\,
            PADIN => \N__12128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4602\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRnW_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12121\,
            DIN => \N__12120\,
            DOUT => \N__12119\,
            PACKAGEPIN => \PRnW_wire\
        );

    \PRnW_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12121\,
            PADOUT => \N__12120\,
            PADIN => \N__12119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8250\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12112\,
            DIN => \N__12111\,
            DOUT => \N__12110\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12112\,
            PADOUT => \N__12111\,
            PADIN => \N__12110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12103\,
            DIN => \N__12102\,
            DOUT => \N__12101\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12103\,
            PADOUT => \N__12102\,
            PADIN => \N__12101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4601\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12094\,
            DIN => \N__12093\,
            DOUT => \N__12092\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12094\,
            PADOUT => \N__12093\,
            PADIN => \N__12092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4539\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12085\,
            DIN => \N__12084\,
            DOUT => \N__12083\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12085\,
            PADOUT => \N__12084\,
            PADIN => \N__12083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12076\,
            DIN => \N__12075\,
            DOUT => \N__12074\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12076\,
            PADOUT => \N__12075\,
            PADIN => \N__12074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12067\,
            DIN => \N__12066\,
            DOUT => \N__12065\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12067\,
            PADOUT => \N__12066\,
            PADIN => \N__12065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12058\,
            DIN => \N__12057\,
            DOUT => \N__12056\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12058\,
            PADOUT => \N__12057\,
            PADIN => \N__12056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BLSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12049\,
            DIN => \N__12048\,
            DOUT => \N__12047\,
            PACKAGEPIN => \BLSn_wire\
        );

    \BLSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12049\,
            PADOUT => \N__12048\,
            PADIN => \N__12047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7458\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12040\,
            DIN => \N__12039\,
            DOUT => \N__12038\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12040\,
            PADOUT => \N__12039\,
            PADIN => \N__12038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12031\,
            DIN => \N__12030\,
            DOUT => \N__12029\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12031\,
            PADOUT => \N__12030\,
            PADIN => \N__12029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12022\,
            DIN => \N__12021\,
            DOUT => \N__12020\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12022\,
            PADOUT => \N__12021\,
            PADIN => \N__12020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8805\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12013\,
            DIN => \N__12012\,
            DOUT => \N__12011\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12013\,
            PADOUT => \N__12012\,
            PADIN => \N__12011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10083\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12004\,
            DIN => \N__12003\,
            DOUT => \N__12002\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12004\,
            PADOUT => \N__12003\,
            PADIN => \N__12002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11995\,
            DIN => \N__11994\,
            DOUT => \N__11993\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11995\,
            PADOUT => \N__11994\,
            PADIN => \N__11993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11986\,
            DIN => \N__11985\,
            DOUT => \N__11984\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11986\,
            PADOUT => \N__11985\,
            PADIN => \N__11984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11977\,
            DIN => \N__11976\,
            DOUT => \N__11975\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11977\,
            PADOUT => \N__11976\,
            PADIN => \N__11975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5774\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2876\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11955\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__11955\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\
        );

    \I__2874\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11949\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__11949\,
            I => \U712_BYTE_ENABLE.N_455\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__11946\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_\
        );

    \I__2871\ : IoInMux
    port map (
            O => \N__11943\,
            I => \N__11940\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__11940\,
            I => \N__11937\
        );

    \I__2869\ : Span4Mux_s1_h
    port map (
            O => \N__11937\,
            I => \N__11934\
        );

    \I__2868\ : Sp12to4
    port map (
            O => \N__11934\,
            I => \N__11931\
        );

    \I__2867\ : Span12Mux_s11_v
    port map (
            O => \N__11931\,
            I => \N__11928\
        );

    \I__2866\ : Span12Mux_h
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__11925\,
            I => \N_209_i\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__11922\,
            I => \N__11918\
        );

    \I__2863\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11915\
        );

    \I__2862\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__11915\,
            I => \U712_BYTE_ENABLE.N_331_i\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__11912\,
            I => \U712_BYTE_ENABLE.N_331_i\
        );

    \I__2859\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11894\
        );

    \I__2858\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11894\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11894\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__11904\,
            I => \N__11890\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__11903\,
            I => \N__11887\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11883\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11880\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__11894\,
            I => \N__11877\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11865\
        );

    \I__2850\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11860\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11856\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11853\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11848\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__11880\,
            I => \N__11848\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__11877\,
            I => \N__11845\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11840\
        );

    \I__2843\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11840\
        );

    \I__2842\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11832\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11832\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11832\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11825\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11825\
        );

    \I__2837\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11825\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11822\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11819\
        );

    \I__2834\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11814\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11814\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__11860\,
            I => \N__11810\
        );

    \I__2831\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11807\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11804\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11799\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__11848\,
            I => \N__11799\
        );

    \I__2827\ : Span4Mux_h
    port map (
            O => \N__11845\,
            I => \N__11794\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11794\
        );

    \I__2825\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11791\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11788\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11825\,
            I => \N__11779\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11822\,
            I => \N__11779\
        );

    \I__2821\ : Span4Mux_h
    port map (
            O => \N__11819\,
            I => \N__11779\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11814\,
            I => \N__11779\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11776\
        );

    \I__2818\ : Odrv12
    port map (
            O => \N__11810\,
            I => \CPU_CYCLEm\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__11807\,
            I => \CPU_CYCLEm\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__11804\,
            I => \CPU_CYCLEm\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__11799\,
            I => \CPU_CYCLEm\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__11794\,
            I => \CPU_CYCLEm\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11791\,
            I => \CPU_CYCLEm\
        );

    \I__2812\ : Odrv12
    port map (
            O => \N__11788\,
            I => \CPU_CYCLEm\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__11779\,
            I => \CPU_CYCLEm\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__11776\,
            I => \CPU_CYCLEm\
        );

    \I__2809\ : IoInMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2807\ : IoSpan4Mux
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__2806\ : Span4Mux_s3_v
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__11745\,
            I => \N__11742\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__11742\,
            I => \N_205\
        );

    \I__2803\ : IoInMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__2801\ : Span4Mux_s3_v
    port map (
            O => \N__11733\,
            I => \N__11730\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__11730\,
            I => \N_411_i\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11721\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11714\
        );

    \I__2797\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11714\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11714\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11706\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11714\,
            I => \N__11706\
        );

    \I__2793\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11701\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11701\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11698\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__11706\,
            I => \N__11695\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11701\,
            I => \N__11690\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__11698\,
            I => \N__11690\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__11695\,
            I => \N__11684\
        );

    \I__2786\ : Span4Mux_v
    port map (
            O => \N__11690\,
            I => \N__11684\
        );

    \I__2785\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11681\
        );

    \I__2784\ : Sp12to4
    port map (
            O => \N__11684\,
            I => \N__11676\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__11681\,
            I => \N__11676\
        );

    \I__2782\ : Span12Mux_h
    port map (
            O => \N__11676\,
            I => \N__11673\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__11673\,
            I => \A_c_1\
        );

    \I__2780\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11666\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11658\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11666\,
            I => \N__11655\
        );

    \I__2777\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11650\
        );

    \I__2776\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11650\
        );

    \I__2775\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11645\
        );

    \I__2774\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11645\
        );

    \I__2773\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11642\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11658\,
            I => \N__11639\
        );

    \I__2771\ : Span4Mux_h
    port map (
            O => \N__11655\,
            I => \N__11633\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11633\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11645\,
            I => \N__11628\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11628\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__11639\,
            I => \N__11625\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11622\
        );

    \I__2765\ : Span4Mux_v
    port map (
            O => \N__11633\,
            I => \N__11616\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__11628\,
            I => \N__11616\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__11625\,
            I => \N__11611\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__11622\,
            I => \N__11611\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11608\
        );

    \I__2760\ : Sp12to4
    port map (
            O => \N__11616\,
            I => \N__11605\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__11611\,
            I => \N__11602\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11608\,
            I => \N__11599\
        );

    \I__2757\ : Span12Mux_h
    port map (
            O => \N__11605\,
            I => \N__11592\
        );

    \I__2756\ : Sp12to4
    port map (
            O => \N__11602\,
            I => \N__11592\
        );

    \I__2755\ : Span12Mux_s10_v
    port map (
            O => \N__11599\,
            I => \N__11592\
        );

    \I__2754\ : Odrv12
    port map (
            O => \N__11592\,
            I => \A_c_0\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__11589\,
            I => \N__11584\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__11588\,
            I => \N__11579\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \N__11576\
        );

    \I__2750\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11570\
        );

    \I__2749\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11570\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__11582\,
            I => \N__11567\
        );

    \I__2747\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11562\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11562\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \N__11559\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__11570\,
            I => \N__11555\
        );

    \I__2743\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11552\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__11562\,
            I => \N__11548\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11545\
        );

    \I__2740\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11542\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__11555\,
            I => \N__11537\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__11552\,
            I => \N__11537\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11533\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__11548\,
            I => \N__11530\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11545\,
            I => \N__11525\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11542\,
            I => \N__11525\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__11537\,
            I => \N__11522\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11519\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11516\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__11530\,
            I => \N__11511\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__11525\,
            I => \N__11511\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__11522\,
            I => \N__11508\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11503\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__11516\,
            I => \N__11503\
        );

    \I__2725\ : Span4Mux_v
    port map (
            O => \N__11511\,
            I => \N__11500\
        );

    \I__2724\ : Sp12to4
    port map (
            O => \N__11508\,
            I => \N__11495\
        );

    \I__2723\ : Span12Mux_v
    port map (
            O => \N__11503\,
            I => \N__11495\
        );

    \I__2722\ : Sp12to4
    port map (
            O => \N__11500\,
            I => \N__11492\
        );

    \I__2721\ : Span12Mux_h
    port map (
            O => \N__11495\,
            I => \N__11489\
        );

    \I__2720\ : Span12Mux_h
    port map (
            O => \N__11492\,
            I => \N__11486\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__11489\,
            I => \SIZ_c_1\
        );

    \I__2718\ : Odrv12
    port map (
            O => \N__11486\,
            I => \SIZ_c_1\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11477\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11474\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__11477\,
            I => \N__11465\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__11474\,
            I => \N__11465\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11462\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11457\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11457\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11454\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__11465\,
            I => \N__11448\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11462\,
            I => \N__11448\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11457\,
            I => \N__11443\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11454\,
            I => \N__11443\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11440\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__11448\,
            I => \N__11437\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__11443\,
            I => \N__11434\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11431\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__11437\,
            I => \N__11427\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__11434\,
            I => \N__11422\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__11431\,
            I => \N__11422\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11419\
        );

    \I__2697\ : Sp12to4
    port map (
            O => \N__11427\,
            I => \N__11416\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__11422\,
            I => \N__11413\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11410\
        );

    \I__2694\ : Span12Mux_h
    port map (
            O => \N__11416\,
            I => \N__11403\
        );

    \I__2693\ : Sp12to4
    port map (
            O => \N__11413\,
            I => \N__11403\
        );

    \I__2692\ : Span12Mux_v
    port map (
            O => \N__11410\,
            I => \N__11403\
        );

    \I__2691\ : Odrv12
    port map (
            O => \N__11403\,
            I => \SIZ_c_0\
        );

    \I__2690\ : IoInMux
    port map (
            O => \N__11400\,
            I => \N__11397\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11397\,
            I => \N__11394\
        );

    \I__2688\ : Span4Mux_s3_v
    port map (
            O => \N__11394\,
            I => \N__11391\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__11391\,
            I => \N_213\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11385\,
            I => \U712_BYTE_ENABLE.N_464\
        );

    \I__2684\ : IoInMux
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11379\,
            I => \N__11376\
        );

    \I__2682\ : Sp12to4
    port map (
            O => \N__11376\,
            I => \N__11373\
        );

    \I__2681\ : Span12Mux_h
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__2680\ : Span12Mux_v
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__2679\ : Odrv12
    port map (
            O => \N__11367\,
            I => \N_40_i\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11361\,
            I => \U712_BYTE_ENABLE.N_452\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11352\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11352\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11352\,
            I => \N__11346\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11343\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11340\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__11349\,
            I => \N__11336\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__11346\,
            I => \N__11333\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11343\,
            I => \N__11328\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11340\,
            I => \N__11328\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11323\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11323\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__11333\,
            I => \N__11318\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__11328\,
            I => \N__11318\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11315\
        );

    \I__2662\ : Span4Mux_h
    port map (
            O => \N__11318\,
            I => \N__11310\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__11315\,
            I => \N__11310\
        );

    \I__2660\ : Sp12to4
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__2659\ : Span12Mux_h
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__2658\ : Span12Mux_v
    port map (
            O => \N__11304\,
            I => \N__11301\
        );

    \I__2657\ : Odrv12
    port map (
            O => \N__11301\,
            I => \CASUn_c\
        );

    \I__2656\ : IoInMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__2654\ : Span4Mux_s3_h
    port map (
            O => \N__11292\,
            I => \N__11289\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__11289\,
            I => \N__11286\
        );

    \I__2652\ : Span4Mux_h
    port map (
            O => \N__11286\,
            I => \N__11283\
        );

    \I__2651\ : Span4Mux_h
    port map (
            O => \N__11283\,
            I => \N__11280\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__11280\,
            I => \N_208_i\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11273\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__11276\,
            I => \N__11269\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11273\,
            I => \N__11264\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11261\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11255\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11255\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11252\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__11264\,
            I => \N__11247\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11261\,
            I => \N__11247\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11244\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11255\,
            I => \N__11241\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11252\,
            I => \N__11238\
        );

    \I__2637\ : Sp12to4
    port map (
            O => \N__11247\,
            I => \N__11235\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11232\
        );

    \I__2635\ : Span12Mux_h
    port map (
            O => \N__11241\,
            I => \N__11229\
        );

    \I__2634\ : Span12Mux_v
    port map (
            O => \N__11238\,
            I => \N__11226\
        );

    \I__2633\ : Span12Mux_h
    port map (
            O => \N__11235\,
            I => \N__11223\
        );

    \I__2632\ : Span12Mux_v
    port map (
            O => \N__11232\,
            I => \N__11220\
        );

    \I__2631\ : Span12Mux_v
    port map (
            O => \N__11229\,
            I => \N__11217\
        );

    \I__2630\ : Span12Mux_h
    port map (
            O => \N__11226\,
            I => \N__11214\
        );

    \I__2629\ : Span12Mux_v
    port map (
            O => \N__11223\,
            I => \N__11209\
        );

    \I__2628\ : Span12Mux_h
    port map (
            O => \N__11220\,
            I => \N__11209\
        );

    \I__2627\ : Odrv12
    port map (
            O => \N__11217\,
            I => \CASLn_c\
        );

    \I__2626\ : Odrv12
    port map (
            O => \N__11214\,
            I => \CASLn_c\
        );

    \I__2625\ : Odrv12
    port map (
            O => \N__11209\,
            I => \CASLn_c\
        );

    \I__2624\ : IoInMux
    port map (
            O => \N__11202\,
            I => \N__11199\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__11199\,
            I => \N__11195\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11191\
        );

    \I__2621\ : IoSpan4Mux
    port map (
            O => \N__11195\,
            I => \N__11186\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11183\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11178\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11178\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11175\
        );

    \I__2616\ : Span4Mux_s2_v
    port map (
            O => \N__11186\,
            I => \N__11172\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__11183\,
            I => \N__11165\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11178\,
            I => \N__11165\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11165\
        );

    \I__2612\ : Sp12to4
    port map (
            O => \N__11172\,
            I => \N__11162\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__11165\,
            I => \N__11159\
        );

    \I__2610\ : Span12Mux_v
    port map (
            O => \N__11162\,
            I => \N__11155\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__11159\,
            I => \N__11152\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11149\
        );

    \I__2607\ : Odrv12
    port map (
            O => \N__11155\,
            I => \DBENn_c\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__11152\,
            I => \DBENn_c\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11149\,
            I => \DBENn_c\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__11142\,
            I => \N__11136\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11133\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11130\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11127\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11123\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__11133\,
            I => \N__11118\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__11130\,
            I => \N__11118\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__11127\,
            I => \N__11115\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11112\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11108\
        );

    \I__2594\ : Span4Mux_h
    port map (
            O => \N__11118\,
            I => \N__11101\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__11115\,
            I => \N__11101\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11101\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11098\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__11108\,
            I => \N__11094\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__11101\,
            I => \N__11089\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__11098\,
            I => \N__11089\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11097\,
            I => \N__11085\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__11094\,
            I => \N__11082\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__11089\,
            I => \N__11079\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11076\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11073\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__11082\,
            I => \DMA_CYCLEm\
        );

    \I__2581\ : Odrv4
    port map (
            O => \N__11079\,
            I => \DMA_CYCLEm\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__11076\,
            I => \DMA_CYCLEm\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__11073\,
            I => \DMA_CYCLEm\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__11061\,
            I => \U712_BYTE_ENABLE.N_456\
        );

    \I__2576\ : IoInMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2574\ : Span4Mux_s0_v
    port map (
            O => \N__11052\,
            I => \N__11049\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__11046\,
            I => \N_412_i\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__11043\,
            I => \N__11039\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11030\
        );

    \I__2569\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11027\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11038\,
            I => \N__11024\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11037\,
            I => \N__11021\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11016\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__11035\,
            I => \N__11011\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__11034\,
            I => \N__11007\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__11033\,
            I => \N__11002\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__10998\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11027\,
            I => \N__10995\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__10989\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__11021\,
            I => \N__10989\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11020\,
            I => \N__10986\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11019\,
            I => \N__10983\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__10977\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11015\,
            I => \N__10974\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10963\
        );

    \I__2553\ : InMux
    port map (
            O => \N__11011\,
            I => \N__10963\
        );

    \I__2552\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10963\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11007\,
            I => \N__10963\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10963\
        );

    \I__2549\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10960\
        );

    \I__2548\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10955\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10955\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__10998\,
            I => \N__10950\
        );

    \I__2545\ : Span4Mux_v
    port map (
            O => \N__10995\,
            I => \N__10950\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10947\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__10989\,
            I => \N__10940\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10986\,
            I => \N__10940\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10940\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10937\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10934\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10931\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10928\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10919\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10919\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10960\,
            I => \N__10919\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10919\
        );

    \I__2532\ : Sp12to4
    port map (
            O => \N__10950\,
            I => \N__10915\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10904\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__10940\,
            I => \N__10904\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10904\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10904\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10904\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__10928\,
            I => \N__10899\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__10919\,
            I => \N__10899\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10896\
        );

    \I__2523\ : Span12Mux_h
    port map (
            O => \N__10915\,
            I => \N__10891\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__10904\,
            I => \N__10891\
        );

    \I__2521\ : Sp12to4
    port map (
            O => \N__10899\,
            I => \N__10888\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10885\
        );

    \I__2519\ : Span12Mux_v
    port map (
            O => \N__10891\,
            I => \N__10882\
        );

    \I__2518\ : Span12Mux_h
    port map (
            O => \N__10888\,
            I => \N__10879\
        );

    \I__2517\ : Span12Mux_v
    port map (
            O => \N__10885\,
            I => \N__10876\
        );

    \I__2516\ : Span12Mux_h
    port map (
            O => \N__10882\,
            I => \N__10873\
        );

    \I__2515\ : Span12Mux_v
    port map (
            O => \N__10879\,
            I => \N__10868\
        );

    \I__2514\ : Span12Mux_h
    port map (
            O => \N__10876\,
            I => \N__10868\
        );

    \I__2513\ : Odrv12
    port map (
            O => \N__10873\,
            I => \AGNUS_REV_c\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__10868\,
            I => \AGNUS_REV_c\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10858\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10855\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10851\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10848\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10855\,
            I => \N__10845\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10842\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10851\,
            I => \N__10839\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__10848\,
            I => \N__10836\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__10845\,
            I => \N__10831\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10842\,
            I => \N__10831\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__10839\,
            I => \N__10828\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__10836\,
            I => \N__10823\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__10831\,
            I => \N__10823\
        );

    \I__2498\ : Sp12to4
    port map (
            O => \N__10828\,
            I => \N__10820\
        );

    \I__2497\ : Sp12to4
    port map (
            O => \N__10823\,
            I => \N__10817\
        );

    \I__2496\ : Span12Mux_h
    port map (
            O => \N__10820\,
            I => \N__10814\
        );

    \I__2495\ : Span12Mux_h
    port map (
            O => \N__10817\,
            I => \N__10811\
        );

    \I__2494\ : Span12Mux_v
    port map (
            O => \N__10814\,
            I => \N__10808\
        );

    \I__2493\ : Span12Mux_v
    port map (
            O => \N__10811\,
            I => \N__10805\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__10808\,
            I => \DRA_c_9\
        );

    \I__2491\ : Odrv12
    port map (
            O => \N__10805\,
            I => \DRA_c_9\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10800\,
            I => \N__10797\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10797\,
            I => \N__10794\
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__10794\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2487\ : ClkMux
    port map (
            O => \N__10791\,
            I => \N__10773\
        );

    \I__2486\ : ClkMux
    port map (
            O => \N__10790\,
            I => \N__10773\
        );

    \I__2485\ : ClkMux
    port map (
            O => \N__10789\,
            I => \N__10773\
        );

    \I__2484\ : ClkMux
    port map (
            O => \N__10788\,
            I => \N__10773\
        );

    \I__2483\ : ClkMux
    port map (
            O => \N__10787\,
            I => \N__10773\
        );

    \I__2482\ : ClkMux
    port map (
            O => \N__10786\,
            I => \N__10773\
        );

    \I__2481\ : GlobalMux
    port map (
            O => \N__10773\,
            I => \N__10770\
        );

    \I__2480\ : gio2CtrlBuf
    port map (
            O => \N__10770\,
            I => \C3_c_g\
        );

    \I__2479\ : CEMux
    port map (
            O => \N__10767\,
            I => \N__10731\
        );

    \I__2478\ : CEMux
    port map (
            O => \N__10766\,
            I => \N__10731\
        );

    \I__2477\ : CEMux
    port map (
            O => \N__10765\,
            I => \N__10731\
        );

    \I__2476\ : CEMux
    port map (
            O => \N__10764\,
            I => \N__10731\
        );

    \I__2475\ : CEMux
    port map (
            O => \N__10763\,
            I => \N__10731\
        );

    \I__2474\ : CEMux
    port map (
            O => \N__10762\,
            I => \N__10731\
        );

    \I__2473\ : CEMux
    port map (
            O => \N__10761\,
            I => \N__10731\
        );

    \I__2472\ : CEMux
    port map (
            O => \N__10760\,
            I => \N__10731\
        );

    \I__2471\ : CEMux
    port map (
            O => \N__10759\,
            I => \N__10731\
        );

    \I__2470\ : CEMux
    port map (
            O => \N__10758\,
            I => \N__10731\
        );

    \I__2469\ : CEMux
    port map (
            O => \N__10757\,
            I => \N__10731\
        );

    \I__2468\ : CEMux
    port map (
            O => \N__10756\,
            I => \N__10731\
        );

    \I__2467\ : GlobalMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__2466\ : gio2CtrlBuf
    port map (
            O => \N__10728\,
            I => \DBRn_c_i_0_g\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10715\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10712\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10709\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10704\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10704\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10699\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10699\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10696\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10715\,
            I => \N__10693\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10678\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10669\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10661\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10699\,
            I => \N__10658\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10696\,
            I => \N__10643\
        );

    \I__2451\ : Glb2LocalMux
    port map (
            O => \N__10693\,
            I => \N__10557\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__10692\,
            I => \N__10557\
        );

    \I__2449\ : SRMux
    port map (
            O => \N__10691\,
            I => \N__10557\
        );

    \I__2448\ : SRMux
    port map (
            O => \N__10690\,
            I => \N__10557\
        );

    \I__2447\ : SRMux
    port map (
            O => \N__10689\,
            I => \N__10557\
        );

    \I__2446\ : SRMux
    port map (
            O => \N__10688\,
            I => \N__10557\
        );

    \I__2445\ : SRMux
    port map (
            O => \N__10687\,
            I => \N__10557\
        );

    \I__2444\ : SRMux
    port map (
            O => \N__10686\,
            I => \N__10557\
        );

    \I__2443\ : SRMux
    port map (
            O => \N__10685\,
            I => \N__10557\
        );

    \I__2442\ : SRMux
    port map (
            O => \N__10684\,
            I => \N__10557\
        );

    \I__2441\ : SRMux
    port map (
            O => \N__10683\,
            I => \N__10557\
        );

    \I__2440\ : SRMux
    port map (
            O => \N__10682\,
            I => \N__10557\
        );

    \I__2439\ : SRMux
    port map (
            O => \N__10681\,
            I => \N__10557\
        );

    \I__2438\ : Glb2LocalMux
    port map (
            O => \N__10678\,
            I => \N__10557\
        );

    \I__2437\ : SRMux
    port map (
            O => \N__10677\,
            I => \N__10557\
        );

    \I__2436\ : SRMux
    port map (
            O => \N__10676\,
            I => \N__10557\
        );

    \I__2435\ : SRMux
    port map (
            O => \N__10675\,
            I => \N__10557\
        );

    \I__2434\ : SRMux
    port map (
            O => \N__10674\,
            I => \N__10557\
        );

    \I__2433\ : SRMux
    port map (
            O => \N__10673\,
            I => \N__10557\
        );

    \I__2432\ : SRMux
    port map (
            O => \N__10672\,
            I => \N__10557\
        );

    \I__2431\ : Glb2LocalMux
    port map (
            O => \N__10669\,
            I => \N__10557\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__10668\,
            I => \N__10557\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__10667\,
            I => \N__10557\
        );

    \I__2428\ : SRMux
    port map (
            O => \N__10666\,
            I => \N__10557\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__10665\,
            I => \N__10557\
        );

    \I__2426\ : SRMux
    port map (
            O => \N__10664\,
            I => \N__10557\
        );

    \I__2425\ : Glb2LocalMux
    port map (
            O => \N__10661\,
            I => \N__10557\
        );

    \I__2424\ : Glb2LocalMux
    port map (
            O => \N__10658\,
            I => \N__10557\
        );

    \I__2423\ : SRMux
    port map (
            O => \N__10657\,
            I => \N__10557\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__10656\,
            I => \N__10557\
        );

    \I__2421\ : SRMux
    port map (
            O => \N__10655\,
            I => \N__10557\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__10654\,
            I => \N__10557\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__10653\,
            I => \N__10557\
        );

    \I__2418\ : SRMux
    port map (
            O => \N__10652\,
            I => \N__10557\
        );

    \I__2417\ : SRMux
    port map (
            O => \N__10651\,
            I => \N__10557\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__10650\,
            I => \N__10557\
        );

    \I__2415\ : SRMux
    port map (
            O => \N__10649\,
            I => \N__10557\
        );

    \I__2414\ : SRMux
    port map (
            O => \N__10648\,
            I => \N__10557\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__10647\,
            I => \N__10557\
        );

    \I__2412\ : SRMux
    port map (
            O => \N__10646\,
            I => \N__10557\
        );

    \I__2411\ : Glb2LocalMux
    port map (
            O => \N__10643\,
            I => \N__10557\
        );

    \I__2410\ : SRMux
    port map (
            O => \N__10642\,
            I => \N__10557\
        );

    \I__2409\ : GlobalMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__2408\ : gio2CtrlBuf
    port map (
            O => \N__10554\,
            I => \RESETn_c_i_g\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10547\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10544\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10547\,
            I => \N__10539\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10544\,
            I => \N__10539\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__2402\ : Sp12to4
    port map (
            O => \N__10536\,
            I => \N__10533\
        );

    \I__2401\ : Span12Mux_h
    port map (
            O => \N__10533\,
            I => \N__10530\
        );

    \I__2400\ : Odrv12
    port map (
            O => \N__10530\,
            I => \RAS0n_c\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10524\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10524\,
            I => \N__10521\
        );

    \I__2397\ : Sp12to4
    port map (
            O => \N__10521\,
            I => \N__10518\
        );

    \I__2396\ : Span12Mux_v
    port map (
            O => \N__10518\,
            I => \N__10515\
        );

    \I__2395\ : Span12Mux_h
    port map (
            O => \N__10515\,
            I => \N__10512\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__10512\,
            I => \RAS1n_c\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10493\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10488\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10488\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10485\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10480\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10480\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10473\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__10502\,
            I => \N__10468\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10461\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10461\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10461\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10456\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10456\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10447\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10436\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10488\,
            I => \N__10436\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10485\,
            I => \N__10436\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10480\,
            I => \N__10436\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10431\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10431\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10426\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10426\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10422\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10417\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10417\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10414\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10461\,
            I => \N__10409\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10409\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10398\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10398\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10398\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10398\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10398\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \N__10395\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10447\,
            I => \N__10391\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10386\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10386\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10379\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10431\,
            I => \N__10379\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10426\,
            I => \N__10379\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10376\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__10422\,
            I => \N__10366\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10366\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10366\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__10409\,
            I => \N__10360\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10398\,
            I => \N__10360\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10357\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10354\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10341\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10341\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__10379\,
            I => \N__10336\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10336\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10331\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10331\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10328\
        );

    \I__2338\ : Span4Mux_v
    port map (
            O => \N__10366\,
            I => \N__10325\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10322\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__10360\,
            I => \N__10315\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10357\,
            I => \N__10315\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10315\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10310\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10310\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10297\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10297\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10297\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10297\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10297\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10297\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__10341\,
            I => \N__10292\
        );

    \I__2324\ : Span4Mux_v
    port map (
            O => \N__10336\,
            I => \N__10292\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10289\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10286\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__10325\,
            I => \N__10282\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10322\,
            I => \N__10273\
        );

    \I__2319\ : Sp12to4
    port map (
            O => \N__10315\,
            I => \N__10273\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10273\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10273\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__10292\,
            I => \N__10266\
        );

    \I__2315\ : Span4Mux_v
    port map (
            O => \N__10289\,
            I => \N__10266\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__10286\,
            I => \N__10266\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10263\
        );

    \I__2312\ : Sp12to4
    port map (
            O => \N__10282\,
            I => \N__10254\
        );

    \I__2311\ : Span12Mux_v
    port map (
            O => \N__10273\,
            I => \N__10254\
        );

    \I__2310\ : Sp12to4
    port map (
            O => \N__10266\,
            I => \N__10254\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10263\,
            I => \N__10254\
        );

    \I__2308\ : Span12Mux_h
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__2307\ : Odrv12
    port map (
            O => \N__10251\,
            I => \RESETn_c\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10245\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10239\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10233\,
            I => \N__10188\
        );

    \I__2300\ : ClkMux
    port map (
            O => \N__10232\,
            I => \N__10095\
        );

    \I__2299\ : ClkMux
    port map (
            O => \N__10231\,
            I => \N__10095\
        );

    \I__2298\ : ClkMux
    port map (
            O => \N__10230\,
            I => \N__10095\
        );

    \I__2297\ : ClkMux
    port map (
            O => \N__10229\,
            I => \N__10095\
        );

    \I__2296\ : ClkMux
    port map (
            O => \N__10228\,
            I => \N__10095\
        );

    \I__2295\ : ClkMux
    port map (
            O => \N__10227\,
            I => \N__10095\
        );

    \I__2294\ : ClkMux
    port map (
            O => \N__10226\,
            I => \N__10095\
        );

    \I__2293\ : ClkMux
    port map (
            O => \N__10225\,
            I => \N__10095\
        );

    \I__2292\ : ClkMux
    port map (
            O => \N__10224\,
            I => \N__10095\
        );

    \I__2291\ : ClkMux
    port map (
            O => \N__10223\,
            I => \N__10095\
        );

    \I__2290\ : ClkMux
    port map (
            O => \N__10222\,
            I => \N__10095\
        );

    \I__2289\ : ClkMux
    port map (
            O => \N__10221\,
            I => \N__10095\
        );

    \I__2288\ : ClkMux
    port map (
            O => \N__10220\,
            I => \N__10095\
        );

    \I__2287\ : ClkMux
    port map (
            O => \N__10219\,
            I => \N__10095\
        );

    \I__2286\ : ClkMux
    port map (
            O => \N__10218\,
            I => \N__10095\
        );

    \I__2285\ : ClkMux
    port map (
            O => \N__10217\,
            I => \N__10095\
        );

    \I__2284\ : ClkMux
    port map (
            O => \N__10216\,
            I => \N__10095\
        );

    \I__2283\ : ClkMux
    port map (
            O => \N__10215\,
            I => \N__10095\
        );

    \I__2282\ : ClkMux
    port map (
            O => \N__10214\,
            I => \N__10095\
        );

    \I__2281\ : ClkMux
    port map (
            O => \N__10213\,
            I => \N__10095\
        );

    \I__2280\ : ClkMux
    port map (
            O => \N__10212\,
            I => \N__10095\
        );

    \I__2279\ : ClkMux
    port map (
            O => \N__10211\,
            I => \N__10095\
        );

    \I__2278\ : ClkMux
    port map (
            O => \N__10210\,
            I => \N__10095\
        );

    \I__2277\ : ClkMux
    port map (
            O => \N__10209\,
            I => \N__10095\
        );

    \I__2276\ : ClkMux
    port map (
            O => \N__10208\,
            I => \N__10095\
        );

    \I__2275\ : ClkMux
    port map (
            O => \N__10207\,
            I => \N__10095\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__10206\,
            I => \N__10095\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__10205\,
            I => \N__10095\
        );

    \I__2272\ : ClkMux
    port map (
            O => \N__10204\,
            I => \N__10095\
        );

    \I__2271\ : ClkMux
    port map (
            O => \N__10203\,
            I => \N__10095\
        );

    \I__2270\ : ClkMux
    port map (
            O => \N__10202\,
            I => \N__10095\
        );

    \I__2269\ : ClkMux
    port map (
            O => \N__10201\,
            I => \N__10095\
        );

    \I__2268\ : ClkMux
    port map (
            O => \N__10200\,
            I => \N__10095\
        );

    \I__2267\ : ClkMux
    port map (
            O => \N__10199\,
            I => \N__10095\
        );

    \I__2266\ : ClkMux
    port map (
            O => \N__10198\,
            I => \N__10095\
        );

    \I__2265\ : ClkMux
    port map (
            O => \N__10197\,
            I => \N__10095\
        );

    \I__2264\ : ClkMux
    port map (
            O => \N__10196\,
            I => \N__10095\
        );

    \I__2263\ : ClkMux
    port map (
            O => \N__10195\,
            I => \N__10095\
        );

    \I__2262\ : ClkMux
    port map (
            O => \N__10194\,
            I => \N__10095\
        );

    \I__2261\ : ClkMux
    port map (
            O => \N__10193\,
            I => \N__10095\
        );

    \I__2260\ : ClkMux
    port map (
            O => \N__10192\,
            I => \N__10095\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__10191\,
            I => \N__10095\
        );

    \I__2258\ : Glb2LocalMux
    port map (
            O => \N__10188\,
            I => \N__10095\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__10187\,
            I => \N__10095\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__10186\,
            I => \N__10095\
        );

    \I__2255\ : GlobalMux
    port map (
            O => \N__10095\,
            I => \CLK80_PLL\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10089\,
            I => \U712_BYTE_ENABLE.N_467\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__10086\,
            I => \U712_BYTE_ENABLE.N_455_cascade_\
        );

    \I__2251\ : IoInMux
    port map (
            O => \N__10083\,
            I => \N__10080\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10077\
        );

    \I__2249\ : IoSpan4Mux
    port map (
            O => \N__10077\,
            I => \N__10074\
        );

    \I__2248\ : IoSpan4Mux
    port map (
            O => \N__10074\,
            I => \N__10071\
        );

    \I__2247\ : Span4Mux_s2_v
    port map (
            O => \N__10071\,
            I => \N__10068\
        );

    \I__2246\ : Sp12to4
    port map (
            O => \N__10068\,
            I => \N__10065\
        );

    \I__2245\ : Span12Mux_v
    port map (
            O => \N__10065\,
            I => \N__10062\
        );

    \I__2244\ : Odrv12
    port map (
            O => \N__10062\,
            I => \N_38_i\
        );

    \I__2243\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10056\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__10053\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10046\
        );

    \I__2239\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10043\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__10046\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__10043\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10034\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10031\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10034\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10031\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10023\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10020\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__10020\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10014\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__10011\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__10011\,
            I => \N__10005\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10010\,
            I => \N__10000\
        );

    \I__2225\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10000\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10008\,
            I => \N__9997\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__10005\,
            I => \N__9989\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10000\,
            I => \N__9989\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9986\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__9989\,
            I => \N__9983\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9986\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__9983\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2216\ : IoInMux
    port map (
            O => \N__9978\,
            I => \N__9975\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__2214\ : IoSpan4Mux
    port map (
            O => \N__9972\,
            I => \N__9969\
        );

    \I__2213\ : Sp12to4
    port map (
            O => \N__9969\,
            I => \N__9966\
        );

    \I__2212\ : Span12Mux_s9_v
    port map (
            O => \N__9966\,
            I => \N__9963\
        );

    \I__2211\ : Span12Mux_h
    port map (
            O => \N__9963\,
            I => \N__9960\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__9960\,
            I => \WEn_c\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9952\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9949\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9945\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9940\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9949\,
            I => \N__9940\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9937\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9945\,
            I => \N__9934\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__9940\,
            I => \N__9931\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__9934\,
            I => \N__9925\
        );

    \I__2199\ : Span4Mux_h
    port map (
            O => \N__9931\,
            I => \N__9920\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__9928\,
            I => \N__9920\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__9925\,
            I => \N__9917\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__9920\,
            I => \N__9914\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__9917\,
            I => \N__9909\
        );

    \I__2194\ : Sp12to4
    port map (
            O => \N__9914\,
            I => \N__9909\
        );

    \I__2193\ : Span12Mux_h
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__2192\ : Odrv12
    port map (
            O => \N__9906\,
            I => \DRA_c_4\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__9891\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9884\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9881\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9884\,
            I => \N__9875\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9881\,
            I => \N__9875\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9872\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__9875\,
            I => \N__9868\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9865\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9862\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__9868\,
            I => \N__9859\
        );

    \I__2177\ : Sp12to4
    port map (
            O => \N__9865\,
            I => \N__9854\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9862\,
            I => \N__9854\
        );

    \I__2175\ : Sp12to4
    port map (
            O => \N__9859\,
            I => \N__9849\
        );

    \I__2174\ : Span12Mux_v
    port map (
            O => \N__9854\,
            I => \N__9849\
        );

    \I__2173\ : Span12Mux_h
    port map (
            O => \N__9849\,
            I => \N__9846\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__9846\,
            I => \DRA_c_6\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9840\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9831\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9828\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9825\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__9834\,
            I => \N__9820\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9831\,
            I => \N__9820\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9828\,
            I => \N__9815\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9825\,
            I => \N__9815\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9820\,
            I => \N__9812\
        );

    \I__2161\ : Span12Mux_v
    port map (
            O => \N__9815\,
            I => \N__9807\
        );

    \I__2160\ : Sp12to4
    port map (
            O => \N__9812\,
            I => \N__9807\
        );

    \I__2159\ : Span12Mux_h
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__2158\ : Odrv12
    port map (
            O => \N__9804\,
            I => \DRA_c_5\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__9801\,
            I => \N__9798\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9792\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__9792\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9784\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9779\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9779\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9774\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9774\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__9774\,
            I => \N__9770\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9767\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__9770\,
            I => \N__9764\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9761\
        );

    \I__2144\ : Sp12to4
    port map (
            O => \N__9764\,
            I => \N__9756\
        );

    \I__2143\ : Span12Mux_v
    port map (
            O => \N__9761\,
            I => \N__9756\
        );

    \I__2142\ : Span12Mux_h
    port map (
            O => \N__9756\,
            I => \N__9753\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__9753\,
            I => \DRA_c_3\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9746\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9743\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9746\,
            I => \N__9737\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9734\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9737\,
            I => \N__9729\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9729\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__9729\,
            I => \N__9725\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9722\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__9725\,
            I => \N__9719\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9716\
        );

    \I__2129\ : Sp12to4
    port map (
            O => \N__9719\,
            I => \N__9711\
        );

    \I__2128\ : Span12Mux_v
    port map (
            O => \N__9716\,
            I => \N__9711\
        );

    \I__2127\ : Span12Mux_h
    port map (
            O => \N__9711\,
            I => \N__9708\
        );

    \I__2126\ : Odrv12
    port map (
            O => \N__9708\,
            I => \DRA_c_2\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9702\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9702\,
            I => \N__9699\
        );

    \I__2123\ : Span12Mux_v
    port map (
            O => \N__9699\,
            I => \N__9696\
        );

    \I__2122\ : Odrv12
    port map (
            O => \N__9696\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__9687\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9681\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9675\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9672\,
            I => \bfn_13_12_0_\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9669\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9666\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9663\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9660\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9657\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9654\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9651\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9645\,
            I => \N__9641\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9638\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__9641\,
            I => \N__9635\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9638\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__9635\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__2100\ : ClkMux
    port map (
            O => \N__9630\,
            I => \N__9606\
        );

    \I__2099\ : ClkMux
    port map (
            O => \N__9629\,
            I => \N__9606\
        );

    \I__2098\ : ClkMux
    port map (
            O => \N__9628\,
            I => \N__9606\
        );

    \I__2097\ : ClkMux
    port map (
            O => \N__9627\,
            I => \N__9606\
        );

    \I__2096\ : ClkMux
    port map (
            O => \N__9626\,
            I => \N__9606\
        );

    \I__2095\ : ClkMux
    port map (
            O => \N__9625\,
            I => \N__9606\
        );

    \I__2094\ : ClkMux
    port map (
            O => \N__9624\,
            I => \N__9606\
        );

    \I__2093\ : ClkMux
    port map (
            O => \N__9623\,
            I => \N__9606\
        );

    \I__2092\ : GlobalMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__2091\ : gio2CtrlBuf
    port map (
            O => \N__9603\,
            I => \C1_c_g\
        );

    \I__2090\ : SRMux
    port map (
            O => \N__9600\,
            I => \N__9597\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9594\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__9594\,
            I => \N__9591\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__9591\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9584\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9581\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9584\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9581\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9572\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9569\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9572\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9569\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__9564\,
            I => \N__9560\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9557\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9554\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9545\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9542\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9545\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9542\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9534\,
            I => \U712_REG_SM.N_351\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__9531\,
            I => \N__9528\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__9522\,
            I => \N__9518\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9515\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__9518\,
            I => \U712_REG_SM.N_435\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9515\,
            I => \U712_REG_SM.N_435\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9507\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9503\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9497\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__9503\,
            I => \N__9494\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9491\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9486\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9486\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9497\,
            I => \U712_REG_SM.N_345\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__9494\,
            I => \U712_REG_SM.N_345\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9491\,
            I => \U712_REG_SM.N_345\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9486\,
            I => \U712_REG_SM.N_345\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9474\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9474\,
            I => \N__9469\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9465\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9462\
        );

    \I__2045\ : Span4Mux_h
    port map (
            O => \N__9469\,
            I => \N__9459\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9456\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9465\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9462\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9459\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9456\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9440\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__9446\,
            I => \N__9437\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9433\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9430\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \N__9427\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9440\,
            I => \N__9424\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9419\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9419\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9433\,
            I => \N__9416\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9430\,
            I => \N__9413\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9406\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__9424\,
            I => \N__9403\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9396\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__9416\,
            I => \N__9396\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__9413\,
            I => \N__9396\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9391\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9391\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9386\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9386\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9406\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__9403\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__9396\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9391\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9386\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2015\ : IoInMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9369\
        );

    \I__2013\ : Span4Mux_s1_v
    port map (
            O => \N__9369\,
            I => \N__9366\
        );

    \I__2012\ : Sp12to4
    port map (
            O => \N__9366\,
            I => \N__9363\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9360\,
            I => \ASn_c\
        );

    \I__2009\ : CEMux
    port map (
            O => \N__9357\,
            I => \N__9354\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9351\,
            I => \U712_REG_SM.N_131_0\
        );

    \I__2006\ : IoInMux
    port map (
            O => \N__9348\,
            I => \N__9345\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9345\,
            I => \N__9342\
        );

    \I__2004\ : Odrv12
    port map (
            O => \N__9342\,
            I => \RESETn_c_i\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9333\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9333\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9333\,
            I => \N__9330\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__9327\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9321\,
            I => \N__9318\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__9318\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9311\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9308\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9311\,
            I => \N__9305\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9308\,
            I => \N__9302\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__9305\,
            I => \N__9295\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__9302\,
            I => \N__9295\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9290\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9290\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__9295\,
            I => \N__9287\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9290\,
            I => \N__9284\
        );

    \I__1985\ : Sp12to4
    port map (
            O => \N__9287\,
            I => \N__9281\
        );

    \I__1984\ : Span12Mux_h
    port map (
            O => \N__9284\,
            I => \N__9278\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__9281\,
            I => \DRA_c_8\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__9278\,
            I => \DRA_c_8\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9268\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9265\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9262\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9259\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9254\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9262\,
            I => \N__9254\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__9259\,
            I => \N__9250\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9247\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9244\
        );

    \I__1972\ : Sp12to4
    port map (
            O => \N__9250\,
            I => \N__9237\
        );

    \I__1971\ : Sp12to4
    port map (
            O => \N__9247\,
            I => \N__9237\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9244\,
            I => \N__9237\
        );

    \I__1969\ : Span12Mux_h
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__1968\ : Odrv12
    port map (
            O => \N__9234\,
            I => \DRA_c_7\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9218\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9215\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9218\,
            I => \N__9212\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9215\,
            I => \N__9209\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__9212\,
            I => \N__9204\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__9209\,
            I => \N__9204\
        );

    \I__1958\ : Sp12to4
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__1956\ : Span12Mux_v
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__9195\,
            I => \DRA_c_0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9184\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9181\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9178\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__9184\,
            I => \N__9175\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9181\,
            I => \N__9172\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__9178\,
            I => \N__9169\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__9175\,
            I => \N__9165\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__9172\,
            I => \N__9160\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__9169\,
            I => \N__9160\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9157\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__9165\,
            I => \N__9154\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__9160\,
            I => \N__9149\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__9157\,
            I => \N__9149\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__9154\,
            I => \N__9146\
        );

    \I__1939\ : Sp12to4
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__1938\ : Sp12to4
    port map (
            O => \N__9146\,
            I => \N__9138\
        );

    \I__1937\ : Span12Mux_v
    port map (
            O => \N__9143\,
            I => \N__9138\
        );

    \I__1936\ : Span12Mux_h
    port map (
            O => \N__9138\,
            I => \N__9135\
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__9135\,
            I => \DRA_c_1\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__1932\ : Odrv12
    port map (
            O => \N__9126\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__9114\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9105\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9105\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9105\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__1924\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9098\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9095\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9098\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__9095\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__9090\,
            I => \N__9086\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9083\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9080\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__9083\,
            I => \DBR_SYNC_i_1\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9080\,
            I => \DBR_SYNC_i_1\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9072\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9072\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9065\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9062\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__9065\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9062\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9051\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9051\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9048\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9041\
        );

    \I__1904\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9038\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__9041\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9038\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__9033\,
            I => \N__9030\
        );

    \I__1900\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9027\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9027\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__1898\ : InMux
    port map (
            O => \N__9024\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9021\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__1896\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__9015\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__9012\,
            I => \N__9007\
        );

    \I__1893\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8997\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8997\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8997\
        );

    \I__1890\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8994\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8991\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8988\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8985\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8980\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8975\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8975\
        );

    \I__1883\ : Span4Mux_h
    port map (
            O => \N__8985\,
            I => \N__8971\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8968\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8965\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__8980\,
            I => \N__8960\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__8975\,
            I => \N__8960\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8957\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__8971\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8968\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8965\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__8960\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8957\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8942\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__8945\,
            I => \N__8938\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8935\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8928\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8925\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__8935\,
            I => \N__8922\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8913\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8913\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8913\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8913\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8910\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8925\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__8922\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8913\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8910\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8898\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8892\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8892\,
            I => \N__8889\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__8889\,
            I => \N__8885\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8882\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8885\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8882\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__8871\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__8862\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8856\,
            I => \N__8853\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__8853\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8847\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8837\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8840\,
            I => \N__8834\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__8837\,
            I => \N__8831\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8828\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__8831\,
            I => \N__8823\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8823\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__8823\,
            I => \N__8818\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8815\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8812\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__8818\,
            I => \REG_CYCLEm\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8815\,
            I => \REG_CYCLEm\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8812\,
            I => \REG_CYCLEm\
        );

    \I__1825\ : IoInMux
    port map (
            O => \N__8805\,
            I => \N__8802\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8802\,
            I => \N__8799\
        );

    \I__1823\ : Span4Mux_s2_v
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__8796\,
            I => \N__8793\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__1819\ : Span12Mux_h
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__8784\,
            I => \N_196_i\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8778\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8772\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8772\,
            I => \N__8769\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__8766\,
            I => \U712_CHIP_RAM.N_492\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8758\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8755\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8752\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8758\,
            I => \U712_REG_SM.N_131\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8755\,
            I => \U712_REG_SM.N_131\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8752\,
            I => \U712_REG_SM.N_131\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8742\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_7\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8732\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8729\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__8732\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8729\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8721\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_6\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8709\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8706\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8703\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \N__8700\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__8709\,
            I => \N__8694\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8706\,
            I => \N__8694\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8703\,
            I => \N__8691\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8688\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8685\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__8694\,
            I => \N__8680\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__8691\,
            I => \N__8680\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8688\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8685\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__8680\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1781\ : IoInMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1779\ : Span4Mux_s3_v
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__1777\ : Sp12to4
    port map (
            O => \N__8661\,
            I => \N__8658\
        );

    \I__1776\ : Span12Mux_h
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__8655\,
            I => \CRCSn_c\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1772\ : Span4Mux_h
    port map (
            O => \N__8646\,
            I => \N__8643\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__8643\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8637\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8631\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__8622\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__8613\,
            I => \N__8610\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__8610\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8601\
        );

    \I__1757\ : Span4Mux_h
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__8598\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8592\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8592\,
            I => \N__8586\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8583\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8580\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8577\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__8586\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8583\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8580\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8577\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8565\,
            I => \U712_REG_SM.N_365\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8559\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_4\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8553\,
            I => \U712_REG_SM.N_588\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8547\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8540\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8537\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8540\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8537\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__8532\,
            I => \N__8529\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8521\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8518\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8510\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__8521\,
            I => \N__8505\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8505\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8498\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8498\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8498\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8493\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8493\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__8505\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8498\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8493\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__8484\,
            I => \N__8480\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8476\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8471\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8468\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8476\,
            I => \N__8465\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8460\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8460\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8471\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8468\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8465\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8460\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__8451\,
            I => \U712_REG_SM.N_395_cascade_\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__8448\,
            I => \U712_REG_SM.N_439_cascade_\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8442\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8442\,
            I => \U712_REG_SM.REG_CYCLE_5_iv_0_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8436\,
            I => \U712_REG_SM.N_395\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8419\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8419\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8416\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8424\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8419\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8416\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1693\ : IoInMux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8403\
        );

    \I__1691\ : Span4Mux_s2_v
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__8400\,
            I => \N__8396\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8393\
        );

    \I__1688\ : Span4Mux_h
    port map (
            O => \N__8396\,
            I => \N__8390\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8393\,
            I => \N__8387\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__8390\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1685\ : Odrv12
    port map (
            O => \N__8387\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__8382\,
            I => \N__8375\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8370\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8370\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \N__8366\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8361\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8354\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8351\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8346\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8346\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8343\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8330\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8325\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8325\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8318\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8318\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8318\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8311\
        );

    \I__1667\ : Span4Mux_h
    port map (
            O => \N__8351\,
            I => \N__8311\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8346\,
            I => \N__8311\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8308\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8301\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8301\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8301\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8296\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8296\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8293\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8290\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8287\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8282\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8282\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8330\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__8325\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8318\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__8311\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__8308\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8301\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8296\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8293\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8290\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8287\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__8282\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8256\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8256\,
            I => \N__8253\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__8253\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1640\ : IoInMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1638\ : Span4Mux_s2_v
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1637\ : Sp12to4
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1636\ : Span12Mux_h
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1635\ : Span12Mux_v
    port map (
            O => \N__8235\,
            I => \N__8231\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8228\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__8231\,
            I => \PRnW_c\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8228\,
            I => \PRnW_c\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8215\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8212\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8209\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__8215\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8212\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8209\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8194\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8189\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8186\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__8194\,
            I => \N__8183\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8178\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8178\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8189\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__8183\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8178\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__8169\,
            I => \U712_REG_SM.N_351_cascade_\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8162\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8159\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8156\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8159\,
            I => \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__8156\,
            I => \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8142\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8142\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8142\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8142\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8135\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8132\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8127\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8132\,
            I => \N__8127\
        );

    \I__1599\ : Span12Mux_h
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1598\ : Span12Mux_v
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__8121\,
            I => \TSn_c\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8111\
        );

    \I__1594\ : IoInMux
    port map (
            O => \N__8114\,
            I => \N__8108\
        );

    \I__1593\ : Span12Mux_h
    port map (
            O => \N__8111\,
            I => \N__8105\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8102\
        );

    \I__1591\ : Span12Mux_v
    port map (
            O => \N__8105\,
            I => \N__8099\
        );

    \I__1590\ : IoSpan4Mux
    port map (
            O => \N__8102\,
            I => \N__8096\
        );

    \I__1589\ : Odrv12
    port map (
            O => \N__8099\,
            I => \RAMENn_c\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__8096\,
            I => \RAMENn_c\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__8091\,
            I => \U712_CHIP_RAM.N_448_cascade_\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8083\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8078\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8078\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8083\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8078\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8070\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__8061\,
            I => \U712_CHIP_RAM.N_450\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1574\ : Sp12to4
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1573\ : Span12Mux_v
    port map (
            O => \N__8049\,
            I => \N__8046\
        );

    \I__1572\ : Span12Mux_h
    port map (
            O => \N__8046\,
            I => \N__8043\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__8043\,
            I => \A_c_15\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8037\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__8037\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__8034\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__8028\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1565\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__8019\
        );

    \I__1563\ : Sp12to4
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1562\ : Span12Mux_v
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1561\ : Span12Mux_h
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__8010\,
            I => \A_c_13\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7995\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7990\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7990\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7986\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7974\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7974\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7974\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7995\,
            I => \N__7969\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7990\,
            I => \N__7969\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7960\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7950\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7947\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7942\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7942\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7939\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7936\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7974\,
            I => \N__7931\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__7969\,
            I => \N__7931\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7926\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7926\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7921\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7921\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7910\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7910\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7910\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7910\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7910\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7899\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7899\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7899\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7899\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7899\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7950\,
            I => \N__7892\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7947\,
            I => \N__7892\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7942\,
            I => \N__7892\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7939\,
            I => \N__7889\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7936\,
            I => \N__7884\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7931\,
            I => \N__7884\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7879\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7879\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7910\,
            I => \N__7874\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7899\,
            I => \N__7874\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__7892\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__7889\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__7884\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1513\ : Odrv12
    port map (
            O => \N__7879\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__7874\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7860\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7851\
        );

    \I__1507\ : Span4Mux_v
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1506\ : Sp12to4
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1505\ : Span12Mux_h
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__7842\,
            I => \A_c_6\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7836\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1501\ : CEMux
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7826\
        );

    \I__1499\ : CEMux
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__7826\,
            I => \N__7820\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7823\,
            I => \N__7817\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7820\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1495\ : Odrv12
    port map (
            O => \N__7817\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1492\ : Span4Mux_h
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1490\ : Sp12to4
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1489\ : Span12Mux_h
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__7794\,
            I => \A_c_20\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7786\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7781\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7781\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7786\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7781\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7773\,
            I => \N__7769\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7766\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__7769\,
            I => \N__7763\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7766\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7763\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7754\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7751\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7748\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7745\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__7748\,
            I => \N__7742\
        );

    \I__1471\ : Odrv12
    port map (
            O => \N__7745\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__7742\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7733\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7730\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7733\,
            I => \N__7724\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7730\,
            I => \N__7724\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7719\
        );

    \I__1464\ : Span4Mux_h
    port map (
            O => \N__7724\,
            I => \N__7716\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7713\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7710\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7719\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__7716\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7713\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7710\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__7695\,
            I => \N__7691\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7688\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7691\,
            I => \U712_CHIP_RAM.N_461\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7688\,
            I => \U712_CHIP_RAM.N_461\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__7683\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\
        );

    \I__1450\ : IoInMux
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1448\ : Span4Mux_s3_v
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1447\ : Sp12to4
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1446\ : Span12Mux_h
    port map (
            O => \N__7668\,
            I => \N__7664\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7661\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__7664\,
            I => \LATCH_CLK_c\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7661\,
            I => \LATCH_CLK_c\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7653\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7653\,
            I => \U712_REG_SM.N_357\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7650\,
            I => \N__7646\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7643\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7640\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7643\,
            I => \U712_REG_SM.N_353\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7640\,
            I => \U712_REG_SM.N_353\
        );

    \I__1435\ : IoInMux
    port map (
            O => \N__7635\,
            I => \N__7632\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1433\ : Span4Mux_s1_v
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1432\ : Sp12to4
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1431\ : Span12Mux_h
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__7620\,
            I => \CASn_c\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7613\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__7616\,
            I => \N__7607\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7613\,
            I => \N__7604\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7601\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7598\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7593\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7593\
        );

    \I__1422\ : Span4Mux_v
    port map (
            O => \N__7604\,
            I => \N__7583\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7583\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7583\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7583\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7580\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__7583\,
            I => \N__7577\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7580\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__7577\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1414\ : IoInMux
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1412\ : Span4Mux_s2_v
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1411\ : Span4Mux_h
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1410\ : Sp12to4
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1409\ : Span12Mux_v
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1408\ : Odrv12
    port map (
            O => \N__7554\,
            I => \RASn_c\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__7551\,
            I => \N__7548\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7541\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7538\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__7541\,
            I => \N__7535\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7532\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__7535\,
            I => \N__7527\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__7532\,
            I => \N__7527\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__7527\,
            I => \DBRn_c_i\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7520\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7517\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7520\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7517\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7509\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1390\ : Span4Mux_h
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__7497\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1388\ : IoInMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1386\ : IoSpan4Mux
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1385\ : IoSpan4Mux
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1384\ : Span4Mux_s3_h
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__7479\,
            I => \N__7476\
        );

    \I__1382\ : Sp12to4
    port map (
            O => \N__7476\,
            I => \N__7472\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1380\ : Span12Mux_h
    port map (
            O => \N__7472\,
            I => \N__7464\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7469\,
            I => \N__7464\
        );

    \I__1378\ : Span12Mux_h
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1377\ : Odrv12
    port map (
            O => \N__7461\,
            I => \C3_c\
        );

    \I__1376\ : IoInMux
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7455\,
            I => \N__7451\
        );

    \I__1374\ : IoInMux
    port map (
            O => \N__7454\,
            I => \N__7448\
        );

    \I__1373\ : IoSpan4Mux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7448\,
            I => \N__7442\
        );

    \I__1371\ : Span4Mux_s1_v
    port map (
            O => \N__7445\,
            I => \N__7439\
        );

    \I__1370\ : Span4Mux_s1_v
    port map (
            O => \N__7442\,
            I => \N__7436\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__7439\,
            I => \N__7433\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__7436\,
            I => \N__7430\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__7433\,
            I => \N__7427\
        );

    \I__1366\ : Sp12to4
    port map (
            O => \N__7430\,
            I => \N__7424\
        );

    \I__1365\ : Span12Mux_h
    port map (
            O => \N__7427\,
            I => \N__7418\
        );

    \I__1364\ : Span12Mux_h
    port map (
            O => \N__7424\,
            I => \N__7418\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7415\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__7418\,
            I => \BLSn_c\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7415\,
            I => \BLSn_c\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7407\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7407\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__7404\,
            I => \U712_REG_SM.N_345_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7396\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7391\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7391\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7396\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7391\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7383\,
            I => \U712_REG_SM.N_396\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__7380\,
            I => \U712_REG_SM.N_435_cascade_\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7371\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7371\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7371\,
            I => \U712_REG_SM.N_352\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7362\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7362\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7362\,
            I => \U712_CHIP_RAM.N_500\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__7359\,
            I => \N__7350\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7346\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7343\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7340\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7337\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7334\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7331\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7350\,
            I => \N__7326\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7326\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7346\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7343\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7340\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7337\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7334\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7331\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7326\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.N_500_cascade_\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7300\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7293\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7293\
        );

    \I__1322\ : Span4Mux_h
    port map (
            O => \N__7300\,
            I => \N__7290\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7287\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7284\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7293\,
            I => \U712_CHIP_RAM.N_514\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__7290\,
            I => \U712_CHIP_RAM.N_514\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7287\,
            I => \U712_CHIP_RAM.N_514\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7284\,
            I => \U712_CHIP_RAM.N_514\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7275\,
            I => \N__7270\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7267\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7264\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7261\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7267\,
            I => \N__7256\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7264\,
            I => \N__7246\
        );

    \I__1309\ : Span4Mux_h
    port map (
            O => \N__7261\,
            I => \N__7246\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7241\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7241\
        );

    \I__1306\ : Span4Mux_h
    port map (
            O => \N__7256\,
            I => \N__7238\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7233\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7233\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7226\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7226\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7226\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__7246\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7241\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__7238\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7233\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7226\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7211\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7208\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7203\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7203\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__7203\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7197\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7194\
        );

    \I__1288\ : Span4Mux_h
    port map (
            O => \N__7194\,
            I => \N__7190\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7187\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__7190\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7187\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7179\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7176\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__7176\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7168\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__7172\,
            I => \N__7165\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7160\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7168\,
            I => \N__7154\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7151\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7148\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__7163\,
            I => \N__7145\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7160\,
            I => \N__7142\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7139\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__7158\,
            I => \N__7135\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__7157\,
            I => \N__7131\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__7154\,
            I => \N__7125\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7125\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7148\,
            I => \N__7120\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7117\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__7142\,
            I => \N__7112\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7139\,
            I => \N__7112\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7109\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7106\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7101\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7101\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7098\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__7125\,
            I => \N__7095\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7090\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7090\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__7120\,
            I => \N__7087\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__7117\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__7112\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7109\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7106\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7101\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7098\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__7095\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__7090\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__7087\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__7068\,
            I => \N__7062\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7059\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__7066\,
            I => \N__7055\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7050\
        );

    \I__1242\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7050\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7046\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__7058\,
            I => \N__7043\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7039\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7050\,
            I => \N__7036\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__7049\,
            I => \N__7031\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__7046\,
            I => \N__7026\
        );

    \I__1235\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7023\
        );

    \I__1234\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7020\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7039\,
            I => \N__7015\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__7036\,
            I => \N__7015\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7012\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7009\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7004\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7004\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7001\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__7026\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7023\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7020\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__7015\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__7012\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7009\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__7004\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__7001\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6978\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6978\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6978\,
            I => \CPU_TACKm\
        );

    \I__1215\ : CEMux
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__6969\,
            I => \U712_CHIP_RAM.N_248_0\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6962\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6962\,
            I => \N__6953\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6949\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__6953\,
            I => \N__6946\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6943\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6949\,
            I => \N__6939\
        );

    \I__1204\ : Span4Mux_v
    port map (
            O => \N__6946\,
            I => \N__6934\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6934\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6942\,
            I => \N__6931\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__6939\,
            I => \N__6926\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__6934\,
            I => \N__6926\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6923\
        );

    \I__1198\ : Sp12to4
    port map (
            O => \N__6926\,
            I => \N__6918\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6918\
        );

    \I__1196\ : Span12Mux_h
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1195\ : Odrv12
    port map (
            O => \N__6915\,
            I => \RnW_c\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6909\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6898\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6893\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6893\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6898\,
            I => \REG_TACK\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6893\,
            I => \REG_TACK\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6884\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6881\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6878\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6881\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6878\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__6873\,
            I => \U712_CHIP_RAM.N_514_cascade_\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6866\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6863\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6860\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6863\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6860\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6851\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6848\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6851\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6848\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__6843\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\
        );

    \I__1170\ : CEMux
    port map (
            O => \N__6840\,
            I => \N__6837\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__6831\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6820\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6817\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6813\
        );

    \I__1162\ : Span4Mux_h
    port map (
            O => \N__6820\,
            I => \N__6808\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6805\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6802\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6813\,
            I => \N__6799\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6794\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6794\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__6808\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__1155\ : Odrv12
    port map (
            O => \N__6805\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6802\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6799\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6794\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6780\,
            I => \N__6777\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6777\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6767\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6767\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6763\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6760\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6757\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6754\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__6760\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6757\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__6754\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6747\,
            I => \U712_CHIP_RAM.N_481_cascade_\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6744\,
            I => \U712_REG_SM.N_428_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__6732\,
            I => \N__6729\
        );

    \I__1133\ : Sp12to4
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1132\ : Span12Mux_v
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__6723\,
            I => \REGSPACEn_c\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1128\ : Span12Mux_v
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1127\ : Span12Mux_h
    port map (
            O => \N__6711\,
            I => \N__6708\
        );

    \I__1126\ : Odrv12
    port map (
            O => \N__6708\,
            I => \A_c_3\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6696\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6696\,
            I => \N__6693\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1120\ : Sp12to4
    port map (
            O => \N__6690\,
            I => \N__6687\
        );

    \I__1119\ : Span12Mux_h
    port map (
            O => \N__6687\,
            I => \N__6684\
        );

    \I__1118\ : Odrv12
    port map (
            O => \N__6684\,
            I => \A_c_4\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1115\ : Span4Mux_h
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__6672\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1110\ : Span4Mux_h
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1109\ : Sp12to4
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1108\ : Odrv12
    port map (
            O => \N__6654\,
            I => \A_c_7\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6648\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6642\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6642\,
            I => \N__6639\
        );

    \I__1103\ : Span12Mux_h
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__6636\,
            I => \A_c_8\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1098\ : Sp12to4
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1097\ : Span12Mux_h
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6618\,
            I => \A_c_5\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6612\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6606\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6603\
        );

    \I__1091\ : Span12Mux_v
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__1090\ : Span12Mux_v
    port map (
            O => \N__6600\,
            I => \N__6597\
        );

    \I__1089\ : Span12Mux_h
    port map (
            O => \N__6597\,
            I => \N__6594\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__6594\,
            I => \A_c_18\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6588\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6588\,
            I => \N__6585\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__6585\,
            I => \N__6582\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__6582\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__6579\,
            I => \N__6576\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6568\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6568\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6565\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6562\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6568\,
            I => \N__6544\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6565\,
            I => \N__6539\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6539\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6532\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6560\,
            I => \N__6532\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6532\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6527\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6527\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6520\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6520\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6520\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6513\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6513\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6513\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6510\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6505\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6505\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6502\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__6544\,
            I => \N__6499\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6532\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6520\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6505\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6502\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__6499\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6477\,
            I => \N__6468\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6461\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6456\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6456\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6451\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6448\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6445\
        );

    \I__1042\ : Span4Mux_h
    port map (
            O => \N__6468\,
            I => \N__6442\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6435\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6435\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6435\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6432\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6461\,
            I => \N__6427\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6427\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6422\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6422\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6451\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6448\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6445\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__6442\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6435\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6432\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__6427\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6402\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1021\ : Span4Mux_v
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1019\ : Span12Mux_h
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1018\ : Span12Mux_v
    port map (
            O => \N__6384\,
            I => \N__6381\
        );

    \I__1017\ : Odrv12
    port map (
            O => \N__6381\,
            I => \A_c_19\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6375\,
            I => \N__6372\
        );

    \I__1014\ : Span4Mux_s3_h
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1013\ : Sp12to4
    port map (
            O => \N__6369\,
            I => \N__6366\
        );

    \I__1012\ : Span12Mux_v
    port map (
            O => \N__6366\,
            I => \N__6363\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__6360\,
            I => \CMA_c_9\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6353\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6350\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6353\,
            I => \N__6342\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6339\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6328\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6328\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6328\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6328\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6328\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__6342\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6339\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6328\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__6318\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\
        );

    \I__995\ : CEMux
    port map (
            O => \N__6315\,
            I => \N__6311\
        );

    \I__994\ : CEMux
    port map (
            O => \N__6314\,
            I => \N__6308\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6303\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6300\
        );

    \I__991\ : CEMux
    port map (
            O => \N__6307\,
            I => \N__6297\
        );

    \I__990\ : CEMux
    port map (
            O => \N__6306\,
            I => \N__6294\
        );

    \I__989\ : Span4Mux_h
    port map (
            O => \N__6303\,
            I => \N__6289\
        );

    \I__988\ : Span4Mux_v
    port map (
            O => \N__6300\,
            I => \N__6289\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6297\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6294\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__6289\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__984\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6279\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__982\ : Span12Mux_v
    port map (
            O => \N__6276\,
            I => \N__6273\
        );

    \I__981\ : Span12Mux_h
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__980\ : Odrv12
    port map (
            O => \N__6270\,
            I => \A_c_12\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__6267\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__978\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6261\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6261\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__976\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6255\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6252\
        );

    \I__974\ : Span4Mux_h
    port map (
            O => \N__6252\,
            I => \N__6249\
        );

    \I__973\ : Sp12to4
    port map (
            O => \N__6249\,
            I => \N__6246\
        );

    \I__972\ : Span12Mux_v
    port map (
            O => \N__6246\,
            I => \N__6243\
        );

    \I__971\ : Odrv12
    port map (
            O => \N__6243\,
            I => \A_c_2\
        );

    \I__970\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6237\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6237\,
            I => \N__6234\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__6234\,
            I => \N__6231\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__6231\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__966\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6225\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__964\ : Span12Mux_v
    port map (
            O => \N__6222\,
            I => \N__6219\
        );

    \I__963\ : Span12Mux_h
    port map (
            O => \N__6219\,
            I => \N__6216\
        );

    \I__962\ : Odrv12
    port map (
            O => \N__6216\,
            I => \A_c_16\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6213\,
            I => \N__6210\
        );

    \I__960\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6207\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__958\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__6198\,
            I => \N__6195\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__6195\,
            I => \N__6192\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__6189\,
            I => \N__6186\
        );

    \I__952\ : Sp12to4
    port map (
            O => \N__6186\,
            I => \N__6183\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__6183\,
            I => \A_c_17\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__6180\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__949\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6171\
        );

    \I__947\ : Span12Mux_v
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__946\ : Span12Mux_h
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__945\ : Odrv12
    port map (
            O => \N__6165\,
            I => \A_c_14\
        );

    \I__944\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6159\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__6159\,
            I => \U712_CHIP_RAM.N_383\
        );

    \I__942\ : IoInMux
    port map (
            O => \N__6156\,
            I => \N__6153\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__940\ : IoSpan4Mux
    port map (
            O => \N__6150\,
            I => \N__6147\
        );

    \I__939\ : Span4Mux_s2_v
    port map (
            O => \N__6147\,
            I => \N__6144\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__6144\,
            I => \N__6141\
        );

    \I__937\ : Span12Mux_s10_h
    port map (
            O => \N__6141\,
            I => \N__6138\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__6138\,
            I => \N__6135\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__6135\,
            I => \CMA_c_3\
        );

    \I__934\ : IoInMux
    port map (
            O => \N__6132\,
            I => \N__6129\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6129\,
            I => \N__6126\
        );

    \I__932\ : Span12Mux_s11_h
    port map (
            O => \N__6126\,
            I => \N__6123\
        );

    \I__931\ : Span12Mux_v
    port map (
            O => \N__6123\,
            I => \N__6120\
        );

    \I__930\ : Odrv12
    port map (
            O => \N__6120\,
            I => \CMA_c_4\
        );

    \I__929\ : IoInMux
    port map (
            O => \N__6117\,
            I => \N__6114\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6114\,
            I => \N__6111\
        );

    \I__927\ : IoSpan4Mux
    port map (
            O => \N__6111\,
            I => \N__6108\
        );

    \I__926\ : Span4Mux_s2_v
    port map (
            O => \N__6108\,
            I => \N__6105\
        );

    \I__925\ : Sp12to4
    port map (
            O => \N__6105\,
            I => \N__6102\
        );

    \I__924\ : Span12Mux_h
    port map (
            O => \N__6102\,
            I => \N__6099\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__922\ : Odrv12
    port map (
            O => \N__6096\,
            I => \CMA_c_6\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6090\
        );

    \I__920\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6087\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__6087\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__918\ : IoInMux
    port map (
            O => \N__6084\,
            I => \N__6081\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__916\ : Span4Mux_s2_h
    port map (
            O => \N__6078\,
            I => \N__6075\
        );

    \I__915\ : Span4Mux_h
    port map (
            O => \N__6075\,
            I => \N__6072\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__6072\,
            I => \N__6069\
        );

    \I__913\ : Span12Mux_v
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__912\ : Span12Mux_h
    port map (
            O => \N__6066\,
            I => \N__6063\
        );

    \I__911\ : Odrv12
    port map (
            O => \N__6063\,
            I => \CMA_c_7\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6060\,
            I => \N__6054\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__6059\,
            I => \N__6046\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__6058\,
            I => \N__6043\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__6057\,
            I => \N__6040\
        );

    \I__906\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6037\
        );

    \I__905\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6033\
        );

    \I__904\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6028\
        );

    \I__903\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6028\
        );

    \I__902\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6023\
        );

    \I__901\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6023\
        );

    \I__900\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6016\
        );

    \I__899\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6016\
        );

    \I__898\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6016\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6013\
        );

    \I__896\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6010\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6033\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6028\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6023\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__6016\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__6013\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__6010\,
            I => \U712_CHIP_RAM.N_343\
        );

    \I__889\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5994\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__887\ : IoInMux
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5988\,
            I => \N__5985\
        );

    \I__885\ : Span4Mux_s2_h
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__883\ : Span12Mux_v
    port map (
            O => \N__5979\,
            I => \N__5976\
        );

    \I__882\ : Span12Mux_h
    port map (
            O => \N__5976\,
            I => \N__5973\
        );

    \I__881\ : Odrv12
    port map (
            O => \N__5973\,
            I => \CMA_c_8\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5970\,
            I => \U712_REG_SM.N_352_cascade_\
        );

    \I__879\ : IoInMux
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5964\,
            I => \N__5960\
        );

    \I__877\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5957\
        );

    \I__876\ : IoSpan4Mux
    port map (
            O => \N__5960\,
            I => \N__5954\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5957\,
            I => \N__5951\
        );

    \I__874\ : IoSpan4Mux
    port map (
            O => \N__5954\,
            I => \N__5948\
        );

    \I__873\ : Span12Mux_h
    port map (
            O => \N__5951\,
            I => \N__5945\
        );

    \I__872\ : IoSpan4Mux
    port map (
            O => \N__5948\,
            I => \N__5942\
        );

    \I__871\ : Odrv12
    port map (
            O => \N__5945\,
            I => \C1_c\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5942\,
            I => \C1_c\
        );

    \I__869\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5931\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__866\ : IoInMux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__864\ : Span4Mux_s2_v
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__863\ : Span4Mux_v
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__861\ : Span12Mux_h
    port map (
            O => \N__5913\,
            I => \N__5909\
        );

    \I__860\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5906\
        );

    \I__859\ : Odrv12
    port map (
            O => \N__5909\,
            I => \UDSn_c\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5906\,
            I => \UDSn_c\
        );

    \I__857\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5898\,
            I => \U712_REG_SM.N_429\
        );

    \I__855\ : IoInMux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__853\ : Span4Mux_s3_v
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__851\ : Sp12to4
    port map (
            O => \N__5883\,
            I => \N__5879\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__5882\,
            I => \N__5876\
        );

    \I__849\ : Span12Mux_h
    port map (
            O => \N__5879\,
            I => \N__5873\
        );

    \I__848\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__847\ : Odrv12
    port map (
            O => \N__5873\,
            I => \LDSn_c\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5870\,
            I => \LDSn_c\
        );

    \I__845\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5862\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5862\,
            I => \U712_REG_SM.N_493\
        );

    \I__843\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5852\
        );

    \I__842\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5852\
        );

    \I__841\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5849\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5846\,
            I => \U712_CHIP_RAM.N_590\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.N_590\
        );

    \I__836\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5834\
        );

    \I__835\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5831\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5834\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5831\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__5826\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__5823\,
            I => \U712_CHIP_RAM.N_248_cascade_\
        );

    \I__830\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5817\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5814\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__827\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__5805\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__823\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5793\
        );

    \I__822\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5793\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5793\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__820\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5784\
        );

    \I__819\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5784\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__5781\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__5778\,
            I => \U712_CYCLE_TERM.N_358_i_cascade_\
        );

    \I__815\ : IoInMux
    port map (
            O => \N__5775\,
            I => \N__5771\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__5774\,
            I => \N__5767\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5764\
        );

    \I__812\ : IoInMux
    port map (
            O => \N__5770\,
            I => \N__5761\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5767\,
            I => \N__5758\
        );

    \I__810\ : IoSpan4Mux
    port map (
            O => \N__5764\,
            I => \N__5755\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5752\
        );

    \I__808\ : Span12Mux_s7_v
    port map (
            O => \N__5758\,
            I => \N__5749\
        );

    \I__807\ : Sp12to4
    port map (
            O => \N__5755\,
            I => \N__5746\
        );

    \I__806\ : IoSpan4Mux
    port map (
            O => \N__5752\,
            I => \N__5743\
        );

    \I__805\ : Span12Mux_h
    port map (
            O => \N__5749\,
            I => \N__5740\
        );

    \I__804\ : Span12Mux_s7_v
    port map (
            O => \N__5746\,
            I => \N__5737\
        );

    \I__803\ : Sp12to4
    port map (
            O => \N__5743\,
            I => \N__5734\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__5740\,
            I => \N__5728\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__5737\,
            I => \N__5728\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__5734\,
            I => \N__5725\
        );

    \I__799\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5722\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__5728\,
            I => \TACK_EN\
        );

    \I__797\ : Odrv12
    port map (
            O => \N__5725\,
            I => \TACK_EN\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5722\,
            I => \TACK_EN\
        );

    \I__795\ : InMux
    port map (
            O => \N__5715\,
            I => \N__5707\
        );

    \I__794\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5707\
        );

    \I__793\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5704\
        );

    \I__792\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5701\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5698\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5695\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5701\,
            I => \N__5692\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5689\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__5695\,
            I => \N__5684\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__5692\,
            I => \N__5684\
        );

    \I__785\ : Span4Mux_h
    port map (
            O => \N__5689\,
            I => \N__5681\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__5684\,
            I => \N__5678\
        );

    \I__783\ : Sp12to4
    port map (
            O => \N__5681\,
            I => \N__5673\
        );

    \I__782\ : Span12Mux_h
    port map (
            O => \N__5678\,
            I => \N__5673\
        );

    \I__781\ : Span12Mux_v
    port map (
            O => \N__5673\,
            I => \N__5670\
        );

    \I__780\ : Odrv12
    port map (
            O => \N__5670\,
            I => \CLK40_PLL_i\
        );

    \I__779\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5661\
        );

    \I__778\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5654\
        );

    \I__777\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5654\
        );

    \I__776\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5654\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5661\,
            I => \N__5651\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5654\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__5651\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__772\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5642\
        );

    \I__771\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5639\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5642\,
            I => \N__5636\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5633\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__5636\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__5633\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__766\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5624\
        );

    \I__765\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5621\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5618\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5615\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__5618\,
            I => \N__5612\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__5615\,
            I => \N__5609\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__5612\,
            I => \N__5606\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__5609\,
            I => \N__5603\
        );

    \I__758\ : Sp12to4
    port map (
            O => \N__5606\,
            I => \N__5598\
        );

    \I__757\ : Span12Mux_h
    port map (
            O => \N__5603\,
            I => \N__5598\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__5598\,
            I => \DBRn_c\
        );

    \I__755\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5586\
        );

    \I__754\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5586\
        );

    \I__753\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5586\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5586\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__751\ : IoInMux
    port map (
            O => \N__5583\,
            I => \N__5580\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__749\ : IoSpan4Mux
    port map (
            O => \N__5577\,
            I => \N__5574\
        );

    \I__748\ : IoSpan4Mux
    port map (
            O => \N__5574\,
            I => \N__5571\
        );

    \I__747\ : Sp12to4
    port map (
            O => \N__5571\,
            I => \N__5568\
        );

    \I__746\ : Span12Mux_s7_h
    port map (
            O => \N__5568\,
            I => \N__5565\
        );

    \I__745\ : Span12Mux_h
    port map (
            O => \N__5565\,
            I => \N__5562\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__5562\,
            I => \DRDDIR_c\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__5559\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\
        );

    \I__742\ : CEMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__5550\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__5547\,
            I => \N__5543\
        );

    \I__738\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5537\
        );

    \I__737\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5534\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__5542\,
            I => \N__5528\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5541\,
            I => \N__5522\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5519\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5515\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5512\
        );

    \I__731\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5507\
        );

    \I__730\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5507\
        );

    \I__729\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5503\
        );

    \I__728\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5500\
        );

    \I__727\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5497\
        );

    \I__726\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5494\
        );

    \I__725\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5485\
        );

    \I__724\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5485\
        );

    \I__723\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5485\
        );

    \I__722\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5485\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5478\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__5512\,
            I => \N__5478\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5478\
        );

    \I__718\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5475\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5503\,
            I => \N__5470\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5470\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5497\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5494\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5475\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__5470\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__5457\,
            I => \U712_CHIP_RAM.N_503_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5451\,
            I => \U712_CHIP_RAM.N_420\
        );

    \I__706\ : CEMux
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5445\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\
        );

    \I__704\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5438\
        );

    \I__703\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5435\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5432\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5435\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5432\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__699\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__5421\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5408\
        );

    \I__693\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5405\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__5408\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5405\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__689\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5390\
        );

    \I__688\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5385\
        );

    \I__687\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5382\
        );

    \I__686\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5379\
        );

    \I__685\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5376\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5373\
        );

    \I__683\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5370\
        );

    \I__682\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5367\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5360\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5382\,
            I => \N__5360\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5379\,
            I => \N__5360\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5370\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5367\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__5360\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.N_366_cascade_\
        );

    \I__672\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5343\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5340\
        );

    \I__670\ : Span4Mux_v
    port map (
            O => \N__5340\,
            I => \N__5336\
        );

    \I__669\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5333\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__5328\,
            I => \U712_CHIP_RAM.DBENn_8_1_cascade_\
        );

    \I__665\ : IoInMux
    port map (
            O => \N__5325\,
            I => \N__5322\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__663\ : IoSpan4Mux
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__662\ : Span4Mux_s2_v
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__661\ : Sp12to4
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__660\ : Span12Mux_s11_v
    port map (
            O => \N__5310\,
            I => \N__5306\
        );

    \I__659\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5303\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__5306\,
            I => \DBDIR_c\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5303\,
            I => \DBDIR_c\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__5298\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_\
        );

    \I__655\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5289\
        );

    \I__654\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5289\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5285\
        );

    \I__652\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5282\
        );

    \I__651\ : Span4Mux_h
    port map (
            O => \N__5285\,
            I => \N__5277\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5277\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__648\ : Sp12to4
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__647\ : Span12Mux_h
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__5268\,
            I => \AWEn_c\
        );

    \I__645\ : IoInMux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__643\ : Span4Mux_s2_v
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__642\ : Sp12to4
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__641\ : Span12Mux_h
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__640\ : Span12Mux_v
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__639\ : Odrv12
    port map (
            O => \N__5247\,
            I => \DMA_LATCH_EN_c\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__5244\,
            I => \U712_CHIP_RAM.N_343_cascade_\
        );

    \I__637\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5238\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__635\ : IoInMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__633\ : IoSpan4Mux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__632\ : Span4Mux_s2_v
    port map (
            O => \N__5226\,
            I => \N__5222\
        );

    \I__631\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5219\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__5222\,
            I => \N__5216\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5219\,
            I => \N__5213\
        );

    \I__628\ : Span12Mux_s8_v
    port map (
            O => \N__5216\,
            I => \N__5210\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__5213\,
            I => \N__5207\
        );

    \I__626\ : Span12Mux_v
    port map (
            O => \N__5210\,
            I => \N__5202\
        );

    \I__625\ : Sp12to4
    port map (
            O => \N__5207\,
            I => \N__5202\
        );

    \I__624\ : Span12Mux_h
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__623\ : Odrv12
    port map (
            O => \N__5199\,
            I => \A_c_10\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__5196\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__621\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5190\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__619\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5184\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__617\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5177\
        );

    \I__616\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5174\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5171\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__5174\,
            I => \N__5168\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__5171\,
            I => \U712_CHIP_RAM.N_334\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__5168\,
            I => \U712_CHIP_RAM.N_334\
        );

    \I__611\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5159\
        );

    \I__610\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5156\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5159\,
            I => \N__5153\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5156\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0\
        );

    \I__606\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5145\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5145\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1\
        );

    \I__604\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5138\
        );

    \I__603\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5135\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5138\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5135\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__600\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5126\
        );

    \I__599\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5123\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5123\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__5118\,
            I => \N__5114\
        );

    \I__595\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5111\
        );

    \I__594\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5108\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__5111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5108\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__591\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5099\
        );

    \I__590\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__5099\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5096\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__5091\,
            I => \U712_CHIP_RAM.N_332_cascade_\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \U712_CHIP_RAM.N_510_cascade_\
        );

    \I__585\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5082\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__583\ : IoInMux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__581\ : Span4Mux_s1_v
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__580\ : Sp12to4
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__579\ : Span12Mux_h
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__578\ : Span12Mux_v
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__5061\,
            I => \CMA_c_0\
        );

    \I__576\ : IoInMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__574\ : IoSpan4Mux
    port map (
            O => \N__5052\,
            I => \N__5049\
        );

    \I__573\ : Span4Mux_s2_v
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__572\ : Sp12to4
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__571\ : Odrv12
    port map (
            O => \N__5043\,
            I => \CMA_c_1\
        );

    \I__570\ : IoInMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__568\ : IoSpan4Mux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__567\ : IoSpan4Mux
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__565\ : Span12Mux_s7_h
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__564\ : Span12Mux_h
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__563\ : Odrv12
    port map (
            O => \N__5019\,
            I => \CMA_c_5\
        );

    \I__562\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5013\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__560\ : InMux
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__5007\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__5004\,
            I => \U712_CHIP_RAM.N_583_cascade_\
        );

    \I__557\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4998\,
            I => \U712_CHIP_RAM.N_591\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__4995\,
            I => \U712_CHIP_RAM.N_402_cascade_\
        );

    \I__554\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4983\
        );

    \I__553\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4976\
        );

    \I__552\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4976\
        );

    \I__551\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4976\
        );

    \I__550\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4969\
        );

    \I__549\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4969\
        );

    \I__548\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4969\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4983\,
            I => \U712_CHIP_RAM.N_375_0_i\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4976\,
            I => \U712_CHIP_RAM.N_375_0_i\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4969\,
            I => \U712_CHIP_RAM.N_375_0_i\
        );

    \I__544\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4959\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4956\,
            I => \U712_CHIP_RAM.N_375_0_i_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4950\,
            I => \U712_CHIP_RAM.N_402\
        );

    \I__539\ : CEMux
    port map (
            O => \N__4947\,
            I => \N__4943\
        );

    \I__538\ : CEMux
    port map (
            O => \N__4946\,
            I => \N__4940\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4943\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4940\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__535\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4932\,
            I => \U712_CHIP_RAM.N_426\
        );

    \I__533\ : IoInMux
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__531\ : IoSpan4Mux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__530\ : Span4Mux_s1_h
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__528\ : Span12Mux_h
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__4908\,
            I => \CLK_EN_c\
        );

    \I__525\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4901\
        );

    \I__524\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4898\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4893\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4893\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__4893\,
            I => \U712_CHIP_RAM.N_586\
        );

    \I__520\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__4884\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__4881\,
            I => \U712_CHIP_RAM.N_586_cascade_\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__4878\,
            I => \U712_CHIP_RAM.N_419_cascade_\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_349_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4866\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4866\,
            I => \U712_CHIP_RAM.N_349\
        );

    \I__511\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4860\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__508\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4849\
        );

    \I__507\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4846\
        );

    \I__506\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4843\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4849\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__4836\,
            I => \U712_CHIP_RAM.N_509_cascade_\
        );

    \I__501\ : IoInMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4826\
        );

    \I__499\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4823\
        );

    \I__498\ : Span12Mux_s4_v
    port map (
            O => \N__4826\,
            I => \N__4820\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__496\ : Span12Mux_h
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__495\ : Span4Mux_v
    port map (
            O => \N__4817\,
            I => \N__4811\
        );

    \I__494\ : Span12Mux_v
    port map (
            O => \N__4814\,
            I => \N__4808\
        );

    \I__493\ : Sp12to4
    port map (
            O => \N__4811\,
            I => \N__4805\
        );

    \I__492\ : Odrv12
    port map (
            O => \N__4808\,
            I => \A_c_9\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__4805\,
            I => \A_c_9\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__4800\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__489\ : IoInMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__487\ : Span12Mux_s8_v
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__4788\,
            I => \VBENn_c\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__483\ : Span12Mux_s6_v
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__482\ : Span12Mux_h
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__481\ : Odrv12
    port map (
            O => \N__4773\,
            I => \CMA_c_10\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__478\ : IoSpan4Mux
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__477\ : Span4Mux_s2_v
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__476\ : Sp12to4
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__475\ : Span12Mux_s8_v
    port map (
            O => \N__4755\,
            I => \N__4751\
        );

    \I__474\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__4751\,
            I => \N__4745\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4748\,
            I => \N__4742\
        );

    \I__471\ : Span12Mux_h
    port map (
            O => \N__4745\,
            I => \N__4737\
        );

    \I__470\ : Span12Mux_v
    port map (
            O => \N__4742\,
            I => \N__4737\
        );

    \I__469\ : Odrv12
    port map (
            O => \N__4737\,
            I => \A_c_11\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4734\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__4731\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__466\ : IoInMux
    port map (
            O => \N__4728\,
            I => \N__4725\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4725\,
            I => \N__4722\
        );

    \I__464\ : Span4Mux_s3_v
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__463\ : Sp12to4
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__462\ : Span12Mux_h
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__461\ : Span12Mux_v
    port map (
            O => \N__4713\,
            I => \N__4710\
        );

    \I__460\ : Odrv12
    port map (
            O => \N__4710\,
            I => \CMA_c_2\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__4707\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER19_cascade_\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__4704\,
            I => \U712_CHIP_RAM.N_335_cascade_\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4701\,
            I => \U712_CHIP_RAM.N_507_cascade_\
        );

    \I__456\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4695\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__4692\,
            I => \U712_CHIP_RAM.N_477\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__4689\,
            I => \U712_CHIP_RAM.N_477_cascade_\
        );

    \I__452\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4679\
        );

    \I__451\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4679\
        );

    \I__450\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4676\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4679\,
            I => \N__4673\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4676\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__4673\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__4668\,
            I => \U712_CYCLE_TERM.N_406_cascade_\
        );

    \I__445\ : IoInMux
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__443\ : Span4Mux_s3_h
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__441\ : Span12Mux_v
    port map (
            O => \N__4653\,
            I => \N__4649\
        );

    \I__440\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__4649\,
            I => \TACK_OUT\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4646\,
            I => \TACK_OUT\
        );

    \I__437\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0\
        );

    \I__435\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4632\,
            I => \U712_CHIP_RAM.N_478\
        );

    \I__433\ : InMux
    port map (
            O => \N__4629\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__432\ : InMux
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__431\ : InMux
    port map (
            O => \N__4623\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__430\ : InMux
    port map (
            O => \N__4620\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__429\ : InMux
    port map (
            O => \N__4617\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__428\ : InMux
    port map (
            O => \N__4614\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__427\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__4605\,
            I => \U712_CHIP_RAM.N_483\
        );

    \I__424\ : IoInMux
    port map (
            O => \N__4602\,
            I => \N__4598\
        );

    \I__423\ : IoInMux
    port map (
            O => \N__4601\,
            I => \N__4595\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4598\,
            I => \N__4592\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__420\ : IoSpan4Mux
    port map (
            O => \N__4592\,
            I => \N__4584\
        );

    \I__419\ : IoSpan4Mux
    port map (
            O => \N__4589\,
            I => \N__4584\
        );

    \I__418\ : Span4Mux_s3_v
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__417\ : Sp12to4
    port map (
            O => \N__4581\,
            I => \N__4577\
        );

    \I__416\ : IoInMux
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__4577\,
            I => \N__4571\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__413\ : Span12Mux_h
    port map (
            O => \N__4571\,
            I => \N__4563\
        );

    \I__412\ : Span12Mux_s5_h
    port map (
            O => \N__4568\,
            I => \N__4563\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__4563\,
            I => \CLK40_PLL_i_i\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__4560\,
            I => \U712_CHIP_RAM.N_592_cascade_\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__4557\,
            I => \U712_CHIP_RAM.N_482_cascade_\
        );

    \I__408\ : InMux
    port map (
            O => \N__4554\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__405\ : Span4Mux_s3_h
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__4542\,
            I => \DBRn_c_i_0\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__4533\,
            I => \N__4530\
        );

    \I__400\ : Span4Mux_s2_v
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4524\,
            I => \CLK80_PLL_iso_i\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__395\ : Span4Mux_s0_v
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__393\ : Sp12to4
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__392\ : Span12Mux_h
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__391\ : Span12Mux_v
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__4500\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__9627\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__9624\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__9625\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__9626\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__9629\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__9628\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__9630\
        );

    \INVU712_CYCLE_TERM.TACK_STATE_1C\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_STATE_1C_net\,
            I => \N__10220\
        );

    \INVU712_CYCLE_TERM.TACK_OUTC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            I => \N__10228\
        );

    \INVU712_CYCLE_TERM.TACK_STATE_3C\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_STATE_3C_net\,
            I => \N__10231\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5967\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9348\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4551\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7494\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7544\,
            in2 => \_gnd_net_\,
            in3 => \N__10725\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10236\,
            lcout => \CLK80_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5628\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5646\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_3C_net\,
            ce => 'H',
            sr => \N__10673\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4684\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_3C_net\,
            ce => 'H',
            sr => \N__10673\
        );

    \pll_RNI8MQ3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5506\,
            in1 => \N__7130\,
            in2 => \_gnd_net_\,
            in3 => \N__6548\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5858\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__4698\,
            in2 => \N__4560\,
            in3 => \N__8699\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110000"
        )
    port map (
            in0 => \N__6472\,
            in1 => \N__6549\,
            in2 => \N__7158\,
            in3 => \N__8338\,
            lcout => \U712_CHIP_RAM.N_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__5859\,
            in1 => \N__10445\,
            in2 => \N__5400\,
            in3 => \N__8339\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__4611\,
            in1 => \N__6773\,
            in2 => \N__4557\,
            in3 => \N__9996\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8335\,
            in2 => \_gnd_net_\,
            in3 => \N__11097\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4989\,
            in1 => \N__7138\,
            in2 => \_gnd_net_\,
            in3 => \N__4554\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6574\,
            in2 => \_gnd_net_\,
            in3 => \N__4629\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4990\,
            in1 => \N__6473\,
            in2 => \_gnd_net_\,
            in3 => \N__4626\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4986\,
            in1 => \N__5117\,
            in2 => \_gnd_net_\,
            in3 => \N__4623\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4991\,
            in1 => \N__5130\,
            in2 => \_gnd_net_\,
            in3 => \N__4620\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4987\,
            in1 => \N__5142\,
            in2 => \_gnd_net_\,
            in3 => \N__4617\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__5103\,
            in1 => \N__4988\,
            in2 => \_gnd_net_\,
            in3 => \N__4614\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10218\,
            ce => \N__4947\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__8364\,
            in2 => \_gnd_net_\,
            in3 => \N__6552\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4852\,
            in1 => \N__8359\,
            in2 => \N__7049\,
            in3 => \N__5533\,
            lcout => \U712_CHIP_RAM.N_483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2EV43_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5532\,
            in1 => \N__6551\,
            in2 => \N__7157\,
            in3 => \N__7030\,
            lcout => \U712_CHIP_RAM.N_590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8357\,
            in2 => \_gnd_net_\,
            in3 => \N__7134\,
            lcout => \U712_CHIP_RAM.N_335\,
            ltout => \U712_CHIP_RAM.N_335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10501\,
            in1 => \N__6471\,
            in2 => \N__4704\,
            in3 => \N__6553\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5EAU6_3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__5163\,
            in1 => \N__7042\,
            in2 => \N__4701\,
            in3 => \N__5181\,
            lcout => \U712_CHIP_RAM.N_477\,
            ltout => \U712_CHIP_RAM.N_477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__4635\,
            in1 => \N__6766\,
            in2 => \N__4689\,
            in3 => \N__7592\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIN90C1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11088\,
            in1 => \N__10499\,
            in2 => \N__5547\,
            in3 => \N__8358\,
            lcout => \U712_CHIP_RAM.N_504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4685\,
            in2 => \_gnd_net_\,
            in3 => \N__5645\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__5712\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__10496\,
            in1 => \N__4686\,
            in2 => \N__4668\,
            in3 => \N__4652\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7159\,
            in1 => \N__4641\,
            in2 => \N__7058\,
            in3 => \N__5546\,
            lcout => \U712_CHIP_RAM.N_478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4829\,
            in1 => \N__6240\,
            in2 => \_gnd_net_\,
            in3 => \N__8002\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8003\,
            in1 => \N__11893\,
            in2 => \N__4800\,
            in3 => \N__8652\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11902\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__8000\,
            in1 => \N__6051\,
            in2 => \N__8712\,
            in3 => \_gnd_net_\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10204\,
            ce => \N__6315\,
            sr => \N__10686\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7998\,
            in1 => \N__4754\,
            in2 => \_gnd_net_\,
            in3 => \N__6681\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__11901\,
            in1 => \N__7999\,
            in2 => \N__4734\,
            in3 => \N__8859\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__6356\,
            in1 => \N__6052\,
            in2 => \N__4731\,
            in3 => \N__9705\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10204\,
            ce => \N__6315\,
            sr => \N__10686\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8342\,
            in1 => \N__4904\,
            in2 => \N__7163\,
            in3 => \N__6561\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10451\,
            in2 => \N__4707\,
            in3 => \N__5525\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10210\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIGDNC1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100010111"
        )
    port map (
            in0 => \N__8340\,
            in1 => \N__6559\,
            in2 => \N__5540\,
            in3 => \N__5389\,
            lcout => \U712_CHIP_RAM.N_349\,
            ltout => \U712_CHIP_RAM.N_349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI6NJS1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10455\,
            in2 => \N__4872\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8341\,
            in1 => \N__6560\,
            in2 => \N__5541\,
            in3 => \N__6816\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10452\,
            in2 => \_gnd_net_\,
            in3 => \N__5518\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__10454\,
            in1 => \N__4853\,
            in2 => \_gnd_net_\,
            in3 => \N__4869\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10453\,
            in2 => \_gnd_net_\,
            in3 => \N__6464\,
            lcout => \U712_CHIP_RAM.N_501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__4863\,
            in1 => \N__6870\,
            in2 => \N__4857\,
            in3 => \N__4992\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10214\,
            ce => \N__4946\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILQND1_3_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6466\,
            in1 => \N__10497\,
            in2 => \_gnd_net_\,
            in3 => \N__6557\,
            lcout => \U712_CHIP_RAM.N_509\,
            ltout => \U712_CHIP_RAM.N_509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__7274\,
            in1 => \N__7200\,
            in2 => \N__4836\,
            in3 => \N__7356\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7F93_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__6465\,
            in1 => \N__10498\,
            in2 => \N__7066\,
            in3 => \N__7173\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_583_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI615I6_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5010\,
            in1 => \N__6812\,
            in2 => \N__5004\,
            in3 => \N__5339\,
            lcout => \U712_CHIP_RAM.N_402\,
            ltout => \U712_CHIP_RAM.N_402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISSQMA_3_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__6467\,
            in1 => \N__5001\,
            in2 => \N__4995\,
            in3 => \N__4935\,
            lcout => \U712_CHIP_RAM.N_375_0_i\,
            ltout => \U712_CHIP_RAM.N_375_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__8259\,
            in2 => \N__4956\,
            in3 => \N__4953\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10214\,
            ce => \N__4946\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGB4P1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6811\,
            in1 => \N__6558\,
            in2 => \_gnd_net_\,
            in3 => \N__5527\,
            lcout => \U712_CHIP_RAM.N_426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6556\,
            in1 => \N__7124\,
            in2 => \N__8378\,
            in3 => \N__4905\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10219\,
            ce => \N__5556\,
            sr => \N__10665\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6454\,
            in2 => \_gnd_net_\,
            in3 => \N__7035\,
            lcout => \U712_CHIP_RAM.N_586\,
            ltout => \U712_CHIP_RAM.N_586_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8360\,
            in1 => \N__4890\,
            in2 => \N__4881\,
            in3 => \N__10471\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIADE59_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6824\,
            in1 => \N__6555\,
            in2 => \N__4878\,
            in3 => \N__7354\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOV5BI_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__7729\,
            in2 => \N__4875\,
            in3 => \N__10472\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__5129\,
            in2 => \N__5118\,
            in3 => \N__5102\,
            lcout => \U712_CHIP_RAM.N_332\,
            ltout => \U712_CHIP_RAM.N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6455\,
            in1 => \N__7123\,
            in2 => \N__5091\,
            in3 => \N__5531\,
            lcout => \U712_CHIP_RAM.N_510\,
            ltout => \U712_CHIP_RAM.N_510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8365\,
            in1 => \N__6554\,
            in2 => \N__5088\,
            in3 => \N__5395\,
            lcout => \U712_CHIP_RAM.N_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7275\,
            in1 => \N__7308\,
            in2 => \_gnd_net_\,
            in3 => \N__7358\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10224\,
            ce => \N__5448\,
            sr => \N__10654\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11621\,
            in1 => \N__11558\,
            in2 => \N__6942\,
            in3 => \N__11430\,
            lcout => \U712_REG_SM.N_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__6357\,
            in1 => \N__8640\,
            in2 => \N__6060\,
            in3 => \N__5085\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10193\,
            ce => \N__6314\,
            sr => \N__10691\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5241\,
            in1 => \N__5187\,
            in2 => \_gnd_net_\,
            in3 => \N__5193\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10196\,
            ce => \N__6307\,
            sr => \N__10687\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__6162\,
            in1 => \N__6053\,
            in2 => \N__8007\,
            in3 => \N__5016\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10196\,
            ce => \N__6307\,
            sr => \N__10687\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11869\,
            in1 => \N__6651\,
            in2 => \_gnd_net_\,
            in3 => \N__7506\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7611\,
            in2 => \_gnd_net_\,
            in3 => \N__10009\,
            lcout => \U712_CHIP_RAM.N_343\,
            ltout => \U712_CHIP_RAM.N_343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__9339\,
            in1 => \N__11868\,
            in2 => \N__5244\,
            in3 => \N__7963\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5225\,
            in1 => \N__6705\,
            in2 => \_gnd_net_\,
            in3 => \N__7958\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7964\,
            in1 => \N__11871\,
            in2 => \N__5196\,
            in3 => \N__8868\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__10010\,
            in1 => \N__7612\,
            in2 => \_gnd_net_\,
            in3 => \N__7959\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110000101"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__9338\,
            in2 => \N__7989\,
            in3 => \N__11870\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__5180\,
            in1 => \N__5162\,
            in2 => \N__7068\,
            in3 => \N__5148\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8336\,
            in1 => \N__5388\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__7273\,
            in1 => \N__6966\,
            in2 => \_gnd_net_\,
            in3 => \N__5295\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__6869\,
            in2 => \N__5349\,
            in3 => \N__7304\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10205\,
            ce => 'H',
            sr => \N__10674\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5346\,
            in1 => \N__7303\,
            in2 => \_gnd_net_\,
            in3 => \N__7065\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DBENn_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__11158\,
            in1 => \N__5415\,
            in2 => \N__5328\,
            in3 => \N__9132\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10205\,
            ce => 'H',
            sr => \N__10674\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5294\,
            in1 => \N__5309\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10205\,
            ce => 'H',
            sr => \N__10674\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5394\,
            in2 => \_gnd_net_\,
            in3 => \N__6547\,
            lcout => \U712_CHIP_RAM.N_350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQS0H1_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__6476\,
            in2 => \N__7172\,
            in3 => \N__11813\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN2IA4_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6854\,
            in1 => \N__5526\,
            in2 => \N__5298\,
            in3 => \N__7034\,
            lcout => \U712_CHIP_RAM.N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__5288\,
            in1 => \N__5593\,
            in2 => \N__10502\,
            in3 => \N__5441\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__5594\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__11268\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001111111"
        )
    port map (
            in0 => \N__11358\,
            in1 => \N__6965\,
            in2 => \N__11276\,
            in3 => \N__5595\,
            lcout => \DRDDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__6573\,
            in1 => \N__5837\,
            in2 => \N__8382\,
            in3 => \N__7723\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5559\,
            in3 => \N__10723\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7164\,
            in1 => \N__8333\,
            in2 => \N__5542\,
            in3 => \N__7029\,
            lcout => \U712_CHIP_RAM.N_503\,
            ltout => \U712_CHIP_RAM.N_503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNILPRG5_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__7254\,
            in2 => \N__5457\,
            in3 => \N__6823\,
            lcout => \U712_CHIP_RAM.N_420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5411\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7299\,
            in1 => \N__7255\,
            in2 => \_gnd_net_\,
            in3 => \N__7353\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIAGI99_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__5427\,
            in1 => \N__7758\,
            in2 => \N__5418\,
            in3 => \N__7722\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__8334\,
            in1 => \N__5396\,
            in2 => \_gnd_net_\,
            in3 => \N__6480\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__5857\,
            in1 => \N__5838\,
            in2 => \N__5826\,
            in3 => \N__7694\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5823\,
            in3 => \N__10721\,
            lcout => \U712_CHIP_RAM.N_248_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__5666\,
            in1 => \N__5714\,
            in2 => \N__5802\,
            in3 => \N__5820\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_1C_net\,
            ce => 'H',
            sr => \N__10651\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__5665\,
            in1 => \N__5790\,
            in2 => \N__5814\,
            in3 => \N__5811\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_1C_net\,
            ce => 'H',
            sr => \N__10651\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__6902\,
            in1 => \N__5798\,
            in2 => \_gnd_net_\,
            in3 => \N__6984\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_358_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5789\,
            in2 => \N__5778\,
            in3 => \N__5733\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_1C_net\,
            ce => 'H',
            sr => \N__10651\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__5715\,
            in1 => \N__5664\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_1C_net\,
            ce => 'H',
            sr => \N__10651\
        );

    \DBR_SYNC_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5627\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10225\,
            ce => 'H',
            sr => \N__10649\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10225\,
            ce => 'H',
            sr => \N__10649\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8513\,
            in2 => \_gnd_net_\,
            in3 => \N__9409\,
            lcout => \U712_REG_SM.N_352\,
            ltout => \U712_REG_SM.N_352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10503\,
            in1 => \N__8198\,
            in2 => \N__5970\,
            in3 => \N__7401\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8514\,
            in2 => \_gnd_net_\,
            in3 => \N__9410\,
            lcout => \U712_REG_SM.N_353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => 'H',
            sr => \N__10647\
        );

    \U712_REG_SM.UDSn_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__5912\,
            in1 => \N__8762\,
            in2 => \N__9446\,
            in3 => \N__5865\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => 'H',
            sr => \N__10647\
        );

    \U712_REG_SM.LDSn_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__5901\,
            in1 => \N__9436\,
            in2 => \N__5882\,
            in3 => \N__8763\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10232\,
            ce => 'H',
            sr => \N__10647\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__6952\,
            in1 => \N__11638\,
            in2 => \N__11575\,
            in3 => \N__11453\,
            lcout => \U712_REG_SM.N_493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7967\,
            in1 => \N__11873\,
            in2 => \N__6213\,
            in3 => \N__7512\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7965\,
            in1 => \N__6591\,
            in2 => \_gnd_net_\,
            in3 => \N__6228\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__7966\,
            in2 => \_gnd_net_\,
            in3 => \N__7776\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__11874\,
            in1 => \N__7968\,
            in2 => \N__6180\,
            in3 => \N__7523\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6177\,
            in1 => \N__11872\,
            in2 => \_gnd_net_\,
            in3 => \N__8607\,
            lcout => \U712_CHIP_RAM.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__6345\,
            in1 => \N__8619\,
            in2 => \N__6057\,
            in3 => \N__6264\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__6049\,
            in1 => \N__6346\,
            in2 => \N__9903\,
            in3 => \N__8073\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__6347\,
            in1 => \N__9324\,
            in2 => \N__6058\,
            in3 => \N__8031\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__6050\,
            in1 => \N__6348\,
            in2 => \N__6093\,
            in3 => \N__8877\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__6349\,
            in1 => \N__8628\,
            in2 => \N__6059\,
            in3 => \N__5997\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__6405\,
            in1 => \N__6399\,
            in2 => \N__11903\,
            in3 => \N__10800\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10194\,
            ce => \N__6306\,
            sr => \N__10682\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11863\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10008\,
            in1 => \N__7953\,
            in2 => \N__7616\,
            in3 => \N__8713\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__7954\,
            in1 => \N__7610\,
            in2 => \N__6321\,
            in3 => \N__8714\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6318\,
            in3 => \N__10724\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__10425\,
            in1 => \N__8946\,
            in2 => \N__8067\,
            in3 => \N__9005\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6282\,
            in1 => \N__6615\,
            in2 => \_gnd_net_\,
            in3 => \N__7956\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7957\,
            in1 => \N__11864\,
            in2 => \N__6267\,
            in3 => \N__9123\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6258\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6669\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6645\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6609\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10200\,
            ce => \N__7829\,
            sr => \N__10666\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6475\,
            in1 => \N__8369\,
            in2 => \N__6579\,
            in3 => \N__11839\,
            lcout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6575\,
            in2 => \_gnd_net_\,
            in3 => \N__6474\,
            lcout => \U712_CHIP_RAM.N_514\,
            ltout => \U712_CHIP_RAM.N_514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7260\,
            in1 => \N__7357\,
            in2 => \N__6873\,
            in3 => \N__7368\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10206\,
            ce => \N__6840\,
            sr => \N__10655\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIVM1I4_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7367\,
            in1 => \N__7259\,
            in2 => \_gnd_net_\,
            in3 => \N__7355\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10720\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6855\,
            in1 => \N__7736\,
            in2 => \N__8379\,
            in3 => \N__7789\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6843\,
            in3 => \N__10719\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8151\,
            in1 => \N__7252\,
            in2 => \N__7359\,
            in3 => \N__6828\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_481_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__6772\,
            in2 => \N__6747\,
            in3 => \N__7981\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6888\,
            in2 => \_gnd_net_\,
            in3 => \N__8219\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__10477\,
            in1 => \N__8138\,
            in2 => \N__6744\,
            in3 => \N__6741\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8149\,
            in1 => \N__7214\,
            in2 => \_gnd_net_\,
            in3 => \N__8086\,
            lcout => \U712_CHIP_RAM.N_500\,
            ltout => \U712_CHIP_RAM.N_500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7251\,
            in1 => \N__7349\,
            in2 => \N__7311\,
            in3 => \N__7298\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__10476\,
            in2 => \N__11142\,
            in3 => \N__7253\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__8087\,
            in1 => \N__8150\,
            in2 => \_gnd_net_\,
            in3 => \N__7215\,
            lcout => \U712_CHIP_RAM.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__7182\,
            in1 => \N__7171\,
            in2 => \_gnd_net_\,
            in3 => \N__7067\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10215\,
            ce => \N__6975\,
            sr => \N__10650\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__8591\,
            in1 => \N__7399\,
            in2 => \_gnd_net_\,
            in3 => \N__6958\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \DBR_SYNC_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6912\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.REG_TACK_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__8556\,
            in2 => \N__6906\,
            in3 => \N__8568\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.START_RST_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__7400\,
            in1 => \N__6887\,
            in2 => \_gnd_net_\,
            in3 => \N__8197\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.C3_SYNC_0_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7475\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.REGENn_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__7423\,
            in2 => \_gnd_net_\,
            in3 => \N__9506\,
            lcout => \BLSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.C3_SYNC_1_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7410\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10221\,
            ce => 'H',
            sr => \N__10648\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8516\,
            in2 => \_gnd_net_\,
            in3 => \N__9412\,
            lcout => \U712_REG_SM.N_345\,
            ltout => \U712_REG_SM.N_345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9477\,
            in2 => \N__7404\,
            in3 => \N__8223\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__7656\,
            in1 => \N__7386\,
            in2 => \N__9443\,
            in3 => \N__10506\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__8193\,
            in1 => \N__8544\,
            in2 => \_gnd_net_\,
            in3 => \N__7377\,
            lcout => \U712_REG_SM.N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8474\,
            in1 => \N__8515\,
            in2 => \_gnd_net_\,
            in3 => \N__9411\,
            lcout => \U712_REG_SM.N_435\,
            ltout => \U712_REG_SM.N_435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__8192\,
            in1 => \_gnd_net_\,
            in2 => \N__7380\,
            in3 => \N__7376\,
            lcout => \U712_REG_SM.N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8983\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \U712_REG_SM.N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8590\,
            in1 => \N__8475\,
            in2 => \N__7650\,
            in3 => \N__8821\,
            lcout => \U712_REG_SM.REG_CYCLE_5_iv_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__8745\,
            in1 => \N__7649\,
            in2 => \N__8484\,
            in3 => \N__10509\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10187\,
            ce => 'H',
            sr => \N__10692\
        );

    \U712_CHIP_RAM.RASn_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7617\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10191\,
            ce => 'H',
            sr => \N__10688\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__11042\,
            in1 => \N__10862\,
            in2 => \N__7551\,
            in3 => \N__7524\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__10683\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11038\,
            in1 => \N__10863\,
            in2 => \_gnd_net_\,
            in3 => \N__9315\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10757\,
            sr => \N__10675\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9273\,
            in1 => \N__11037\,
            in2 => \_gnd_net_\,
            in3 => \N__9888\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10757\,
            sr => \N__10675\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__7863\,
            in1 => \N__11876\,
            in2 => \N__9801\,
            in3 => \N__7984\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8895\,
            in1 => \N__8850\,
            in2 => \_gnd_net_\,
            in3 => \N__9004\,
            lcout => \U712_CHIP_RAM.N_450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8058\,
            in1 => \N__8040\,
            in2 => \_gnd_net_\,
            in3 => \N__7983\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__11875\,
            in1 => \N__7985\,
            in2 => \N__8034\,
            in3 => \N__9231\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8025\,
            in1 => \N__7839\,
            in2 => \_gnd_net_\,
            in3 => \N__7982\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7857\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10198\,
            ce => \N__7833\,
            sr => \N__10656\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__7772\,
            in2 => \N__11043\,
            in3 => \N__7791\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10201\,
            ce => 'H',
            sr => \N__10652\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7757\,
            in1 => \N__7737\,
            in2 => \_gnd_net_\,
            in3 => \N__7701\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__7667\,
            in1 => \N__11111\,
            in2 => \N__7683\,
            in3 => \N__8381\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10201\,
            ce => 'H',
            sr => \N__10652\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8380\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.PRnW_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110100110001"
        )
    port map (
            in0 => \N__8595\,
            in1 => \N__8165\,
            in2 => \N__8532\,
            in3 => \N__8234\,
            lcout => \PRnW_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10201\,
            ce => 'H',
            sr => \N__10652\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9468\,
            in2 => \_gnd_net_\,
            in3 => \N__8218\,
            lcout => \U712_REG_SM.N_351\,
            ltout => \U712_REG_SM.N_351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110001"
        )
    port map (
            in0 => \N__8525\,
            in1 => \N__8202\,
            in2 => \N__8169\,
            in3 => \N__9444\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__9648\,
            in1 => \N__10026\,
            in2 => \N__10450\,
            in3 => \N__10059\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11859\,
            in2 => \_gnd_net_\,
            in3 => \N__8088\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__8139\,
            in1 => \N__8118\,
            in2 => \N__8091\,
            in3 => \N__10394\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8974\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8589\,
            in1 => \N__8428\,
            in2 => \_gnd_net_\,
            in3 => \N__8483\,
            lcout => \U712_REG_SM.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10479\,
            in2 => \_gnd_net_\,
            in3 => \N__8562\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8429\,
            in1 => \N__10478\,
            in2 => \_gnd_net_\,
            in3 => \N__9501\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8427\,
            in2 => \_gnd_net_\,
            in3 => \N__9500\,
            lcout => \U712_REG_SM.N_588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_2_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__8735\,
            in1 => \N__9521\,
            in2 => \_gnd_net_\,
            in3 => \N__9472\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__8543\,
            in1 => \N__8524\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \U712_REG_SM.N_395\,
            ltout => \U712_REG_SM.N_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8479\,
            in2 => \N__8451\,
            in3 => \N__9447\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_439_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__10504\,
            in1 => \N__8822\,
            in2 => \N__8448\,
            in3 => \N__8445\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__10505\,
            in1 => \N__9502\,
            in2 => \N__8433\,
            in3 => \N__8439\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10718\,
            in2 => \_gnd_net_\,
            in3 => \N__8761\,
            lcout => \U712_REG_SM.N_131_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8724\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8739\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8718\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10186\,
            ce => 'H',
            sr => \N__10681\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11036\,
            in1 => \N__9750\,
            in2 => \_gnd_net_\,
            in3 => \N__9192\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10762\,
            sr => \N__10672\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9222\,
            in1 => \N__11006\,
            in2 => \_gnd_net_\,
            in3 => \N__9187\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10760\,
            sr => \N__10664\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9301\,
            in1 => \N__11014\,
            in2 => \_gnd_net_\,
            in3 => \N__10861\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10760\,
            sr => \N__10664\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9789\,
            in1 => \_gnd_net_\,
            in2 => \N__11034\,
            in3 => \N__9957\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10760\,
            sr => \N__10664\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11010\,
            in1 => \N__9887\,
            in2 => \_gnd_net_\,
            in3 => \N__9843\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10760\,
            sr => \N__10664\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9272\,
            in1 => \_gnd_net_\,
            in2 => \N__11035\,
            in3 => \N__9300\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10790\,
            ce => \N__10760\,
            sr => \N__10664\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9742\,
            in1 => \N__11001\,
            in2 => \_gnd_net_\,
            in3 => \N__9787\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10758\,
            sr => \N__10653\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9788\,
            in1 => \_gnd_net_\,
            in2 => \N__11033\,
            in3 => \N__9956\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10758\,
            sr => \N__10653\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__9068\,
            in2 => \N__8941\,
            in3 => \N__9102\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_196_i_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__11277\,
            in1 => \N__11351\,
            in2 => \N__8840\,
            in3 => \N__11886\,
            lcout => \N_196_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9111\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__8933\,
            in1 => \N__10348\,
            in2 => \N__9033\,
            in3 => \N__9011\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8781\,
            in1 => \N__9110\,
            in2 => \_gnd_net_\,
            in3 => \N__8931\,
            lcout => \U712_CHIP_RAM.N_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__8932\,
            in1 => \N__10347\,
            in2 => \N__9057\,
            in3 => \N__9010\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10346\,
            in1 => \N__9075\,
            in2 => \N__9012\,
            in3 => \N__8934\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10350\,
            in2 => \_gnd_net_\,
            in3 => \N__9693\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9018\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9101\,
            in2 => \N__9090\,
            in3 => \N__9089\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9069\,
            in2 => \_gnd_net_\,
            in3 => \N__9048\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9045\,
            in2 => \_gnd_net_\,
            in3 => \N__9024\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8888\,
            in2 => \_gnd_net_\,
            in3 => \N__9021\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11350\,
            in1 => \N__10353\,
            in2 => \_gnd_net_\,
            in3 => \N__11267\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__10352\,
            in1 => \N__9006\,
            in2 => \N__8945\,
            in3 => \N__8901\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__9537\,
            in1 => \N__9473\,
            in2 => \N__9531\,
            in3 => \N__9510\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10203\,
            ce => 'H',
            sr => \N__10646\
        );

    \U712_REG_SM.ASn_ess_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9445\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10217\,
            ce => \N__9357\,
            sr => \N__10642\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10365\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9188\,
            in1 => \N__11015\,
            in2 => \_gnd_net_\,
            in3 => \N__9749\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => \N__10765\,
            sr => \N__10684\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9880\,
            in1 => \N__11005\,
            in2 => \_gnd_net_\,
            in3 => \N__9271\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => \N__10763\,
            sr => \N__10676\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9314\,
            in1 => \N__10994\,
            in2 => \_gnd_net_\,
            in3 => \N__9253\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10761\,
            sr => \N__10667\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__10980\,
            in2 => \_gnd_net_\,
            in3 => \N__9168\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10756\,
            sr => \N__10657\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10981\,
            in1 => \N__9839\,
            in2 => \_gnd_net_\,
            in3 => \N__9948\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10756\,
            sr => \N__10657\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9678\,
            in2 => \_gnd_net_\,
            in3 => \N__9672\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9549\,
            in2 => \_gnd_net_\,
            in3 => \N__9669\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9576\,
            in2 => \_gnd_net_\,
            in3 => \N__9666\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9588\,
            in2 => \_gnd_net_\,
            in3 => \N__9663\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9563\,
            in2 => \_gnd_net_\,
            in3 => \N__9660\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10038\,
            in2 => \_gnd_net_\,
            in3 => \N__9657\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10050\,
            in2 => \_gnd_net_\,
            in3 => \N__9654\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9644\,
            in2 => \_gnd_net_\,
            in3 => \N__9651\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9623\,
            ce => 'H',
            sr => \N__9600\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__9587\,
            in1 => \N__9575\,
            in2 => \N__9564\,
            in3 => \N__9548\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10049\,
            in2 => \_gnd_net_\,
            in3 => \N__10037\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10017\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10192\,
            ce => 'H',
            sr => \N__10689\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9955\,
            in1 => \N__11020\,
            in2 => \_gnd_net_\,
            in3 => \N__9838\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => \N__10766\,
            sr => \N__10685\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9871\,
            in1 => \N__10982\,
            in2 => \_gnd_net_\,
            in3 => \N__9837\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10764\,
            sr => \N__10677\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__9773\,
            in2 => \_gnd_net_\,
            in3 => \N__9728\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10788\,
            ce => \N__10759\,
            sr => \N__10668\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10375\,
            in2 => \_gnd_net_\,
            in3 => \N__9684\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10242\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11480\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11536\,
            lcout => \U712_BYTE_ENABLE.N_331_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_412_i_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__11711\,
            in1 => \N__11669\,
            in2 => \N__11551\,
            in3 => \N__11470\,
            lcout => \N_412_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__11019\,
            in2 => \_gnd_net_\,
            in3 => \N__10854\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10786\,
            ce => \N__10767\,
            sr => \N__10690\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10551\,
            in1 => \N__10373\,
            in2 => \_gnd_net_\,
            in3 => \N__10527\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10285\,
            in2 => \_gnd_net_\,
            in3 => \N__10248\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__11727\,
            in1 => \N__11670\,
            in2 => \N__11904\,
            in3 => \N__11921\,
            lcout => \U712_BYTE_ENABLE.N_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11126\,
            in1 => \N__11272\,
            in2 => \_gnd_net_\,
            in3 => \N__11189\,
            lcout => \U712_BYTE_ENABLE.N_467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100000000"
        )
    port map (
            in0 => \N__11481\,
            in1 => \_gnd_net_\,
            in2 => \N__11589\,
            in3 => \N__11907\,
            lcout => \U712_BYTE_ENABLE.N_455\,
            ltout => \U712_BYTE_ENABLE.N_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_38_i_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__11725\,
            in1 => \N__10092\,
            in2 => \N__10086\,
            in3 => \N__11958\,
            lcout => \N_38_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__11906\,
            in1 => \N__11665\,
            in2 => \_gnd_net_\,
            in3 => \N__11583\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_209_i_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__11952\,
            in1 => \N__11724\,
            in2 => \N__11946\,
            in3 => \N__11064\,
            lcout => \N_209_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__11664\,
            in1 => \N__11726\,
            in2 => \N__11922\,
            in3 => \N__11905\,
            lcout => \U712_BYTE_ENABLE.N_464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_i_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111000000"
        )
    port map (
            in0 => \N__11661\,
            in1 => \N__11689\,
            in2 => \N__11582\,
            in3 => \N__11473\,
            lcout => \N_205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_411_i_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__11713\,
            in1 => \N__11663\,
            in2 => \N__11588\,
            in3 => \N__11472\,
            lcout => \N_411_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101010000"
        )
    port map (
            in0 => \N__11712\,
            in1 => \N__11662\,
            in2 => \N__11587\,
            in3 => \N__11471\,
            lcout => \N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_40_i_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__11141\,
            in1 => \N__11388\,
            in2 => \N__11198\,
            in3 => \N__11339\,
            lcout => \N_40_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_208_i_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__11140\,
            in1 => \N__11364\,
            in2 => \N__11349\,
            in3 => \N__11190\,
            lcout => \N_208_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11260\,
            in1 => \N__11194\,
            in2 => \_gnd_net_\,
            in3 => \N__11139\,
            lcout => \U712_BYTE_ENABLE.N_456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 9 2025 17:04:52

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    CIACS1n : out std_logic;
    TICK50 : out std_logic;
    RAMSPACEn : out std_logic;
    TICK60 : out std_logic;
    CLKCIA : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    BUFENn : out std_logic;
    TSn : in std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2499\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_CIA.g0Z0Z_2_cascade_\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_CIA.g0Z0Z_10\ : std_logic;
signal \U409_CIA.g0Z0Z_8_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U409_CIA.g0Z0Z_11\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_20\ : std_logic;
signal \A_c_21\ : std_logic;
signal \CIA_SPACEm_3\ : std_logic;
signal \A_c_22\ : std_logic;
signal \CIA_SPACEm_6\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \A_c_31\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \A_c_23\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un5_RAMSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE_HIROM\ : std_logic;
signal \OVL_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \U409_TICK.TICK503_8\ : std_logic;
signal \U409_TICK.TICK503_11_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_132_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_132\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_359_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5376\,
            RESETB => \N__4596\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6392\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6394\,
            DIN => \N__6393\,
            DOUT => \N__6392\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6394\,
            PADOUT => \N__6393\,
            PADIN => \N__6392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6382\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6384\,
            DIN => \N__6383\,
            DOUT => \N__6382\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6384\,
            PADOUT => \N__6383\,
            PADIN => \N__6382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6373\,
            DIN => \N__6372\,
            DOUT => \N__6371\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6373\,
            PADOUT => \N__6372\,
            PADIN => \N__6371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6364\,
            DIN => \N__6363\,
            DOUT => \N__6362\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6364\,
            PADOUT => \N__6363\,
            PADIN => \N__6362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5169\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6355\,
            DIN => \N__6354\,
            DOUT => \N__6353\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6355\,
            PADOUT => \N__6354\,
            PADIN => \N__6353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6346\,
            DIN => \N__6345\,
            DOUT => \N__6344\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6346\,
            PADOUT => \N__6345\,
            PADIN => \N__6344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6337\,
            DIN => \N__6336\,
            DOUT => \N__6335\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6337\,
            PADOUT => \N__6336\,
            PADIN => \N__6335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3720\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6328\,
            DIN => \N__6327\,
            DOUT => \N__6326\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6328\,
            PADOUT => \N__6327\,
            PADIN => \N__6326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3090\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6319\,
            DIN => \N__6318\,
            DOUT => \N__6317\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6319\,
            PADOUT => \N__6318\,
            PADIN => \N__6317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6310\,
            DIN => \N__6309\,
            DOUT => \N__6308\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6310\,
            PADOUT => \N__6309\,
            PADIN => \N__6308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6301\,
            DIN => \N__6300\,
            DOUT => \N__6299\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6301\,
            PADOUT => \N__6300\,
            PADIN => \N__6299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2961\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6292\,
            DIN => \N__6291\,
            DOUT => \N__6290\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6292\,
            PADOUT => \N__6291\,
            PADIN => \N__6290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5811\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__6045\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6283\,
            DIN => \N__6282\,
            DOUT => \N__6281\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6283\,
            PADOUT => \N__6282\,
            PADIN => \N__6281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6274\,
            DIN => \N__6273\,
            DOUT => \N__6272\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6274\,
            PADOUT => \N__6273\,
            PADIN => \N__6272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4782\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6265\,
            DIN => \N__6264\,
            DOUT => \N__6263\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6265\,
            PADOUT => \N__6264\,
            PADIN => \N__6263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6256\,
            DIN => \N__6255\,
            DOUT => \N__6254\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6256\,
            PADOUT => \N__6255\,
            PADIN => \N__6254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6247\,
            DIN => \N__6246\,
            DOUT => \N__6245\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6247\,
            PADOUT => \N__6246\,
            PADIN => \N__6245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3771\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6238\,
            DIN => \N__6237\,
            DOUT => \N__6236\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6238\,
            PADOUT => \N__6237\,
            PADIN => \N__6236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2997\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6229\,
            DIN => \N__6228\,
            DOUT => \N__6227\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6229\,
            PADOUT => \N__6228\,
            PADIN => \N__6227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6220\,
            DIN => \N__6219\,
            DOUT => \N__6218\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6220\,
            PADOUT => \N__6219\,
            PADIN => \N__6218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6211\,
            DIN => \N__6210\,
            DOUT => \N__6209\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6211\,
            PADOUT => \N__6210\,
            PADIN => \N__6209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6202\,
            DIN => \N__6201\,
            DOUT => \N__6200\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6202\,
            PADOUT => \N__6201\,
            PADIN => \N__6200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6193\,
            DIN => \N__6192\,
            DOUT => \N__6191\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6193\,
            PADOUT => \N__6192\,
            PADIN => \N__6191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6184\,
            DIN => \N__6183\,
            DOUT => \N__6182\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6184\,
            PADOUT => \N__6183\,
            PADIN => \N__6182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6175\,
            DIN => \N__6174\,
            DOUT => \N__6173\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6175\,
            PADOUT => \N__6174\,
            PADIN => \N__6173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6166\,
            DIN => \N__6165\,
            DOUT => \N__6164\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6166\,
            PADOUT => \N__6165\,
            PADIN => \N__6164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6157\,
            DIN => \N__6156\,
            DOUT => \N__6155\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6157\,
            PADOUT => \N__6156\,
            PADIN => \N__6155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6148\,
            DIN => \N__6147\,
            DOUT => \N__6146\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6148\,
            PADOUT => \N__6147\,
            PADIN => \N__6146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3681\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6139\,
            DIN => \N__6138\,
            DOUT => \N__6137\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6139\,
            PADOUT => \N__6138\,
            PADIN => \N__6137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6130\,
            DIN => \N__6129\,
            DOUT => \N__6128\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6130\,
            PADOUT => \N__6129\,
            PADIN => \N__6128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6121\,
            DIN => \N__6120\,
            DOUT => \N__6119\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6121\,
            PADOUT => \N__6120\,
            PADIN => \N__6119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6112\,
            DIN => \N__6111\,
            DOUT => \N__6110\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6112\,
            PADOUT => \N__6111\,
            PADIN => \N__6110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6103\,
            DIN => \N__6102\,
            DOUT => \N__6101\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6103\,
            PADOUT => \N__6102\,
            PADIN => \N__6101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6094\,
            DIN => \N__6093\,
            DOUT => \N__6092\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6094\,
            PADOUT => \N__6093\,
            PADIN => \N__6092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6085\,
            DIN => \N__6084\,
            DOUT => \N__6083\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6085\,
            PADOUT => \N__6084\,
            PADIN => \N__6083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6076\,
            DIN => \N__6075\,
            DOUT => \N__6074\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6076\,
            PADOUT => \N__6075\,
            PADIN => \N__6074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6067\,
            DIN => \N__6066\,
            DOUT => \N__6065\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6067\,
            PADOUT => \N__6066\,
            PADIN => \N__6065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__6048\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__1403\ : IoInMux
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__6039\
        );

    \I__1401\ : Span12Mux_s1_v
    port map (
            O => \N__6039\,
            I => \N__6036\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__6036\,
            I => \N__6032\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6029\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__6032\,
            I => \TACK_OUTn\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6029\,
            I => \TACK_OUTn\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6017\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6014\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6011\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6006\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6006\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6017\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6014\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6011\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6006\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1387\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__5991\,
            I => \N__5987\
        );

    \I__1384\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5984\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__5987\,
            I => \N__5981\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__5984\,
            I => \N__5978\
        );

    \I__1381\ : Span4Mux_h
    port map (
            O => \N__5981\,
            I => \N__5962\
        );

    \I__1380\ : Span4Mux_v
    port map (
            O => \N__5978\,
            I => \N__5962\
        );

    \I__1379\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5959\
        );

    \I__1378\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5956\
        );

    \I__1377\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5949\
        );

    \I__1376\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5949\
        );

    \I__1375\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5949\
        );

    \I__1374\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5946\
        );

    \I__1373\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5941\
        );

    \I__1372\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5941\
        );

    \I__1371\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5938\
        );

    \I__1370\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5935\
        );

    \I__1369\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5932\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__5962\,
            I => \N__5925\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5925\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5956\,
            I => \N__5925\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__5949\,
            I => \N__5918\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5918\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5941\,
            I => \N__5918\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5915\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5935\,
            I => \N__5912\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__5932\,
            I => \N__5909\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__5925\,
            I => \N__5906\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__5918\,
            I => \N__5901\
        );

    \I__1357\ : Span4Mux_v
    port map (
            O => \N__5915\,
            I => \N__5901\
        );

    \I__1356\ : Span12Mux_h
    port map (
            O => \N__5912\,
            I => \N__5898\
        );

    \I__1355\ : Span12Mux_h
    port map (
            O => \N__5909\,
            I => \N__5895\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__5906\,
            I => \N__5890\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__5901\,
            I => \N__5890\
        );

    \I__1352\ : Span12Mux_v
    port map (
            O => \N__5898\,
            I => \N__5887\
        );

    \I__1351\ : Span12Mux_v
    port map (
            O => \N__5895\,
            I => \N__5884\
        );

    \I__1350\ : Span12Mux_h
    port map (
            O => \N__5890\,
            I => \N__5881\
        );

    \I__1349\ : Span12Mux_h
    port map (
            O => \N__5887\,
            I => \N__5878\
        );

    \I__1348\ : Span12Mux_h
    port map (
            O => \N__5884\,
            I => \N__5873\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__5881\,
            I => \N__5873\
        );

    \I__1346\ : Odrv12
    port map (
            O => \N__5878\,
            I => \RESETn_c\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__5873\,
            I => \RESETn_c\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__1343\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5858\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5855\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5848\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5848\
        );

    \I__1339\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5848\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5858\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5855\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5848\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5837\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5834\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5837\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__5834\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1331\ : CEMux
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__5826\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__5814\,
            I => \TACK_EN_i\
        );

    \I__1325\ : IoInMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__1323\ : IoSpan4Mux
    port map (
            O => \N__5805\,
            I => \N__5802\
        );

    \I__1322\ : Span4Mux_s3_v
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__5793\,
            I => \N_359_i\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__5790\,
            I => \N__5786\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__5789\,
            I => \N__5783\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5780\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5777\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5766\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5763\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5758\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5758\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5766\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5763\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__5758\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5745\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5745\,
            I => \U409_TRANSFER_ACK.N_132\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5735\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5726\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5726\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5726\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5726\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5735\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5726\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5707\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5707\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5707\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5707\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5702\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5702\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5707\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5702\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__5697\,
            I => \N__5690\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5680\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5680\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5680\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5680\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5675\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5675\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5680\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5675\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5656\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5656\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5656\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5651\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5651\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5656\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5651\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1270\ : SRMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5643\,
            I => \N__5636\
        );

    \I__1268\ : SRMux
    port map (
            O => \N__5642\,
            I => \N__5633\
        );

    \I__1267\ : SRMux
    port map (
            O => \N__5641\,
            I => \N__5630\
        );

    \I__1266\ : SRMux
    port map (
            O => \N__5640\,
            I => \N__5627\
        );

    \I__1265\ : SRMux
    port map (
            O => \N__5639\,
            I => \N__5624\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__5636\,
            I => \N__5619\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5633\,
            I => \N__5619\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5630\,
            I => \N__5615\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5627\,
            I => \N__5612\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5607\
        );

    \I__1259\ : Sp12to4
    port map (
            O => \N__5619\,
            I => \N__5607\
        );

    \I__1258\ : SRMux
    port map (
            O => \N__5618\,
            I => \N__5604\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__5615\,
            I => \N__5601\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__5612\,
            I => \N__5598\
        );

    \I__1255\ : Span12Mux_h
    port map (
            O => \N__5607\,
            I => \N__5593\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5593\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__5601\,
            I => \RESETn_c_i\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__5598\,
            I => \RESETn_c_i\
        );

    \I__1251\ : Odrv12
    port map (
            O => \N__5593\,
            I => \RESETn_c_i\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5582\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5579\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5582\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5579\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5570\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5567\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5564\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5567\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__5564\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__5559\,
            I => \N__5555\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5552\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5549\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5540\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5537\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5540\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5537\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__5532\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5523\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5516\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5516\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5516\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__5523\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5516\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__5511\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__5508\,
            I => \N__5504\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5500\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5495\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5495\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5500\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__5490\,
            I => \U409_TRANSFER_ACK.m9_am_cascade_\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5484\,
            I => \U409_TRANSFER_ACK.m9_bm\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5478\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5478\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5472\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__5463\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5456\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5452\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5449\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5446\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5452\,
            I => \N__5443\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__5449\,
            I => \N__5438\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5438\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__5443\,
            I => \N__5433\
        );

    \I__1200\ : Span4Mux_h
    port map (
            O => \N__5438\,
            I => \N__5433\
        );

    \I__1199\ : Span4Mux_h
    port map (
            O => \N__5433\,
            I => \N__5429\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5426\
        );

    \I__1197\ : Sp12to4
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5426\,
            I => \N__5420\
        );

    \I__1195\ : Span12Mux_v
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__1194\ : Sp12to4
    port map (
            O => \N__5420\,
            I => \N__5414\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__5417\,
            I => \TSn_c\
        );

    \I__1192\ : Odrv12
    port map (
            O => \N__5414\,
            I => \TSn_c\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5405\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5397\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5397\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__5397\,
            I => \N__5394\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__5394\,
            I => \N__5391\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__5391\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5384\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5381\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5384\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5381\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1180\ : IoInMux
    port map (
            O => \N__5376\,
            I => \N__5373\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5373\,
            I => \N__5369\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__5372\,
            I => \N__5366\
        );

    \I__1177\ : IoSpan4Mux
    port map (
            O => \N__5369\,
            I => \N__5362\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5359\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5356\
        );

    \I__1174\ : Span4Mux_s0_v
    port map (
            O => \N__5362\,
            I => \N__5351\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5346\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5346\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__5355\,
            I => \N__5343\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5354\,
            I => \N__5339\
        );

    \I__1169\ : Sp12to4
    port map (
            O => \N__5351\,
            I => \N__5335\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__5346\,
            I => \N__5332\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5327\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5327\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5324\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5321\
        );

    \I__1163\ : Span12Mux_v
    port map (
            O => \N__5335\,
            I => \N__5310\
        );

    \I__1162\ : Sp12to4
    port map (
            O => \N__5332\,
            I => \N__5310\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5310\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5324\,
            I => \N__5310\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5321\,
            I => \N__5310\
        );

    \I__1158\ : Span12Mux_v
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__5307\,
            I => \CLK40_IN_c\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5304\,
            I => \N__5294\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5291\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5282\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5282\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5282\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5282\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5275\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5275\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5275\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5291\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5282\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5275\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5254\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5254\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5254\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5254\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5249\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5249\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5254\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5229\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5229\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5229\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5229\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5222\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5222\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5222\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5222\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__5217\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5208\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5199\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5196\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5191\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5191\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5199\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5191\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1116\ : ClkMux
    port map (
            O => \N__5184\,
            I => \N__5175\
        );

    \I__1115\ : ClkMux
    port map (
            O => \N__5183\,
            I => \N__5175\
        );

    \I__1114\ : ClkMux
    port map (
            O => \N__5182\,
            I => \N__5175\
        );

    \I__1113\ : GlobalMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__1112\ : gio2CtrlBuf
    port map (
            O => \N__5172\,
            I => \CLK28_IN_c_g\
        );

    \I__1111\ : IoInMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__1109\ : Span12Mux_s4_v
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__1108\ : Span12Mux_v
    port map (
            O => \N__5160\,
            I => \N__5155\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5152\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5149\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__5155\,
            I => \CLKCIA_c\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5152\,
            I => \CLKCIA_c\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5149\,
            I => \CLKCIA_c\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__5142\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__5139\,
            I => \U409_TRANSFER_ACK.N_132_cascade_\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5131\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5126\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5126\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5131\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5112\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5112\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5112\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5106\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5085\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5085\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5085\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__5082\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__5079\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5070\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5065\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5065\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5062\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5070\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5065\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__5055\,
            I => \N__5051\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__5054\,
            I => \N__5047\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5041\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5041\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5036\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5036\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5036\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5023\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5023\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5018\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5018\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5003\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5000\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5003\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5000\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4995\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4989\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4989\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4982\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4979\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4982\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4979\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4971\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4964\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4961\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4964\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4961\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4944\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4944\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4939\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4939\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4930\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4930\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4930\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4930\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4944\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4930\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__4923\,
            I => \N__4915\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4902\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4902\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4902\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4902\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4902\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4895\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4895\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4895\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4902\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4895\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__4890\,
            I => \N__4885\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__4889\,
            I => \N__4877\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__4888\,
            I => \N__4874\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4871\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4862\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4862\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4862\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4862\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4855\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4855\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4855\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4871\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4855\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4845\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4835\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4832\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4832\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__997\ : ClkMux
    port map (
            O => \N__4827\,
            I => \N__4800\
        );

    \I__996\ : ClkMux
    port map (
            O => \N__4826\,
            I => \N__4800\
        );

    \I__995\ : ClkMux
    port map (
            O => \N__4825\,
            I => \N__4800\
        );

    \I__994\ : ClkMux
    port map (
            O => \N__4824\,
            I => \N__4800\
        );

    \I__993\ : ClkMux
    port map (
            O => \N__4823\,
            I => \N__4800\
        );

    \I__992\ : ClkMux
    port map (
            O => \N__4822\,
            I => \N__4800\
        );

    \I__991\ : ClkMux
    port map (
            O => \N__4821\,
            I => \N__4800\
        );

    \I__990\ : ClkMux
    port map (
            O => \N__4820\,
            I => \N__4800\
        );

    \I__989\ : ClkMux
    port map (
            O => \N__4819\,
            I => \N__4800\
        );

    \I__988\ : GlobalMux
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__987\ : gio2CtrlBuf
    port map (
            O => \N__4797\,
            I => \CLK6_c_g\
        );

    \I__986\ : InMux
    port map (
            O => \N__4794\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__985\ : InMux
    port map (
            O => \N__4791\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__984\ : InMux
    port map (
            O => \N__4788\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__983\ : InMux
    port map (
            O => \N__4785\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__982\ : IoInMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__980\ : Span12Mux_s1_v
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__979\ : Span12Mux_v
    port map (
            O => \N__4773\,
            I => \N__4769\
        );

    \I__978\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__4769\,
            I => \ROMENn_c\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4766\,
            I => \ROMENn_c\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4761\,
            I => \N__4756\
        );

    \I__974\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4753\
        );

    \I__973\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4748\
        );

    \I__972\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4748\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4753\,
            I => \N__4741\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4748\,
            I => \N__4741\
        );

    \I__969\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4736\
        );

    \I__968\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4736\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__4741\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__965\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4724\
        );

    \I__964\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4724\
        );

    \I__963\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4721\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4721\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__959\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4704\
        );

    \I__958\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4704\
        );

    \I__957\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4701\
        );

    \I__956\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4696\
        );

    \I__955\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4696\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4704\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4701\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4696\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__4689\,
            I => \N__4682\
        );

    \I__950\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4676\
        );

    \I__949\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4676\
        );

    \I__948\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4667\
        );

    \I__947\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4667\
        );

    \I__946\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4667\
        );

    \I__945\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4667\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4676\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4667\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__942\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4658\
        );

    \I__941\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4658\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4655\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__938\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4646\
        );

    \I__937\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4646\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4643\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__934\ : SRMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4631\
        );

    \I__932\ : SRMux
    port map (
            O => \N__4634\,
            I => \N__4628\
        );

    \I__931\ : Span4Mux_v
    port map (
            O => \N__4631\,
            I => \N__4621\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4628\,
            I => \N__4621\
        );

    \I__929\ : SRMux
    port map (
            O => \N__4627\,
            I => \N__4618\
        );

    \I__928\ : SRMux
    port map (
            O => \N__4626\,
            I => \N__4615\
        );

    \I__927\ : Span4Mux_h
    port map (
            O => \N__4621\,
            I => \N__4610\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4610\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4615\,
            I => \N__4607\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__4607\,
            I => \N__4601\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4604\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4601\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__920\ : IoInMux
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__918\ : Span4Mux_s2_v
    port map (
            O => \N__4590\,
            I => \N__4587\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__4584\,
            I => \CONSTANT_ONE_NET\
        );

    \I__915\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4578\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__913\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4571\
        );

    \I__912\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4568\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__4563\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__908\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4557\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__906\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4550\
        );

    \I__905\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4547\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__902\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4538\
        );

    \I__901\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4535\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4535\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__897\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4523\
        );

    \I__896\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4520\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4523\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4520\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__4515\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__892\ : IoInMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__890\ : Span4Mux_s2_v
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__889\ : Sp12to4
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__888\ : Span12Mux_h
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__887\ : Span12Mux_v
    port map (
            O => \N__4497\,
            I => \N__4493\
        );

    \I__886\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4490\
        );

    \I__885\ : Odrv12
    port map (
            O => \N__4493\,
            I => \TICK60_c\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4490\,
            I => \TICK60_c\
        );

    \I__883\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4481\
        );

    \I__882\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4478\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4481\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4478\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__879\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4469\
        );

    \I__878\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4469\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4466\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__874\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4454\
        );

    \I__873\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4451\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4454\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__870\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4442\
        );

    \I__869\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4439\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4442\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4439\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4434\,
            I => \N__4430\
        );

    \I__865\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4417\
        );

    \I__864\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4417\
        );

    \I__863\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4417\
        );

    \I__862\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4408\
        );

    \I__861\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4408\
        );

    \I__860\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4408\
        );

    \I__859\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4408\
        );

    \I__858\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4405\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4417\,
            I => \U409_TICK.TICK603_10\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4408\,
            I => \U409_TICK.TICK603_10\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4405\,
            I => \U409_TICK.TICK603_10\
        );

    \I__854\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4394\
        );

    \I__853\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4391\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4394\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4391\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__850\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4382\
        );

    \I__849\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4379\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4382\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4379\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__845\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4367\
        );

    \I__844\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4364\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4367\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__841\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4356\,
            I => \N__4352\
        );

    \I__839\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4349\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__4352\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4349\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__4344\,
            I => \N__4337\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__4343\,
            I => \N__4333\
        );

    \I__834\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4324\
        );

    \I__833\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4324\
        );

    \I__832\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4324\
        );

    \I__831\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4315\
        );

    \I__830\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4315\
        );

    \I__829\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4315\
        );

    \I__828\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4315\
        );

    \I__827\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4312\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4324\,
            I => \U409_TICK.TICK603_9\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4315\,
            I => \U409_TICK.TICK603_9\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4312\,
            I => \U409_TICK.TICK603_9\
        );

    \I__823\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4299\
        );

    \I__822\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4299\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__4293\,
            I => \CIA_ENABLEm\
        );

    \I__818\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4285\
        );

    \I__817\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4280\
        );

    \I__816\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4280\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4285\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4280\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__813\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4269\
        );

    \I__812\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4269\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4269\,
            I => \N__4265\
        );

    \I__810\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4262\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__4265\,
            I => \N__4259\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4262\,
            I => \N__4256\
        );

    \I__807\ : Sp12to4
    port map (
            O => \N__4259\,
            I => \N__4251\
        );

    \I__806\ : Span12Mux_h
    port map (
            O => \N__4256\,
            I => \N__4251\
        );

    \I__805\ : Odrv12
    port map (
            O => \N__4251\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4248\,
            I => \N__4243\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \N__4240\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__4246\,
            I => \N__4237\
        );

    \I__801\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4232\
        );

    \I__800\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4232\
        );

    \I__799\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4229\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4224\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4224\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__794\ : Span12Mux_h
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__4215\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__792\ : InMux
    port map (
            O => \N__4212\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__4209\,
            I => \N__4206\
        );

    \I__790\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4202\
        );

    \I__789\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4199\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4196\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4199\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__4196\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__785\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4188\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__783\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4182\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__780\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4173\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__778\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4166\
        );

    \I__777\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4163\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__774\ : InMux
    port map (
            O => \N__4158\,
            I => \N__4154\
        );

    \I__773\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4151\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4154\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4151\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__4146\,
            I => \N__4142\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__4145\,
            I => \N__4139\
        );

    \I__768\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4133\
        );

    \I__767\ : InMux
    port map (
            O => \N__4139\,
            I => \N__4133\
        );

    \I__766\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4130\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4133\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4130\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__763\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4121\
        );

    \I__762\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4121\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4118\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__759\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__758\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4109\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4106\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4101\,
            I => \N__4097\
        );

    \I__754\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4094\
        );

    \I__753\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4091\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4094\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4086\,
            I => \N__4082\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \N__4077\
        );

    \I__748\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4072\
        );

    \I__747\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4072\
        );

    \I__746\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4069\
        );

    \I__745\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4066\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4072\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4069\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4066\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__741\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4056\,
            I => \U409_TICK.TICK603_11\
        );

    \I__739\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4049\
        );

    \I__738\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4046\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4049\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4046\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__4041\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__734\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4034\
        );

    \I__733\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4034\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__730\ : InMux
    port map (
            O => \N__4026\,
            I => \N__4013\
        );

    \I__729\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4013\
        );

    \I__728\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4013\
        );

    \I__727\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4004\
        );

    \I__726\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4004\
        );

    \I__725\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4004\
        );

    \I__724\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4004\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4013\,
            I => \U409_TICK.TICK603_14\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U409_TICK.TICK603_14\
        );

    \I__721\ : InMux
    port map (
            O => \N__3999\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__720\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3992\
        );

    \I__719\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3989\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3992\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3989\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__716\ : InMux
    port map (
            O => \N__3984\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__715\ : InMux
    port map (
            O => \N__3981\,
            I => \bfn_11_7_0_\
        );

    \I__714\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3975\,
            I => \N__3971\
        );

    \I__712\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3968\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__3971\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3968\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__709\ : InMux
    port map (
            O => \N__3963\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__708\ : InMux
    port map (
            O => \N__3960\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__707\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3950\
        );

    \I__705\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3947\
        );

    \I__704\ : Odrv4
    port map (
            O => \N__3950\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3947\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__702\ : InMux
    port map (
            O => \N__3942\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__701\ : InMux
    port map (
            O => \N__3939\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__700\ : InMux
    port map (
            O => \N__3936\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__699\ : InMux
    port map (
            O => \N__3933\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__698\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3927\,
            I => \U409_TICK.TICK503_8\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__3924\,
            I => \U409_TICK.TICK503_11_cascade_\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__3921\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__694\ : IoInMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__692\ : Span12Mux_s10_v
    port map (
            O => \N__3912\,
            I => \N__3908\
        );

    \I__691\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3905\
        );

    \I__690\ : Odrv12
    port map (
            O => \N__3908\,
            I => \TICK50_c\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3905\,
            I => \TICK50_c\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__687\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3890\
        );

    \I__686\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3890\
        );

    \I__685\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3887\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3890\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3887\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__3882\,
            I => \N__3878\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3881\,
            I => \N__3873\
        );

    \I__680\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3870\
        );

    \I__679\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3865\
        );

    \I__678\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3865\
        );

    \I__677\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3862\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3870\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3865\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3862\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__673\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3851\
        );

    \I__672\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3848\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3851\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3848\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__669\ : InMux
    port map (
            O => \N__3843\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__668\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3836\
        );

    \I__667\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3833\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3836\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3833\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__664\ : InMux
    port map (
            O => \N__3828\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__663\ : InMux
    port map (
            O => \N__3825\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__662\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3818\
        );

    \I__661\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3815\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3818\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3815\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__658\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3807\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3807\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__656\ : InMux
    port map (
            O => \N__3804\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__654\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3795\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__652\ : InMux
    port map (
            O => \N__3792\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__651\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__648\ : Sp12to4
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__647\ : Span12Mux_h
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__3774\,
            I => \TACKn_in\
        );

    \I__645\ : IoInMux
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__643\ : Span4Mux_s1_v
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__642\ : Sp12to4
    port map (
            O => \N__3762\,
            I => \N__3758\
        );

    \I__641\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3755\
        );

    \I__640\ : Span12Mux_s11_h
    port map (
            O => \N__3758\,
            I => \N__3752\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3755\,
            I => \N__3749\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__3752\,
            I => \N__3746\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__3749\,
            I => \N__3743\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__3746\,
            I => \BUFENn_c\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3743\,
            I => \BUFENn_c\
        );

    \I__634\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3735\,
            I => \N__3732\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__3729\,
            I => \N__3726\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__3723\,
            I => \A_c_13\
        );

    \I__628\ : IoInMux
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__626\ : Span4Mux_s1_h
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__625\ : Sp12to4
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__624\ : Span12Mux_s9_v
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__622\ : Odrv12
    port map (
            O => \N__3702\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__621\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3696\,
            I => \N__3693\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__618\ : Sp12to4
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__617\ : Span12Mux_h
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__3684\,
            I => \A_c_12\
        );

    \I__615\ : IoInMux
    port map (
            O => \N__3681\,
            I => \N__3678\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__613\ : IoSpan4Mux
    port map (
            O => \N__3675\,
            I => \N__3672\
        );

    \I__612\ : Span4Mux_s3_h
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__611\ : Sp12to4
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__610\ : Span12Mux_h
    port map (
            O => \N__3666\,
            I => \N__3663\
        );

    \I__609\ : Odrv12
    port map (
            O => \N__3663\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3660\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__3657\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__605\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3647\
        );

    \I__604\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3644\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3647\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3644\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\
        );

    \I__601\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3634\
        );

    \I__600\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3631\
        );

    \I__599\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3628\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3634\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3631\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3628\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__3621\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\
        );

    \I__594\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3615\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11\
        );

    \I__592\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3605\
        );

    \I__591\ : InMux
    port map (
            O => \N__3611\,
            I => \N__3605\
        );

    \I__590\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3602\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3605\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3602\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3597\,
            I => \N__3592\
        );

    \I__586\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3586\
        );

    \I__585\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3586\
        );

    \I__584\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3581\
        );

    \I__583\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3581\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3586\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3581\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__580\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3567\
        );

    \I__579\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3567\
        );

    \I__578\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3564\
        );

    \I__577\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3559\
        );

    \I__576\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3559\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3567\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3564\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3559\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__3552\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_\
        );

    \I__571\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3546\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3546\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\
        );

    \I__569\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3535\
        );

    \I__568\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3530\
        );

    \I__567\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3530\
        );

    \I__566\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3527\
        );

    \I__565\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3522\
        );

    \I__564\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3522\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3535\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3530\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3527\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3522\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__559\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3507\
        );

    \I__558\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3504\
        );

    \I__557\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3499\
        );

    \I__556\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3499\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3507\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3504\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3499\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__552\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3489\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5\
        );

    \I__550\ : InMux
    port map (
            O => \N__3486\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__549\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3480\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__546\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3471\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3471\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__543\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3462\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__3459\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3456\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\
        );

    \I__539\ : InMux
    port map (
            O => \N__3453\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__538\ : InMux
    port map (
            O => \N__3450\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__537\ : InMux
    port map (
            O => \N__3447\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__536\ : InMux
    port map (
            O => \N__3444\,
            I => \bfn_10_9_0_\
        );

    \I__535\ : InMux
    port map (
            O => \N__3441\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__534\ : InMux
    port map (
            O => \N__3438\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__533\ : InMux
    port map (
            O => \N__3435\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__532\ : InMux
    port map (
            O => \N__3432\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__531\ : InMux
    port map (
            O => \N__3429\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__530\ : InMux
    port map (
            O => \N__3426\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__529\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3414\
        );

    \I__528\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3414\
        );

    \I__527\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3414\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3414\,
            I => \N__3411\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__3411\,
            I => \U409_ADDRESS_DECODE_un5_RAMSPACEn\
        );

    \I__524\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3398\
        );

    \I__523\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3398\
        );

    \I__522\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3398\
        );

    \I__521\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3395\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3398\,
            I => \N__3392\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3395\,
            I => \N__3389\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__3392\,
            I => \N__3385\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__3389\,
            I => \N__3382\
        );

    \I__516\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3379\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__3385\,
            I => \N__3371\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__3382\,
            I => \N__3371\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3379\,
            I => \N__3371\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__3378\,
            I => \N__3368\
        );

    \I__511\ : Span12Mux_h
    port map (
            O => \N__3371\,
            I => \N__3365\
        );

    \I__510\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3362\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__3365\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3362\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__506\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3351\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__3348\,
            I => \N__3345\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__3345\,
            I => \U409_ADDRESS_DECODE_HIROM\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__3342\,
            I => \N__3338\
        );

    \I__501\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3330\
        );

    \I__500\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3330\
        );

    \I__499\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3330\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3330\,
            I => \N__3327\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__496\ : Sp12to4
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__495\ : Span12Mux_h
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__494\ : Span12Mux_v
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__3315\,
            I => \OVL_c\
        );

    \I__492\ : InMux
    port map (
            O => \N__3312\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__491\ : InMux
    port map (
            O => \N__3309\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__490\ : InMux
    port map (
            O => \N__3306\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__489\ : InMux
    port map (
            O => \N__3303\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3300\,
            I => \N__3296\
        );

    \I__487\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3293\
        );

    \I__486\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3290\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3293\,
            I => \N__3286\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3290\,
            I => \N__3283\
        );

    \I__483\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3280\
        );

    \I__482\ : Odrv4
    port map (
            O => \N__3286\,
            I => \CIA_SPACEm_3\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3283\,
            I => \CIA_SPACEm_3\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3280\,
            I => \CIA_SPACEm_3\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__3273\,
            I => \N__3266\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__3272\,
            I => \N__3263\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__3271\,
            I => \N__3259\
        );

    \I__476\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3256\
        );

    \I__475\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3249\
        );

    \I__474\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3249\
        );

    \I__473\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3249\
        );

    \I__472\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3246\
        );

    \I__471\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3243\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3256\,
            I => \N__3240\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3249\,
            I => \N__3231\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3246\,
            I => \N__3231\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3243\,
            I => \N__3231\
        );

    \I__466\ : Sp12to4
    port map (
            O => \N__3240\,
            I => \N__3231\
        );

    \I__465\ : Span12Mux_v
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__464\ : Odrv12
    port map (
            O => \N__3228\,
            I => \A_c_22\
        );

    \I__463\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3221\
        );

    \I__462\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3217\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3214\
        );

    \I__460\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3211\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3217\,
            I => \N__3208\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__3214\,
            I => \N__3203\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3211\,
            I => \N__3203\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__3208\,
            I => \CIA_SPACEm_6\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__3203\,
            I => \CIA_SPACEm_6\
        );

    \I__454\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3195\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3195\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8\
        );

    \I__452\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3189\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3189\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__3186\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_\
        );

    \I__449\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__447\ : Span4Mux_h
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__3174\,
            I => \N__3171\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__3171\,
            I => \TT_c_1\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__443\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3160\
        );

    \I__442\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3157\
        );

    \I__441\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3154\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3160\,
            I => \N__3151\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3157\,
            I => \N__3146\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3154\,
            I => \N__3146\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__3151\,
            I => \N__3143\
        );

    \I__436\ : Span4Mux_v
    port map (
            O => \N__3146\,
            I => \N__3140\
        );

    \I__435\ : Sp12to4
    port map (
            O => \N__3143\,
            I => \N__3137\
        );

    \I__434\ : Span4Mux_h
    port map (
            O => \N__3140\,
            I => \N__3134\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__3137\,
            I => \A_c_31\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__3134\,
            I => \A_c_31\
        );

    \I__431\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3126\,
            I => \N__3123\
        );

    \I__429\ : Span12Mux_h
    port map (
            O => \N__3123\,
            I => \N__3120\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__3120\,
            I => \TT_c_0\
        );

    \I__427\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3114\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3114\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11\
        );

    \I__425\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3108\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3108\,
            I => \N__3104\
        );

    \I__423\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3101\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__3104\,
            I => \N__3098\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3101\,
            I => \N__3095\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3098\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__3095\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\
        );

    \I__418\ : IoInMux
    port map (
            O => \N__3090\,
            I => \N__3087\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__416\ : Span4Mux_s0_v
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__414\ : Span12Mux_s11_h
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__3075\,
            I => \N__3072\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__3072\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__411\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__409\ : Odrv12
    port map (
            O => \N__3063\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__408\ : InMux
    port map (
            O => \N__3060\,
            I => \N__3055\
        );

    \I__407\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3049\
        );

    \I__406\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3046\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3055\,
            I => \N__3043\
        );

    \I__404\ : InMux
    port map (
            O => \N__3054\,
            I => \N__3040\
        );

    \I__403\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3035\
        );

    \I__402\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3035\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3049\,
            I => \N__3032\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3046\,
            I => \N__3029\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__3043\,
            I => \N__3023\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3040\,
            I => \N__3023\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3035\,
            I => \N__3020\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__3032\,
            I => \N__3015\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__3029\,
            I => \N__3015\
        );

    \I__394\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3012\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__3023\,
            I => \N__3007\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__3020\,
            I => \N__3007\
        );

    \I__391\ : Sp12to4
    port map (
            O => \N__3015\,
            I => \N__3000\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3012\,
            I => \N__3000\
        );

    \I__389\ : Sp12to4
    port map (
            O => \N__3007\,
            I => \N__3000\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__3000\,
            I => \A_c_23\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__2997\,
            I => \N__2994\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__385\ : Span12Mux_s11_v
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__2988\,
            I => \PORTSIZE_0_i\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__2985\,
            I => \N__2981\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2984\,
            I => \N__2978\
        );

    \I__381\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2975\
        );

    \I__380\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2972\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2975\,
            I => \N__2969\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2966\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__2969\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__2966\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__2961\,
            I => \N__2958\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__373\ : IoSpan4Mux
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__372\ : Sp12to4
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__371\ : Span12Mux_s7_v
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__2946\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__369\ : InMux
    port map (
            O => \N__2943\,
            I => \N__2937\
        );

    \I__368\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2937\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2937\,
            I => \N__2933\
        );

    \I__366\ : InMux
    port map (
            O => \N__2936\,
            I => \N__2930\
        );

    \I__365\ : Span4Mux_h
    port map (
            O => \N__2933\,
            I => \N__2925\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2930\,
            I => \N__2925\
        );

    \I__363\ : Span4Mux_v
    port map (
            O => \N__2925\,
            I => \N__2922\
        );

    \I__362\ : Span4Mux_v
    port map (
            O => \N__2922\,
            I => \N__2919\
        );

    \I__361\ : Span4Mux_h
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__2916\,
            I => \A_c_28\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2913\,
            I => \U409_CIA.g0Z0Z_2_cascade_\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__2910\,
            I => \N__2906\
        );

    \I__357\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2900\
        );

    \I__356\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2900\
        );

    \I__355\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2897\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2900\,
            I => \N__2892\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2897\,
            I => \N__2892\
        );

    \I__352\ : Span4Mux_v
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__351\ : Span4Mux_v
    port map (
            O => \N__2889\,
            I => \N__2886\
        );

    \I__350\ : Sp12to4
    port map (
            O => \N__2886\,
            I => \N__2883\
        );

    \I__349\ : Odrv12
    port map (
            O => \N__2883\,
            I => \A_c_26\
        );

    \I__348\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2877\,
            I => \N__2873\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2876\,
            I => \N__2870\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__2873\,
            I => \N__2866\
        );

    \I__344\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2861\
        );

    \I__343\ : InMux
    port map (
            O => \N__2869\,
            I => \N__2861\
        );

    \I__342\ : Sp12to4
    port map (
            O => \N__2866\,
            I => \N__2856\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N__2856\
        );

    \I__340\ : Odrv12
    port map (
            O => \N__2856\,
            I => \A_c_27\
        );

    \I__339\ : InMux
    port map (
            O => \N__2853\,
            I => \N__2846\
        );

    \I__338\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2846\
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__2851\,
            I => \N__2843\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2846\,
            I => \N__2840\
        );

    \I__335\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2837\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__2840\,
            I => \N__2832\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2837\,
            I => \N__2832\
        );

    \I__332\ : Span4Mux_h
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__2826\,
            I => \A_c_24\
        );

    \I__329\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2820\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2820\,
            I => \U409_CIA.g0Z0Z_10\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2817\,
            I => \U409_CIA.g0Z0Z_8_cascade_\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2814\,
            I => \N__2810\
        );

    \I__325\ : InMux
    port map (
            O => \N__2813\,
            I => \N__2805\
        );

    \I__324\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2805\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__322\ : Span12Mux_s7_h
    port map (
            O => \N__2802\,
            I => \N__2799\
        );

    \I__321\ : Span12Mux_v
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__320\ : Odrv12
    port map (
            O => \N__2796\,
            I => \A_c_16\
        );

    \I__319\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2787\
        );

    \I__318\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2787\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__316\ : Span4Mux_v
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__315\ : Sp12to4
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__314\ : Span12Mux_v
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__2775\,
            I => \A_c_17\
        );

    \I__312\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__310\ : Span4Mux_h
    port map (
            O => \N__2766\,
            I => \N__2761\
        );

    \I__309\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2758\
        );

    \I__308\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2755\
        );

    \I__307\ : Span4Mux_v
    port map (
            O => \N__2761\,
            I => \N__2752\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2758\,
            I => \N__2747\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2755\,
            I => \N__2747\
        );

    \I__304\ : Odrv4
    port map (
            O => \N__2752\,
            I => \A_c_25\
        );

    \I__303\ : Odrv12
    port map (
            O => \N__2747\,
            I => \A_c_25\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__301\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2735\
        );

    \I__300\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2732\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2735\,
            I => \N__2727\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2732\,
            I => \N__2727\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__296\ : Sp12to4
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__295\ : Span12Mux_h
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__294\ : Span12Mux_v
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2715\,
            I => \A_c_18\
        );

    \I__292\ : InMux
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2709\,
            I => \U409_CIA.g0Z0Z_11\
        );

    \I__290\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2703\,
            I => \N__2698\
        );

    \I__288\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2693\
        );

    \I__287\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2693\
        );

    \I__286\ : Span4Mux_h
    port map (
            O => \N__2698\,
            I => \N__2690\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__2690\,
            I => \N__2684\
        );

    \I__283\ : Span4Mux_h
    port map (
            O => \N__2687\,
            I => \N__2681\
        );

    \I__282\ : Sp12to4
    port map (
            O => \N__2684\,
            I => \N__2676\
        );

    \I__281\ : Sp12to4
    port map (
            O => \N__2681\,
            I => \N__2676\
        );

    \I__280\ : Span12Mux_v
    port map (
            O => \N__2676\,
            I => \N__2673\
        );

    \I__279\ : Odrv12
    port map (
            O => \N__2673\,
            I => \A_c_19\
        );

    \I__278\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2666\
        );

    \I__277\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2663\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2666\,
            I => \N__2660\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2663\,
            I => \N__2656\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__2660\,
            I => \N__2653\
        );

    \I__273\ : InMux
    port map (
            O => \N__2659\,
            I => \N__2650\
        );

    \I__272\ : Span12Mux_v
    port map (
            O => \N__2656\,
            I => \N__2647\
        );

    \I__271\ : Sp12to4
    port map (
            O => \N__2653\,
            I => \N__2642\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2650\,
            I => \N__2642\
        );

    \I__269\ : Odrv12
    port map (
            O => \N__2647\,
            I => \A_c_20\
        );

    \I__268\ : Odrv12
    port map (
            O => \N__2642\,
            I => \A_c_20\
        );

    \I__267\ : InMux
    port map (
            O => \N__2637\,
            I => \N__2631\
        );

    \I__266\ : InMux
    port map (
            O => \N__2636\,
            I => \N__2626\
        );

    \I__265\ : InMux
    port map (
            O => \N__2635\,
            I => \N__2626\
        );

    \I__264\ : InMux
    port map (
            O => \N__2634\,
            I => \N__2623\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2631\,
            I => \N__2616\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2626\,
            I => \N__2616\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2623\,
            I => \N__2616\
        );

    \I__260\ : Span4Mux_v
    port map (
            O => \N__2616\,
            I => \N__2613\
        );

    \I__259\ : Span4Mux_h
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__258\ : Odrv4
    port map (
            O => \N__2610\,
            I => \A_c_21\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2607\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\
        );

    \I__256\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2601\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\
        );

    \I__254\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2591\
        );

    \I__253\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2591\
        );

    \I__252\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2588\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2591\,
            I => \N__2585\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2588\,
            I => \N__2582\
        );

    \I__249\ : Span4Mux_v
    port map (
            O => \N__2585\,
            I => \N__2577\
        );

    \I__248\ : Span4Mux_v
    port map (
            O => \N__2582\,
            I => \N__2577\
        );

    \I__247\ : Sp12to4
    port map (
            O => \N__2577\,
            I => \N__2574\
        );

    \I__246\ : Odrv12
    port map (
            O => \N__2574\,
            I => \A_c_30\
        );

    \I__245\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2565\
        );

    \I__244\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2565\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2565\,
            I => \N__2561\
        );

    \I__242\ : InMux
    port map (
            O => \N__2564\,
            I => \N__2558\
        );

    \I__241\ : Span4Mux_v
    port map (
            O => \N__2561\,
            I => \N__2553\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2558\,
            I => \N__2553\
        );

    \I__239\ : Span4Mux_h
    port map (
            O => \N__2553\,
            I => \N__2550\
        );

    \I__238\ : Span4Mux_v
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__237\ : Odrv4
    port map (
            O => \N__2547\,
            I => \A_c_29\
        );

    \I__236\ : ClkMux
    port map (
            O => \N__2544\,
            I => \N__2499\
        );

    \I__235\ : ClkMux
    port map (
            O => \N__2543\,
            I => \N__2499\
        );

    \I__234\ : ClkMux
    port map (
            O => \N__2542\,
            I => \N__2499\
        );

    \I__233\ : ClkMux
    port map (
            O => \N__2541\,
            I => \N__2499\
        );

    \I__232\ : ClkMux
    port map (
            O => \N__2540\,
            I => \N__2499\
        );

    \I__231\ : ClkMux
    port map (
            O => \N__2539\,
            I => \N__2499\
        );

    \I__230\ : ClkMux
    port map (
            O => \N__2538\,
            I => \N__2499\
        );

    \I__229\ : ClkMux
    port map (
            O => \N__2537\,
            I => \N__2499\
        );

    \I__228\ : ClkMux
    port map (
            O => \N__2536\,
            I => \N__2499\
        );

    \I__227\ : ClkMux
    port map (
            O => \N__2535\,
            I => \N__2499\
        );

    \I__226\ : ClkMux
    port map (
            O => \N__2534\,
            I => \N__2499\
        );

    \I__225\ : ClkMux
    port map (
            O => \N__2533\,
            I => \N__2499\
        );

    \I__224\ : ClkMux
    port map (
            O => \N__2532\,
            I => \N__2499\
        );

    \I__223\ : ClkMux
    port map (
            O => \N__2531\,
            I => \N__2499\
        );

    \I__222\ : ClkMux
    port map (
            O => \N__2530\,
            I => \N__2499\
        );

    \I__221\ : GlobalMux
    port map (
            O => \N__2499\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2543\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__2541\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            I => \N__2540\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__2537\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            I => \N__2535\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__2533\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2531\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2530\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            I => \N__2539\
        );

    \INVU409_TRANSFER_ACK.ROMENnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            I => \N__2536\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__2534\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2532\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2538\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__2544\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2542\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2634\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2670\,
            lcout => \CIA_SPACEm_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_9_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2853\,
            in1 => \N__2765\,
            in2 => \N__3300\,
            in3 => \N__2909\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2869\,
            in1 => \N__2852\,
            in2 => \N__2910\,
            in3 => \N__2764\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2570\,
            in1 => \N__2604\,
            in2 => \N__2607\,
            in3 => \N__2942\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_8_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2943\,
            in1 => \N__2598\,
            in2 => \N__2876\,
            in3 => \N__2571\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3164\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2597\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2564\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3270\,
            in1 => \N__2936\,
            in2 => \N__2913\,
            in3 => \N__2823\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2905\,
            in1 => \N__2880\,
            in2 => \N__2851\,
            in3 => \N__3163\,
            lcout => \U409_CIA.g0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3060\,
            in1 => \N__2793\,
            in2 => \_gnd_net_\,
            in3 => \N__5967\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2712\,
            in1 => \N__2813\,
            in2 => \N__2817\,
            in3 => \N__2702\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2701\,
            in1 => \N__2738\,
            in2 => \N__2814\,
            in3 => \N__2792\,
            lcout => \CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2659\,
            in1 => \N__2772\,
            in2 => \N__2742\,
            in3 => \N__2637\,
            lcout => \U409_CIA.g0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un5_RAMSPACEn_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3269\,
            in1 => \N__2636\,
            in2 => \_gnd_net_\,
            in3 => \N__3053\,
            lcout => \U409_ADDRESS_DECODE_un5_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3289\,
            in1 => \N__3052\,
            in2 => \N__3272\,
            in3 => \N__2706\,
            lcout => \U409_ADDRESS_DECODE_HIROM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__2669\,
            in1 => \N__3220\,
            in2 => \N__3273\,
            in3 => \N__2635\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3224\,
            in1 => \N__3262\,
            in2 => \N__3378\,
            in3 => \N__3299\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_10_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3054\,
            in1 => \N__5997\,
            in2 => \N__3271\,
            in3 => \N__3225\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_14_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3198\,
            in1 => \N__3192\,
            in2 => \N__3186\,
            in3 => \N__3117\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_11_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3183\,
            in1 => \N__5432\,
            in2 => \N__3168\,
            in3 => \N__3129\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3405\,
            in1 => \N__3059\,
            in2 => \_gnd_net_\,
            in3 => \N__3107\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3028\,
            in1 => \N__3388\,
            in2 => \_gnd_net_\,
            in3 => \N__3111\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__3069\,
            in1 => \N__3058\,
            in2 => \N__2984\,
            in3 => \N__5968\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__3421\,
            in1 => \N__3406\,
            in2 => \N__2985\,
            in3 => \N__3337\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__3407\,
            in1 => \_gnd_net_\,
            in2 => \N__3342\,
            in3 => \N__3422\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__3423\,
            in1 => \N__3408\,
            in2 => \N__3357\,
            in3 => \N__3341\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__5455\,
            in1 => \N__4662\,
            in2 => \N__5372\,
            in3 => \N__3543\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__4638\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3650\,
            in1 => \N__3512\,
            in2 => \_gnd_net_\,
            in3 => \N__4713\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__4627\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4138\,
            in2 => \N__4085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4157\,
            in2 => \_gnd_net_\,
            in3 => \N__3312\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__4824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4037\,
            in2 => \_gnd_net_\,
            in3 => \N__3309\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__4824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4101\,
            in3 => \N__3306\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4112\,
            in2 => \_gnd_net_\,
            in3 => \N__3303\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__4824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4355\,
            in2 => \_gnd_net_\,
            in3 => \N__3453\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4457\,
            in2 => \_gnd_net_\,
            in3 => \N__3450\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__4824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4385\,
            in2 => \_gnd_net_\,
            in3 => \N__3447\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4370\,
            in2 => \_gnd_net_\,
            in3 => \N__3444\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4484\,
            in2 => \_gnd_net_\,
            in3 => \N__3441\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__4826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4052\,
            in2 => \_gnd_net_\,
            in3 => \N__3438\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__4826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4169\,
            in2 => \_gnd_net_\,
            in3 => \N__3435\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__4826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4472\,
            in2 => \_gnd_net_\,
            in3 => \N__3432\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__4826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4397\,
            in2 => \_gnd_net_\,
            in3 => \N__3429\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4445\,
            in2 => \_gnd_net_\,
            in3 => \N__3426\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4125\,
            in2 => \_gnd_net_\,
            in3 => \N__3486\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4025\,
            in1 => \N__4341\,
            in2 => \N__4434\,
            in3 => \N__3483\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4827\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4342\,
            in1 => \N__4026\,
            in2 => \N__3477\,
            in3 => \N__4433\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4827\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4340\,
            in1 => \N__4024\,
            in2 => \N__3468\,
            in3 => \N__4429\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4827\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3575\,
            in1 => \N__3542\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__4626\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__3541\,
            in1 => \N__3576\,
            in2 => \N__3597\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__4626\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3574\,
            in2 => \_gnd_net_\,
            in3 => \N__3591\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3638\,
            in1 => \N__3611\,
            in2 => \N__3459\,
            in3 => \N__3492\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_2_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__5365\,
            in1 => \N__5459\,
            in2 => \N__3456\,
            in3 => \N__4649\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3618\,
            in2 => \N__3660\,
            in3 => \N__3612\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__4626\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__3513\,
            in2 => \N__3654\,
            in3 => \N__4715\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__4626\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3572\,
            in1 => \N__3596\,
            in2 => \_gnd_net_\,
            in3 => \N__3539\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U842_4_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4759\,
            in2 => \N__3657\,
            in3 => \N__4685\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIH6AR_6_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__3637\,
            in1 => \N__3510\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4747\,
            in1 => \N__4686\,
            in2 => \N__3621\,
            in3 => \N__4729\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4681\,
            in1 => \N__3538\,
            in2 => \N__4761\,
            in3 => \N__3610\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3595\,
            in1 => \N__3573\,
            in2 => \N__3552\,
            in3 => \N__3549\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_5_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3540\,
            in1 => \N__3511\,
            in2 => \N__4689\,
            in3 => \N__4746\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5990\,
            in1 => \N__3789\,
            in2 => \_gnd_net_\,
            in3 => \N__3761\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4305\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3738\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4304\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3877\,
            in1 => \_gnd_net_\,
            in2 => \N__3900\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4881\,
            in1 => \N__4914\,
            in2 => \N__3882\,
            in3 => \N__4953\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4913\,
            in1 => \N__4956\,
            in2 => \N__3801\,
            in3 => \N__4883\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3822\,
            in1 => \N__3840\,
            in2 => \_gnd_net_\,
            in3 => \N__3876\,
            lcout => \U409_TICK.TICK503_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__3810\,
            in1 => \N__4955\,
            in2 => \N__4923\,
            in3 => \N__4884\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3996\,
            in1 => \N__3855\,
            in2 => \N__4209\,
            in3 => \N__3896\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3930\,
            in1 => \N__3957\,
            in2 => \N__3924\,
            in3 => \N__3978\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__4882\,
            in1 => \N__3911\,
            in2 => \N__3921\,
            in3 => \N__4954\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3895\,
            in2 => \N__3881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3854\,
            in2 => \_gnd_net_\,
            in3 => \N__3843\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__4821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3839\,
            in2 => \_gnd_net_\,
            in3 => \N__3828\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__4821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5006\,
            in2 => \_gnd_net_\,
            in3 => \N__3825\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__4821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3821\,
            in2 => \_gnd_net_\,
            in3 => \N__3804\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4574\,
            in2 => \_gnd_net_\,
            in3 => \N__3792\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4526\,
            in2 => \_gnd_net_\,
            in3 => \N__3999\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__4821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3995\,
            in2 => \_gnd_net_\,
            in3 => \N__3984\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__4821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4838\,
            in2 => \_gnd_net_\,
            in3 => \N__3981\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3974\,
            in2 => \_gnd_net_\,
            in3 => \N__3963\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__4822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4553\,
            in2 => \_gnd_net_\,
            in3 => \N__3960\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3953\,
            in2 => \_gnd_net_\,
            in3 => \N__3942\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__4822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4985\,
            in2 => \_gnd_net_\,
            in3 => \N__3939\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4967\,
            in2 => \_gnd_net_\,
            in3 => \N__3936\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4541\,
            in2 => \_gnd_net_\,
            in3 => \N__3933\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4205\,
            in2 => \_gnd_net_\,
            in3 => \N__4212\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4822\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4021\,
            in1 => \N__4426\,
            in2 => \N__4343\,
            in3 => \N__4191\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4425\,
            in1 => \N__4020\,
            in2 => \N__4086\,
            in3 => \N__4332\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__4428\,
            in2 => \N__4344\,
            in3 => \N__4185\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4427\,
            in1 => \N__4022\,
            in2 => \N__4179\,
            in3 => \N__4336\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4146\,
            in3 => \N__4081\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4170\,
            in1 => \N__4158\,
            in2 => \N__4145\,
            in3 => \N__4124\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4113\,
            in1 => \N__4100\,
            in2 => \_gnd_net_\,
            in3 => \N__4080\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4059\,
            in1 => \N__4053\,
            in2 => \N__4041\,
            in3 => \N__4038\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__4496\,
            in1 => \N__4424\,
            in2 => \N__4515\,
            in3 => \N__4331\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4485\,
            in1 => \N__4473\,
            in2 => \N__4461\,
            in3 => \N__4446\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4398\,
            in1 => \N__4386\,
            in2 => \N__4374\,
            in3 => \N__4359\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5303\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4274\,
            in1 => \N__5202\,
            in2 => \N__4247\,
            in3 => \N__4288\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4275\,
            in1 => \N__5203\,
            in2 => \N__4248\,
            in3 => \N__4289\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4290\,
            in1 => \N__4268\,
            in2 => \N__4246\,
            in3 => \N__5205\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5639\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5529\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__5640\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101011101110"
        )
    port map (
            in0 => \N__4772\,
            in1 => \N__5475\,
            in2 => \N__5789\,
            in3 => \N__5481\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__5641\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4687\,
            in1 => \N__4731\,
            in2 => \N__4716\,
            in3 => \N__4760\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4634\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4730\,
            in1 => \N__4688\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4634\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__5573\,
            in1 => \N__4661\,
            in2 => \_gnd_net_\,
            in3 => \N__4650\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__4634\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4920\,
            in1 => \N__4951\,
            in2 => \N__4890\,
            in3 => \N__4581\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__4575\,
            in2 => \N__4842\,
            in3 => \N__4986\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4918\,
            in1 => \N__4949\,
            in2 => \N__4563\,
            in3 => \N__4560\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4968\,
            in1 => \N__4542\,
            in2 => \N__4530\,
            in3 => \N__5007\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4919\,
            in1 => \N__4880\,
            in2 => \N__4995\,
            in3 => \N__4992\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4950\,
            in1 => \N__4921\,
            in2 => \N__4888\,
            in3 => \N__4974\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4952\,
            in1 => \N__4922\,
            in2 => \N__4889\,
            in3 => \N__4848\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5263\,
            in2 => \N__5304\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5028\,
            in2 => \_gnd_net_\,
            in3 => \N__4794\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__5184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5238\,
            in2 => \_gnd_net_\,
            in3 => \N__4791\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5074\,
            in2 => \_gnd_net_\,
            in3 => \N__4788\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__5184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5050\,
            in2 => \_gnd_net_\,
            in3 => \N__4785\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__5240\,
            in1 => \N__5090\,
            in2 => \N__5103\,
            in3 => \N__5297\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101001100"
        )
    port map (
            in0 => \N__5298\,
            in1 => \N__5100\,
            in2 => \N__5094\,
            in3 => \N__5239\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5264\,
            in1 => \N__5075\,
            in2 => \N__5055\,
            in3 => \N__5029\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5302\,
            in2 => \_gnd_net_\,
            in3 => \N__5267\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5046\,
            in1 => \N__5073\,
            in2 => \_gnd_net_\,
            in3 => \N__5030\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5241\,
            in1 => \N__5299\,
            in2 => \_gnd_net_\,
            in3 => \N__5265\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5158\,
            in2 => \N__5082\,
            in3 => \N__5213\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__5013\,
            in1 => \N__5301\,
            in2 => \N__5079\,
            in3 => \N__5268\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5076\,
            in1 => \N__5243\,
            in2 => \N__5054\,
            in3 => \N__5031\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__5242\,
            in1 => \N__5300\,
            in2 => \_gnd_net_\,
            in3 => \N__5266\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__5204\,
            in1 => \N__5244\,
            in2 => \N__5217\,
            in3 => \N__5214\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5159\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5642\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5136\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5642\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110011"
        )
    port map (
            in0 => \N__5528\,
            in1 => \N__5109\,
            in2 => \N__5508\,
            in3 => \N__5739\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__5740\,
            in1 => \N__5971\,
            in2 => \N__5142\,
            in3 => \N__5772\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5135\,
            in1 => \N__5338\,
            in2 => \N__5121\,
            in3 => \N__5738\,
            lcout => \U409_TRANSFER_ACK.N_132\,
            ltout => \U409_TRANSFER_ACK.N_132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__5770\,
            in1 => \N__5503\,
            in2 => \N__5139\,
            in3 => \N__5526\,
            lcout => \U409_TRANSFER_ACK.m9_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5134\,
            in2 => \_gnd_net_\,
            in3 => \N__5117\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111110011"
        )
    port map (
            in0 => \N__5527\,
            in1 => \N__5769\,
            in2 => \N__5511\,
            in3 => \N__5507\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__5741\,
            in1 => \N__5970\,
            in2 => \N__5490\,
            in3 => \N__5487\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5663\,
            in1 => \N__5689\,
            in2 => \_gnd_net_\,
            in3 => \N__5716\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5717\,
            in1 => \_gnd_net_\,
            in2 => \N__5697\,
            in3 => \N__5664\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5469\,
            in1 => \N__5460\,
            in2 => \N__5355\,
            in3 => \N__5972\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5409\,
            in1 => \N__5387\,
            in2 => \_gnd_net_\,
            in3 => \N__5342\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__5408\,
            in1 => \N__5388\,
            in2 => \N__5354\,
            in3 => \N__5586\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5646\
        );

    \RESETn_ibuf_RNIM9SF_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__5696\,
            in1 => \N__5665\,
            in2 => \N__5790\,
            in3 => \N__5718\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5618\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000001100"
        )
    port map (
            in0 => \N__5771\,
            in1 => \N__5544\,
            in2 => \N__5751\,
            in3 => \N__5742\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5618\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5719\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5693\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5618\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5694\,
            in1 => \N__5666\,
            in2 => \_gnd_net_\,
            in3 => \N__5720\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5618\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100100000"
        )
    port map (
            in0 => \N__5721\,
            in1 => \N__5695\,
            in2 => \N__5670\,
            in3 => \N__5558\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5618\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5974\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5975\,
            in1 => \N__6022\,
            in2 => \_gnd_net_\,
            in3 => \N__5861\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5585\,
            in1 => \N__5574\,
            in2 => \N__5559\,
            in3 => \N__5543\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5863\,
            in1 => \N__5973\,
            in2 => \N__5532\,
            in3 => \N__6023\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6020\,
            in1 => \N__5864\,
            in2 => \_gnd_net_\,
            in3 => \N__5840\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001001100"
        )
    port map (
            in0 => \N__5976\,
            in1 => \N__6035\,
            in2 => \N__6048\,
            in3 => \N__6021\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__6024\,
            in1 => \N__5977\,
            in2 => \N__5868\,
            in3 => \N__5841\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__5829\,
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5823\,
            lcout => \N_359_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

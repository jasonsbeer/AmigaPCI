//iceprog D:\AmigaPCI\U111\U111_icecube\U111_icecube_Implmnt\sbt\outputs\bitmap\U111_TOP_bitmap.bin

module U111_TOP (
    input [1:0] A_040,
    input [1:0] SIZ,
    input CLK40_IN, RESETn, TS_CPUn, RnW, BGn, PORTSIZE, TACKn,

    output [1:0] A_AMIGA,
    output CLK40A, CLK40B, CLK40C, CLK80_CPU, CLKRAMA, CLKRAMB,
    output TSn, TAn, TBI_CPUn, TCI_CPUn, CPUBGn, BUFENn, BUFDIR, DMAn,

    inout [7:0] D_UU_040, //68040 DATA BUS
    inout [7:0] D_UM_040,
    inout [7:0] D_LM_040,
    inout [7:0] D_LL_040,

    inout [7:0] D_UU_AMIGA, //AMIGA DATA BUS
    inout [7:0] D_UM_AMIGA,
    inout [7:0] D_LM_AMIGA,
    inout [7:0] D_LL_AMIGA

    //testbench stuff
    //, input CLK80, CLK40

);

///////////////////////////////
// BUS AND PROCESSOR CLOCKS //
/////////////////////////////

//iCECUBE2 THROWS THIS ERROR, WHICH MUST BE ERRONEOUS?
//An input port (port CLK40_IN) is the target of an assignment - please check if this is intentional

//WE GENERATE THE 40MHz AND 80MHz CLOCKS HERE
wire CLK80;
wire CLK40;

assign CLK40A    = CLK40;
assign CLK40B    = CLK40;
assign CLK40C    = CLK40;
assign CLK80_CPU = CLK80;
assign CLKRAMA   = CLK80;
assign CLKRAMB   = CLK80;

SB_PLL40_2F_PAD #(
    .DIVR (4'b0000),
    .DIVF (7'b0001111),
    .DIVQ (3'b011),
    .FILTER_RANGE (3'b011),
    .FEEDBACK_PATH ("SIMPLE"),
    .PLLOUT_SELECT_PORTA ("GENCLK"),
    .PLLOUT_SELECT_PORTB ("GENCLK_HALF")
) pll (
    .LOCK           (),
    .RESETB         (1'b1),
    .PACKAGEPIN     (CLK40_IN),
    .PLLOUTGLOBALA  (CLK80),
    .PLLOUTGLOBALB  (CLK40)
);

//////////////
// BUFFERS //
////////////

wire CYCLE_EN = 1;
wire LBENn = 1;

U111_BUFFERS U111_BUFFERS (
    //INPUTS
    .RnW (RnW),
    .LBENn (LBENn),
    .CYCLE_EN (CYCLE_EN),
    .BGn (BGn),

    //OUTPUTS
    .CPUBGn (CPUBGn),
    .BUFENn (BUFENn),
    .BUFDIR (BUFDIR),
    .DMAn (DMAn)
);

//////////////////////////////////
// DATA TRANSFER STATE MACHINE //
////////////////////////////////

U111_CYCLE_SM U111_CYCLE_SM (
    //INPUTS
    .CLK80 (CLK80),
    .CLK40 (CLK40),
    .RESETn (RESETn),
    .TS_CPUn (TS_CPUn),
    .RnW (RnW),
    .PORTSIZE (PORTSIZE),
    .TACKn (TACKn),
    .SIZ (SIZ),
    .A_040 (A_040),

    //OUTPUTS
    .TAn (TAn),
    .TBI_CPUn (TBI_CPUn),
    .TCI_CPUn (TCI_CPUn),
    .A_AMIGA (A_AMIGA),
    .TSn (TSn),

    //INOUT
    .D_UU_040 (D_UU_040),
    .D_UM_040 (D_UM_040),
    .D_LM_040 (D_LM_040),
    .D_LL_040 (D_LL_040),
    .D_UU_AMIGA (D_UU_AMIGA),
    .D_UM_AMIGA (D_UM_AMIGA),
    .D_LM_AMIGA (D_LM_AMIGA),
    .D_LL_AMIGA (D_LL_AMIGA)
);


endmodule

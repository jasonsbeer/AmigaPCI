// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 19 2025 16:01:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_UU_AMIGA,
    D_LL_AMIGA,
    D_UM_AMIGA,
    D_LM_AMIGA,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    D_LL_040,
    A_AMIGA,
    A_040,
    SIZ,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    TBIn,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LL_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TEAn;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    input TBIn;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    inout TACKn;
    input BGn;

    wire N__13681;
    wire N__13665;
    wire N__13664;
    wire N__13663;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13647;
    wire N__13646;
    wire N__13645;
    wire N__13638;
    wire N__13637;
    wire N__13636;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13620;
    wire N__13619;
    wire N__13618;
    wire N__13611;
    wire N__13610;
    wire N__13609;
    wire N__13602;
    wire N__13601;
    wire N__13600;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13584;
    wire N__13583;
    wire N__13582;
    wire N__13575;
    wire N__13574;
    wire N__13573;
    wire N__13566;
    wire N__13565;
    wire N__13564;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13539;
    wire N__13538;
    wire N__13537;
    wire N__13530;
    wire N__13529;
    wire N__13528;
    wire N__13521;
    wire N__13520;
    wire N__13519;
    wire N__13512;
    wire N__13511;
    wire N__13510;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13494;
    wire N__13493;
    wire N__13492;
    wire N__13485;
    wire N__13484;
    wire N__13483;
    wire N__13476;
    wire N__13475;
    wire N__13474;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13458;
    wire N__13457;
    wire N__13456;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13440;
    wire N__13439;
    wire N__13438;
    wire N__13431;
    wire N__13430;
    wire N__13429;
    wire N__13422;
    wire N__13421;
    wire N__13420;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13404;
    wire N__13403;
    wire N__13402;
    wire N__13395;
    wire N__13394;
    wire N__13393;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13359;
    wire N__13358;
    wire N__13357;
    wire N__13350;
    wire N__13349;
    wire N__13348;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13332;
    wire N__13331;
    wire N__13330;
    wire N__13323;
    wire N__13322;
    wire N__13321;
    wire N__13314;
    wire N__13313;
    wire N__13312;
    wire N__13305;
    wire N__13304;
    wire N__13303;
    wire N__13296;
    wire N__13295;
    wire N__13294;
    wire N__13287;
    wire N__13286;
    wire N__13285;
    wire N__13278;
    wire N__13277;
    wire N__13276;
    wire N__13269;
    wire N__13268;
    wire N__13267;
    wire N__13260;
    wire N__13259;
    wire N__13258;
    wire N__13251;
    wire N__13250;
    wire N__13249;
    wire N__13242;
    wire N__13241;
    wire N__13240;
    wire N__13233;
    wire N__13232;
    wire N__13231;
    wire N__13224;
    wire N__13223;
    wire N__13222;
    wire N__13215;
    wire N__13214;
    wire N__13213;
    wire N__13206;
    wire N__13205;
    wire N__13204;
    wire N__13197;
    wire N__13196;
    wire N__13195;
    wire N__13188;
    wire N__13187;
    wire N__13186;
    wire N__13179;
    wire N__13178;
    wire N__13177;
    wire N__13170;
    wire N__13169;
    wire N__13168;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13143;
    wire N__13142;
    wire N__13141;
    wire N__13134;
    wire N__13133;
    wire N__13132;
    wire N__13125;
    wire N__13124;
    wire N__13123;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13098;
    wire N__13097;
    wire N__13096;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13062;
    wire N__13061;
    wire N__13060;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13026;
    wire N__13025;
    wire N__13024;
    wire N__13017;
    wire N__13016;
    wire N__13015;
    wire N__13008;
    wire N__13007;
    wire N__13006;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12945;
    wire N__12944;
    wire N__12943;
    wire N__12936;
    wire N__12935;
    wire N__12934;
    wire N__12927;
    wire N__12926;
    wire N__12925;
    wire N__12918;
    wire N__12917;
    wire N__12916;
    wire N__12909;
    wire N__12908;
    wire N__12907;
    wire N__12900;
    wire N__12899;
    wire N__12898;
    wire N__12891;
    wire N__12890;
    wire N__12889;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12873;
    wire N__12872;
    wire N__12871;
    wire N__12864;
    wire N__12863;
    wire N__12862;
    wire N__12855;
    wire N__12854;
    wire N__12853;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12721;
    wire N__12720;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12710;
    wire N__12709;
    wire N__12706;
    wire N__12705;
    wire N__12704;
    wire N__12701;
    wire N__12700;
    wire N__12699;
    wire N__12696;
    wire N__12695;
    wire N__12694;
    wire N__12693;
    wire N__12690;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12679;
    wire N__12678;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12670;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12604;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12596;
    wire N__12595;
    wire N__12594;
    wire N__12593;
    wire N__12592;
    wire N__12591;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12575;
    wire N__12570;
    wire N__12567;
    wire N__12562;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12547;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12541;
    wire N__12534;
    wire N__12529;
    wire N__12528;
    wire N__12527;
    wire N__12526;
    wire N__12521;
    wire N__12516;
    wire N__12509;
    wire N__12506;
    wire N__12505;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12498;
    wire N__12487;
    wire N__12476;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12434;
    wire N__12431;
    wire N__12430;
    wire N__12427;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12419;
    wire N__12416;
    wire N__12415;
    wire N__12414;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12407;
    wire N__12402;
    wire N__12399;
    wire N__12392;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12336;
    wire N__12335;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12305;
    wire N__12302;
    wire N__12295;
    wire N__12292;
    wire N__12285;
    wire N__12280;
    wire N__12277;
    wire N__12270;
    wire N__12263;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12241;
    wire N__12238;
    wire N__12233;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12196;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12172;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12163;
    wire N__12162;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12137;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12128;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12099;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__12074;
    wire N__12073;
    wire N__12072;
    wire N__12071;
    wire N__12070;
    wire N__12069;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12039;
    wire N__12036;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12032;
    wire N__12031;
    wire N__12030;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12012;
    wire N__12009;
    wire N__11998;
    wire N__11995;
    wire N__11992;
    wire N__11991;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11983;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11958;
    wire N__11957;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11932;
    wire N__11929;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11914;
    wire N__11913;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11884;
    wire N__11879;
    wire N__11876;
    wire N__11875;
    wire N__11872;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11830;
    wire N__11829;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11817;
    wire N__11816;
    wire N__11811;
    wire N__11804;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11785;
    wire N__11780;
    wire N__11777;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11754;
    wire N__11747;
    wire N__11746;
    wire N__11743;
    wire N__11742;
    wire N__11737;
    wire N__11730;
    wire N__11721;
    wire N__11716;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11655;
    wire N__11652;
    wire N__11647;
    wire N__11644;
    wire N__11633;
    wire N__11632;
    wire N__11631;
    wire N__11630;
    wire N__11629;
    wire N__11626;
    wire N__11621;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11606;
    wire N__11601;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11585;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11567;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11558;
    wire N__11555;
    wire N__11554;
    wire N__11553;
    wire N__11552;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11548;
    wire N__11545;
    wire N__11536;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11514;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11503;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11483;
    wire N__11482;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11476;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11465;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11408;
    wire N__11401;
    wire N__11398;
    wire N__11393;
    wire N__11390;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11376;
    wire N__11375;
    wire N__11374;
    wire N__11373;
    wire N__11370;
    wire N__11369;
    wire N__11368;
    wire N__11365;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11359;
    wire N__11358;
    wire N__11355;
    wire N__11350;
    wire N__11349;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11321;
    wire N__11316;
    wire N__11309;
    wire N__11308;
    wire N__11305;
    wire N__11298;
    wire N__11289;
    wire N__11280;
    wire N__11275;
    wire N__11264;
    wire N__11257;
    wire N__11254;
    wire N__11249;
    wire N__11246;
    wire N__11241;
    wire N__11234;
    wire N__11233;
    wire N__11232;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11180;
    wire N__11177;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11161;
    wire N__11152;
    wire N__11147;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11127;
    wire N__11124;
    wire N__11117;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11107;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11093;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11089;
    wire N__11088;
    wire N__11087;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11079;
    wire N__11076;
    wire N__11071;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11057;
    wire N__11054;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11022;
    wire N__11017;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11008;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10980;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10931;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10914;
    wire N__10903;
    wire N__10888;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10864;
    wire N__10863;
    wire N__10860;
    wire N__10853;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10842;
    wire N__10841;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10829;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10796;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10788;
    wire N__10785;
    wire N__10774;
    wire N__10771;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10742;
    wire N__10739;
    wire N__10734;
    wire N__10727;
    wire N__10724;
    wire N__10717;
    wire N__10710;
    wire N__10705;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10667;
    wire N__10660;
    wire N__10657;
    wire N__10650;
    wire N__10645;
    wire N__10640;
    wire N__10631;
    wire N__10628;
    wire N__10627;
    wire N__10626;
    wire N__10625;
    wire N__10624;
    wire N__10623;
    wire N__10622;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10615;
    wire N__10614;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10593;
    wire N__10592;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10588;
    wire N__10587;
    wire N__10586;
    wire N__10585;
    wire N__10584;
    wire N__10583;
    wire N__10582;
    wire N__10581;
    wire N__10580;
    wire N__10579;
    wire N__10578;
    wire N__10577;
    wire N__10576;
    wire N__10575;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10448;
    wire N__10445;
    wire N__10444;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10438;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10434;
    wire N__10433;
    wire N__10432;
    wire N__10431;
    wire N__10430;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10424;
    wire N__10423;
    wire N__10422;
    wire N__10421;
    wire N__10420;
    wire N__10419;
    wire N__10418;
    wire N__10417;
    wire N__10416;
    wire N__10415;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10409;
    wire N__10408;
    wire N__10407;
    wire N__10406;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10315;
    wire N__10314;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10310;
    wire N__10309;
    wire N__10308;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10304;
    wire N__10303;
    wire N__10302;
    wire N__10301;
    wire N__10300;
    wire N__10299;
    wire N__10298;
    wire N__10297;
    wire N__10296;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10292;
    wire N__10291;
    wire N__10290;
    wire N__10289;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10285;
    wire N__10284;
    wire N__10283;
    wire N__10282;
    wire N__10281;
    wire N__10280;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10273;
    wire N__10272;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10266;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9625;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__9001;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8997;
    wire N__8994;
    wire N__8993;
    wire N__8988;
    wire N__8985;
    wire N__8984;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8976;
    wire N__8975;
    wire N__8974;
    wire N__8973;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8963;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8953;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8866;
    wire N__8861;
    wire N__8858;
    wire N__8851;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8821;
    wire N__8816;
    wire N__8813;
    wire N__8804;
    wire N__8801;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8785;
    wire N__8780;
    wire N__8775;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8763;
    wire N__8758;
    wire N__8751;
    wire N__8746;
    wire N__8737;
    wire N__8734;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8603;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8491;
    wire N__8488;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8450;
    wire N__8447;
    wire N__8446;
    wire N__8445;
    wire N__8444;
    wire N__8443;
    wire N__8442;
    wire N__8441;
    wire N__8440;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8427;
    wire N__8422;
    wire N__8417;
    wire N__8412;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8404;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8385;
    wire N__8384;
    wire N__8381;
    wire N__8374;
    wire N__8369;
    wire N__8368;
    wire N__8365;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7872;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7861;
    wire N__7858;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7702;
    wire N__7699;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7636;
    wire N__7633;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7537;
    wire N__7534;
    wire N__7533;
    wire N__7530;
    wire N__7525;
    wire N__7520;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7505;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7448;
    wire N__7447;
    wire N__7444;
    wire N__7443;
    wire N__7440;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7141;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6958;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6848;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6829;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6811;
    wire N__6806;
    wire N__6803;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6791;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6779;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6758;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6743;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6650;
    wire N__6647;
    wire N__6646;
    wire N__6645;
    wire N__6640;
    wire N__6637;
    wire N__6636;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6624;
    wire N__6617;
    wire N__6614;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6583;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6442;
    wire N__6441;
    wire N__6440;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6429;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6395;
    wire N__6394;
    wire N__6393;
    wire N__6392;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6379;
    wire N__6374;
    wire N__6369;
    wire N__6362;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6315;
    wire N__6314;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6302;
    wire N__6299;
    wire N__6292;
    wire N__6287;
    wire N__6286;
    wire N__6285;
    wire N__6282;
    wire N__6277;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6247;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6230;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6201;
    wire N__6198;
    wire N__6193;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6182;
    wire N__6179;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6167;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6139;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6115;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6091;
    wire N__6088;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6061;
    wire N__6060;
    wire N__6057;
    wire N__6056;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5987;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire TCIn_c;
    wire VCCG0;
    wire GNDG0;
    wire TAn_in;
    wire N_237_i;
    wire N_240_i;
    wire N_242_i;
    wire N_228_i;
    wire N_241_i;
    wire N_243_i;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_0 ;
    wire N_229_i;
    wire RESETn_c_i;
    wire N_231_i;
    wire N_220_i;
    wire N_230_i;
    wire N_232_i;
    wire N_222_i;
    wire N_221_i;
    wire N_233_i;
    wire N_234_i;
    wire N_235_i;
    wire N_213_i;
    wire N_223_i;
    wire N_224_i;
    wire N_217_i;
    wire N_227_i;
    wire N_226_i;
    wire N_236_i;
    wire N_239_i;
    wire N_238_i;
    wire WRITE_CYCLE_ACTIVE_rep24_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep25_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep28_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep27_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep26_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep30_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep16_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep29_i_ess;
    wire WRITE_CYCLE_ACTIVE_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep17_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep19_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep18_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep20_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep21_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep22_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep9_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep23_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep11_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep1_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep5_i_ess;
    wire N_215_i;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire D_LL_AMIGA_in_7;
    wire un2_D_LL_AMIGA_7;
    wire D_LL_040_in_2;
    wire D_UM_040_in_2;
    wire un1_D_UM_040_2;
    wire WRITE_CYCLE_ACTIVE_rep8_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep10_i_ess;
    wire D_LM_AMIGA_in_7;
    wire un2_D_LM_AMIGA_7;
    wire WRITE_CYCLE_ACTIVE_rep12_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep14_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep6_i_ess;
    wire N_218_i;
    wire D_UU_040_in_7;
    wire D_LM_040_in_7;
    wire un1_D_UU_040_7;
    wire N_219_i;
    wire D_LL_AMIGA_in_5;
    wire un2_D_LL_AMIGA_5;
    wire D_LM_AMIGA_in_1;
    wire un2_D_LM_AMIGA_1;
    wire WRITE_CYCLE_ACTIVE_rep15_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep3_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep7_i_ess;
    wire D_LM_AMIGA_in_3;
    wire un2_D_LM_AMIGA_3;
    wire D_LM_AMIGA_in_5;
    wire un2_D_LM_AMIGA_5;
    wire N_214_i;
    wire D_UU_040_in_1;
    wire D_LM_040_in_1;
    wire un1_D_UU_040_1;
    wire WRITE_CYCLE_ACTIVE_rep0_i_ess;
    wire N_212_i;
    wire WRITE_CYCLE_ACTIVE_rep4_i_ess;
    wire N_216_i;
    wire WRITE_CYCLE_ACTIVE_rep2_i_ess;
    wire N_225_i;
    wire LBENn_c_i;
    wire D_LL_AMIGA_in_0;
    wire un2_D_LL_AMIGA_0;
    wire D_LM_AMIGA_in_2;
    wire un2_D_LM_AMIGA_2;
    wire WRITE_CYCLE_ACTIVE_rep13_i_ess;
    wire D_UU_040_in_5;
    wire D_LM_040_in_5;
    wire un1_D_UU_040_5;
    wire D_LL_AMIGA_in_6;
    wire un2_D_LL_AMIGA_6;
    wire D_LM_AMIGA_in_0;
    wire un2_D_LM_AMIGA_0;
    wire D_LL_AMIGA_in_3;
    wire un2_D_LL_AMIGA_3;
    wire D_LL_AMIGA_in_4;
    wire un2_D_LL_AMIGA_4;
    wire D_LM_AMIGA_in_4;
    wire un2_D_LM_AMIGA_4;
    wire CONSTANT_ONE_NET;
    wire LBENn_c_i_0;
    wire D_LL_AMIGA_in_1;
    wire un2_D_LL_AMIGA_1;
    wire A_040_c_1;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ;
    wire \U111_CYCLE_SM.N_148_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire un1_D_UU_AMIGA_1;
    wire D_LL_AMIGA_in_2;
    wire un2_D_LL_AMIGA_2;
    wire \U111_CYCLE_SM.TS_ENZ0Z6 ;
    wire \U111_CYCLE_SM.N_158_cascade_ ;
    wire \U111_CYCLE_SM.N_130_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.TS_EN_6 ;
    wire \U111_CYCLE_SM.N_160_cascade_ ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U111_CYCLE_SM.PORT_MISMATCH_2_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire \U111_CYCLE_SM.N_142_0 ;
    wire TBIn_c;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ;
    wire \U111_CYCLE_SM.N_149 ;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire \U111_CYCLE_SM.N_132_0_cascade_ ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_ ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2 ;
    wire TACKn_in;
    wire TEAn_c;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire D_LM_AMIGA_in_6;
    wire un2_D_LM_AMIGA_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire D_UM_AMIGA_in_5;
    wire un1_D_UM_AMIGA_5;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire D_UU_AMIGA_in_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire \U111_CYCLE_SM.FLIP_WORD_2 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire \U111_CYCLE_SM.N_160 ;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire un1_D_UM_AMIGA_0;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire PORTSIZE_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire un1_D_UM_AMIGA_2;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire un1_D_UM_AMIGA_6;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire \U111_CYCLE_SM.N_159_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire TAn_1_i;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire D_UM_AMIGA_in_3;
    wire un1_D_UM_AMIGA_3;
    wire D_UM_AMIGA_in_4;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire un1_D_UM_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire D_UU_AMIGA_in_6;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire un1_D_UU_AMIGA_6;
    wire D_LM_040_in_6;
    wire D_UU_040_in_6;
    wire un1_D_UU_040_6;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire D_LL_040_in_4;
    wire D_UM_040_in_4;
    wire un1_D_UM_040_4;
    wire D_UM_040_in_5;
    wire D_LL_040_in_5;
    wire un1_D_UM_040_5;
    wire D_LL_040_in_1;
    wire D_UM_040_in_1;
    wire un1_D_UM_040_1;
    wire D_LM_040_in_2;
    wire D_UU_040_in_2;
    wire un1_D_UU_040_2;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_UM_040_in_3;
    wire D_LL_040_in_3;
    wire un1_D_UM_040_3;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire D_LL_040_in_7;
    wire D_UM_040_in_7;
    wire un1_D_UM_040_7;
    wire READ_CYCLE_ACTIVE_rep4_i_ess;
    wire N_184_i;
    wire READ_CYCLE_ACTIVE_rep2_i_ess;
    wire N_182_i;
    wire READ_CYCLE_ACTIVE_rep0_i_ess;
    wire N_180_i;
    wire READ_CYCLE_ACTIVE_rep7_i_ess;
    wire N_187_i;
    wire READ_CYCLE_ACTIVE_rep6_i_ess;
    wire N_186_i;
    wire N_207_i;
    wire N_205_i;
    wire READ_CYCLE_ACTIVE_rep27_i_ess;
    wire READ_CYCLE_ACTIVE_rep25_i_ess;
    wire N_196_i;
    wire READ_CYCLE_ACTIVE_rep16_i_ess;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire READ_CYCLE_ACTIVE_rep5_i_ess;
    wire N_185_i;
    wire READ_CYCLE_ACTIVE_rep13_i_ess;
    wire N_193_i;
    wire N_208_i;
    wire READ_CYCLE_ACTIVE_rep28_i_ess;
    wire N_204_i;
    wire READ_CYCLE_ACTIVE_rep30_i_ess;
    wire N_210_i;
    wire N_206_i;
    wire N_209_i;
    wire READ_CYCLE_ACTIVE_rep29_i_ess;
    wire READ_CYCLE_ACTIVE_rep24_i_ess;
    wire READ_CYCLE_ACTIVE_rep26_i_ess;
    wire N_197_i;
    wire N_211_i;
    wire N_198_i;
    wire N_199_i;
    wire READ_CYCLE_ACTIVE_rep31_i_ess;
    wire READ_CYCLE_ACTIVE_rep19_i_ess;
    wire READ_CYCLE_ACTIVE_rep18_i_ess;
    wire READ_CYCLE_ACTIVE_rep17_i_ess;
    wire N_200_i;
    wire N_188_i;
    wire READ_CYCLE_ACTIVE_rep21_i_ess;
    wire N_201_i;
    wire READ_CYCLE_ACTIVE_rep20_i_ess;
    wire READ_CYCLE_ACTIVE_rep8_i_ess;
    wire N_190_i;
    wire N_194_i;
    wire READ_CYCLE_ACTIVE_rep14_i_ess;
    wire READ_CYCLE_ACTIVE_rep10_i_ess;
    wire READ_CYCLE_ACTIVE_rep22_i_ess;
    wire N_202_i;
    wire READ_CYCLE_ACTIVE_rep23_i_ess;
    wire N_203_i;
    wire READ_CYCLE_ACTIVE_rep9_i_ess;
    wire N_189_i;
    wire READ_CYCLE_ACTIVE_rep11_i_ess;
    wire N_191_i;
    wire READ_CYCLE_ACTIVE_rep15_i_ess;
    wire N_195_i;
    wire RnW_c;
    wire TS_CPUn_c;
    wire LBENn_c;
    wire BGn_c;
    wire CLK40;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_g_0 ;
    wire RESETn_c_i_g;
    wire READ_CYCLE_ACTIVE_rep1_i_ess;
    wire N_181_i;
    wire READ_CYCLE_ACTIVE_rep12_i_ess;
    wire N_192_i;
    wire READ_CYCLE_ACTIVE_rep3_i_ess;
    wire N_183_i;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__5485),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__13681));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__13681),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__13665),
            .DIN(N__13664),
            .DOUT(N__13663),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__13665),
            .PADOUT(N__13664),
            .PADIN(N__13663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__13656),
            .DIN(N__13655),
            .DOUT(N__13654),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__13656),
            .PADOUT(N__13655),
            .PADIN(N__13654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7811),
            .DIN0(TAn_in),
            .DOUT0(N__6287),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__13647),
            .DIN(N__13646),
            .DOUT(N__13645),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__13647),
            .PADOUT(N__13646),
            .PADIN(N__13645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4184),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__7988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__13638),
            .DIN(N__13637),
            .DOUT(N__13636),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__13638),
            .PADOUT(N__13637),
            .PADIN(N__13636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9527),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__8333),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__13629),
            .DIN(N__13628),
            .DOUT(N__13627),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__13629),
            .PADOUT(N__13628),
            .PADIN(N__13627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__13620),
            .DIN(N__13619),
            .DOUT(N__13618),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__13620),
            .PADOUT(N__13619),
            .PADIN(N__13618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4448),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__9044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__13611),
            .DIN(N__13610),
            .DOUT(N__13609),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__13611),
            .PADOUT(N__13610),
            .PADIN(N__13609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__13602),
            .DIN(N__13601),
            .DOUT(N__13600),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__13602),
            .PADOUT(N__13601),
            .PADIN(N__13600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4280),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__9245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__13593),
            .DIN(N__13592),
            .DOUT(N__13591),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__13593),
            .PADOUT(N__13592),
            .PADIN(N__13591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10082),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__5000),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__13584),
            .DIN(N__13583),
            .DOUT(N__13582),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__13584),
            .PADOUT(N__13583),
            .PADIN(N__13582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__13575),
            .DIN(N__13574),
            .DOUT(N__13573),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__13575),
            .PADOUT(N__13574),
            .PADIN(N__13573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12776),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__6569),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__13566),
            .DIN(N__13565),
            .DOUT(N__13564),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__13566),
            .PADOUT(N__13565),
            .PADIN(N__13564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__13557),
            .DIN(N__13556),
            .DOUT(N__13555),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__13557),
            .PADOUT(N__13556),
            .PADIN(N__13555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4865),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__4883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__13548),
            .DIN(N__13547),
            .DOUT(N__13546),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__13548),
            .PADOUT(N__13547),
            .PADIN(N__13546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12718),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__13539),
            .DIN(N__13538),
            .DOUT(N__13537),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__13539),
            .PADOUT(N__13538),
            .PADIN(N__13537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__13530),
            .DIN(N__13529),
            .DOUT(N__13528),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__13530),
            .PADOUT(N__13529),
            .PADIN(N__13528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__13521),
            .DIN(N__13520),
            .DOUT(N__13519),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__13521),
            .PADOUT(N__13520),
            .PADIN(N__13519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9731),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__5423),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__13512),
            .DIN(N__13511),
            .DOUT(N__13510),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__13512),
            .PADOUT(N__13511),
            .PADIN(N__13510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10157),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__5933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__13503),
            .DIN(N__13502),
            .DOUT(N__13501),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__13503),
            .PADOUT(N__13502),
            .PADIN(N__13501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4085),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__5062),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__13494),
            .DIN(N__13493),
            .DOUT(N__13492),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__13494),
            .PADOUT(N__13493),
            .PADIN(N__13492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9929),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__5249),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__13485),
            .DIN(N__13484),
            .DOUT(N__13483),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__13485),
            .PADOUT(N__13484),
            .PADIN(N__13483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5450),
            .DIN0(TACKn_in),
            .DOUT0(N__4208),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__13476),
            .DIN(N__13475),
            .DOUT(N__13474),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__13476),
            .PADOUT(N__13475),
            .PADIN(N__13474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10004),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__7418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__13467),
            .DIN(N__13466),
            .DOUT(N__13465),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__13467),
            .PADOUT(N__13466),
            .PADIN(N__13465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__13458),
            .DIN(N__13457),
            .DOUT(N__13456),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__13458),
            .PADOUT(N__13457),
            .PADIN(N__13456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4334),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__4693),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__13449),
            .DIN(N__13448),
            .DOUT(N__13447),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__13449),
            .PADOUT(N__13448),
            .PADIN(N__13447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5102),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__9458),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TEAn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__13440),
            .DIN(N__13439),
            .DOUT(N__13438),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__13440),
            .PADOUT(N__13439),
            .PADIN(N__13438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__13431),
            .DIN(N__13430),
            .DOUT(N__13429),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__13431),
            .PADOUT(N__13430),
            .PADIN(N__13429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__13422),
            .DIN(N__13421),
            .DOUT(N__13420),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__13422),
            .PADOUT(N__13421),
            .PADIN(N__13420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5486),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__13413),
            .DIN(N__13412),
            .DOUT(N__13411),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__13413),
            .PADOUT(N__13412),
            .PADIN(N__13411),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9797),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__5666),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__13404),
            .DIN(N__13403),
            .DOUT(N__13402),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__13404),
            .PADOUT(N__13403),
            .PADIN(N__13402),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4127),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__8057),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__13395),
            .DIN(N__13394),
            .DOUT(N__13393),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__13395),
            .PADOUT(N__13394),
            .PADIN(N__13393),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4298),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__9134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__13386),
            .DIN(N__13385),
            .DOUT(N__13384),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__13386),
            .PADOUT(N__13385),
            .PADIN(N__13384),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9593),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__6884),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__13377),
            .DIN(N__13376),
            .DOUT(N__13375),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__13377),
            .PADOUT(N__13376),
            .PADIN(N__13375),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4289),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__9511),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__13368),
            .DIN(N__13367),
            .DOUT(N__13366),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__13368),
            .PADOUT(N__13367),
            .PADIN(N__13366),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6529),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__13359),
            .DIN(N__13358),
            .DOUT(N__13357),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__13359),
            .PADOUT(N__13358),
            .PADIN(N__13357),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9749),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__5585),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__13350),
            .DIN(N__13349),
            .DOUT(N__13348),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__13350),
            .PADOUT(N__13349),
            .PADIN(N__13348),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9962),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__5228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_obuf_iopad (
            .OE(N__13341),
            .DIN(N__13340),
            .DOUT(N__13339),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__13341),
            .PADOUT(N__13340),
            .PADIN(N__13339),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5801),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__13332),
            .DIN(N__13331),
            .DOUT(N__13330),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__13332),
            .PADOUT(N__13331),
            .PADIN(N__13330),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4400),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__8657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__13323),
            .DIN(N__13322),
            .DOUT(N__13321),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__13323),
            .PADOUT(N__13322),
            .PADIN(N__13321),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4478),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__4919),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__13314),
            .DIN(N__13313),
            .DOUT(N__13312),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__13314),
            .PADOUT(N__13313),
            .PADIN(N__13312),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__13305),
            .DIN(N__13304),
            .DOUT(N__13303),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__13305),
            .PADOUT(N__13304),
            .PADIN(N__13303),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4751),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__13296),
            .DIN(N__13295),
            .DOUT(N__13294),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__13296),
            .PADOUT(N__13295),
            .PADIN(N__13294),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10055),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__5510),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__13287),
            .DIN(N__13286),
            .DOUT(N__13285),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__13287),
            .PADOUT(N__13286),
            .PADIN(N__13285),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12734),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__7097),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__13278),
            .DIN(N__13277),
            .DOUT(N__13276),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__13278),
            .PADOUT(N__13277),
            .PADIN(N__13276),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__13269),
            .DIN(N__13268),
            .DOUT(N__13267),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__13269),
            .PADOUT(N__13268),
            .PADIN(N__13267),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4463),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__5399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__13260),
            .DIN(N__13259),
            .DOUT(N__13258),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__13260),
            .PADOUT(N__13259),
            .PADIN(N__13258),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9666),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__13251),
            .DIN(N__13250),
            .DOUT(N__13249),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__13251),
            .PADOUT(N__13250),
            .PADIN(N__13249),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10040),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__7559),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__13242),
            .DIN(N__13241),
            .DOUT(N__13240),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__13242),
            .PADOUT(N__13241),
            .PADIN(N__13240),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4367),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__9173),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__13233),
            .DIN(N__13232),
            .DOUT(N__13231),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__13233),
            .PADOUT(N__13232),
            .PADIN(N__13231),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5351),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__9206),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__13224),
            .DIN(N__13223),
            .DOUT(N__13222),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__13224),
            .PADOUT(N__13223),
            .PADIN(N__13222),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9545),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__6953),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__13215),
            .DIN(N__13214),
            .DOUT(N__13213),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__13215),
            .PADOUT(N__13214),
            .PADIN(N__13213),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam BGn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD BGn_ibuf_iopad (
            .OE(N__13206),
            .DIN(N__13205),
            .DOUT(N__13204),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__13206),
            .PADOUT(N__13205),
            .PADIN(N__13204),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__13197),
            .DIN(N__13196),
            .DOUT(N__13195),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__13197),
            .PADOUT(N__13196),
            .PADIN(N__13195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9821),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__5282),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__13188),
            .DIN(N__13187),
            .DOUT(N__13186),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__13188),
            .PADOUT(N__13187),
            .PADIN(N__13186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4268),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__4631),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__13179),
            .DIN(N__13178),
            .DOUT(N__13177),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__13179),
            .PADOUT(N__13178),
            .PADIN(N__13177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9572),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__7022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__13170),
            .DIN(N__13169),
            .DOUT(N__13168),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__13170),
            .PADOUT(N__13169),
            .PADIN(N__13168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__13161),
            .DIN(N__13160),
            .DOUT(N__13159),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__13161),
            .PADOUT(N__13160),
            .PADIN(N__13159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__13152),
            .DIN(N__13151),
            .DOUT(N__13150),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__13152),
            .PADOUT(N__13151),
            .PADIN(N__13150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4142),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__9416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__13143),
            .DIN(N__13142),
            .DOUT(N__13141),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__13143),
            .PADOUT(N__13142),
            .PADIN(N__13141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6010),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__13134),
            .DIN(N__13133),
            .DOUT(N__13132),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__13134),
            .PADOUT(N__13133),
            .PADIN(N__13132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9642),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__13125),
            .DIN(N__13124),
            .DOUT(N__13123),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__13125),
            .PADOUT(N__13124),
            .PADIN(N__13123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9914),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__5165),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__13116),
            .DIN(N__13115),
            .DOUT(N__13114),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__13116),
            .PADOUT(N__13115),
            .PADIN(N__13114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4238),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__5744),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__13107),
            .DIN(N__13106),
            .DOUT(N__13105),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__13107),
            .PADOUT(N__13106),
            .PADIN(N__13105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10103),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__6473),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__13098),
            .DIN(N__13097),
            .DOUT(N__13096),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__13098),
            .PADOUT(N__13097),
            .PADIN(N__13096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9857),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__7169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__13089),
            .DIN(N__13088),
            .DOUT(N__13087),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__13089),
            .PADOUT(N__13088),
            .PADIN(N__13087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4352),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__9092),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__13080),
            .DIN(N__13079),
            .DOUT(N__13078),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__13080),
            .PADOUT(N__13079),
            .PADIN(N__13078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4790),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__9284),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__13071),
            .DIN(N__13070),
            .DOUT(N__13069),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__13071),
            .PADOUT(N__13070),
            .PADIN(N__13069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9764),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__4835),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__13062),
            .DIN(N__13061),
            .DOUT(N__13060),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__13062),
            .PADOUT(N__13061),
            .PADIN(N__13060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4157),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__8222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__13053),
            .DIN(N__13052),
            .DOUT(N__13051),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__13053),
            .PADOUT(N__13052),
            .PADIN(N__13051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4958),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__8261),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__13044),
            .DIN(N__13043),
            .DOUT(N__13042),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__13044),
            .PADOUT(N__13043),
            .PADIN(N__13042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4253),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__7928),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__13035),
            .DIN(N__13034),
            .DOUT(N__13033),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__13035),
            .PADOUT(N__13034),
            .PADIN(N__13033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9878),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__8579),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__13026),
            .DIN(N__13025),
            .DOUT(N__13024),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__13026),
            .PADOUT(N__13025),
            .PADIN(N__13024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9667),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__13017),
            .DIN(N__13016),
            .DOUT(N__13015),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__13017),
            .PADOUT(N__13016),
            .PADIN(N__13015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9779),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__5894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__13008),
            .DIN(N__13007),
            .DOUT(N__13006),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__13008),
            .PADOUT(N__13007),
            .PADIN(N__13006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__12999),
            .DIN(N__12998),
            .DOUT(N__12997),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__12999),
            .PADOUT(N__12998),
            .PADIN(N__12997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4433),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__8096),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__12990),
            .DIN(N__12989),
            .DOUT(N__12988),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__12990),
            .PADOUT(N__12989),
            .PADIN(N__12988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4223),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__8318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12981),
            .DIN(N__12980),
            .DOUT(N__12979),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12981),
            .PADOUT(N__12980),
            .PADIN(N__12979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__12972),
            .DIN(N__12971),
            .DOUT(N__12970),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__12972),
            .PADOUT(N__12971),
            .PADIN(N__12970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10025),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__5126),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__12963),
            .DIN(N__12962),
            .DOUT(N__12961),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__12963),
            .PADOUT(N__12962),
            .PADIN(N__12961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9992),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__7352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__12954),
            .DIN(N__12953),
            .DOUT(N__12952),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__12954),
            .PADOUT(N__12953),
            .PADIN(N__12952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12755),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__7658),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__12945),
            .DIN(N__12944),
            .DOUT(N__12943),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__12945),
            .PADOUT(N__12944),
            .PADIN(N__12943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4418),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__5699),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__12936),
            .DIN(N__12935),
            .DOUT(N__12934),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__12936),
            .PADOUT(N__12935),
            .PADIN(N__12934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9947),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__4718),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__12927),
            .DIN(N__12926),
            .DOUT(N__12925),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__12927),
            .PADOUT(N__12926),
            .PADIN(N__12925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4172),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__8155),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__12918),
            .DIN(N__12917),
            .DOUT(N__12916),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__12918),
            .PADOUT(N__12917),
            .PADIN(N__12916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12794),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__7733),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__12909),
            .DIN(N__12908),
            .DOUT(N__12907),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__12909),
            .PADOUT(N__12908),
            .PADIN(N__12907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__12900),
            .DIN(N__12899),
            .DOUT(N__12898),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__12900),
            .PADOUT(N__12899),
            .PADIN(N__12898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4307),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__9347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__12891),
            .DIN(N__12890),
            .DOUT(N__12889),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__12891),
            .PADOUT(N__12890),
            .PADIN(N__12889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9698),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__5624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__12882),
            .DIN(N__12881),
            .DOUT(N__12880),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__12882),
            .PADOUT(N__12881),
            .PADIN(N__12880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4385),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__8174),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__12873),
            .DIN(N__12872),
            .DOUT(N__12871),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__12873),
            .PADOUT(N__12872),
            .PADIN(N__12871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4775),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__12864),
            .DIN(N__12863),
            .DOUT(N__12862),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__12864),
            .PADOUT(N__12863),
            .PADIN(N__12862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10136),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__7583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__12855),
            .DIN(N__12854),
            .DOUT(N__12853),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__12855),
            .PADOUT(N__12854),
            .PADIN(N__12853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5375),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__9365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__12846),
            .DIN(N__12845),
            .DOUT(N__12844),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__12846),
            .PADOUT(N__12845),
            .PADIN(N__12844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9842),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__5543),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__12837),
            .DIN(N__12836),
            .DOUT(N__12835),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__12837),
            .PADOUT(N__12836),
            .PADIN(N__12835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4112),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__8723),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__12828),
            .DIN(N__12827),
            .DOUT(N__12826),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__12828),
            .PADOUT(N__12827),
            .PADIN(N__12826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9614),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__8510),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__12819),
            .DIN(N__12818),
            .DOUT(N__12817),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__12819),
            .PADOUT(N__12818),
            .PADIN(N__12817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5330),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__8012),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3259 (
            .O(N__12800),
            .I(N__12797));
    LocalMux I__3258 (
            .O(N__12797),
            .I(READ_CYCLE_ACTIVE_rep3_i_ess));
    IoInMux I__3257 (
            .O(N__12794),
            .I(N__12791));
    LocalMux I__3256 (
            .O(N__12791),
            .I(N__12788));
    Span12Mux_s6_v I__3255 (
            .O(N__12788),
            .I(N__12785));
    Odrv12 I__3254 (
            .O(N__12785),
            .I(N_183_i));
    InMux I__3253 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__3252 (
            .O(N__12779),
            .I(READ_CYCLE_ACTIVE_rep9_i_ess));
    IoInMux I__3251 (
            .O(N__12776),
            .I(N__12773));
    LocalMux I__3250 (
            .O(N__12773),
            .I(N__12770));
    Span4Mux_s3_h I__3249 (
            .O(N__12770),
            .I(N__12767));
    Span4Mux_v I__3248 (
            .O(N__12767),
            .I(N__12764));
    Odrv4 I__3247 (
            .O(N__12764),
            .I(N_189_i));
    InMux I__3246 (
            .O(N__12761),
            .I(N__12758));
    LocalMux I__3245 (
            .O(N__12758),
            .I(READ_CYCLE_ACTIVE_rep11_i_ess));
    IoInMux I__3244 (
            .O(N__12755),
            .I(N__12752));
    LocalMux I__3243 (
            .O(N__12752),
            .I(N__12749));
    Span4Mux_s3_h I__3242 (
            .O(N__12749),
            .I(N__12746));
    Span4Mux_v I__3241 (
            .O(N__12746),
            .I(N__12743));
    Odrv4 I__3240 (
            .O(N__12743),
            .I(N_191_i));
    InMux I__3239 (
            .O(N__12740),
            .I(N__12737));
    LocalMux I__3238 (
            .O(N__12737),
            .I(READ_CYCLE_ACTIVE_rep15_i_ess));
    IoInMux I__3237 (
            .O(N__12734),
            .I(N__12731));
    LocalMux I__3236 (
            .O(N__12731),
            .I(N__12728));
    Span12Mux_s4_h I__3235 (
            .O(N__12728),
            .I(N__12725));
    Odrv12 I__3234 (
            .O(N__12725),
            .I(N_195_i));
    CascadeMux I__3233 (
            .O(N__12722),
            .I(N__12714));
    CascadeMux I__3232 (
            .O(N__12721),
            .I(N__12710));
    CascadeMux I__3231 (
            .O(N__12720),
            .I(N__12706));
    CascadeMux I__3230 (
            .O(N__12719),
            .I(N__12701));
    IoInMux I__3229 (
            .O(N__12718),
            .I(N__12696));
    InMux I__3228 (
            .O(N__12717),
            .I(N__12690));
    InMux I__3227 (
            .O(N__12714),
            .I(N__12686));
    InMux I__3226 (
            .O(N__12713),
            .I(N__12683));
    InMux I__3225 (
            .O(N__12710),
            .I(N__12680));
    CascadeMux I__3224 (
            .O(N__12709),
            .I(N__12674));
    InMux I__3223 (
            .O(N__12706),
            .I(N__12671));
    InMux I__3222 (
            .O(N__12705),
            .I(N__12666));
    CascadeMux I__3221 (
            .O(N__12704),
            .I(N__12663));
    InMux I__3220 (
            .O(N__12701),
            .I(N__12660));
    InMux I__3219 (
            .O(N__12700),
            .I(N__12655));
    InMux I__3218 (
            .O(N__12699),
            .I(N__12655));
    LocalMux I__3217 (
            .O(N__12696),
            .I(N__12652));
    CascadeMux I__3216 (
            .O(N__12695),
            .I(N__12649));
    CascadeMux I__3215 (
            .O(N__12694),
            .I(N__12646));
    CascadeMux I__3214 (
            .O(N__12693),
            .I(N__12643));
    LocalMux I__3213 (
            .O(N__12690),
            .I(N__12637));
    InMux I__3212 (
            .O(N__12689),
            .I(N__12634));
    LocalMux I__3211 (
            .O(N__12686),
            .I(N__12627));
    LocalMux I__3210 (
            .O(N__12683),
            .I(N__12627));
    LocalMux I__3209 (
            .O(N__12680),
            .I(N__12627));
    InMux I__3208 (
            .O(N__12679),
            .I(N__12624));
    InMux I__3207 (
            .O(N__12678),
            .I(N__12621));
    CascadeMux I__3206 (
            .O(N__12677),
            .I(N__12617));
    InMux I__3205 (
            .O(N__12674),
            .I(N__12614));
    LocalMux I__3204 (
            .O(N__12671),
            .I(N__12611));
    InMux I__3203 (
            .O(N__12670),
            .I(N__12608));
    InMux I__3202 (
            .O(N__12669),
            .I(N__12605));
    LocalMux I__3201 (
            .O(N__12666),
            .I(N__12600));
    InMux I__3200 (
            .O(N__12663),
            .I(N__12597));
    LocalMux I__3199 (
            .O(N__12660),
            .I(N__12586));
    LocalMux I__3198 (
            .O(N__12655),
            .I(N__12586));
    Span4Mux_s3_v I__3197 (
            .O(N__12652),
            .I(N__12583));
    InMux I__3196 (
            .O(N__12649),
            .I(N__12580));
    InMux I__3195 (
            .O(N__12646),
            .I(N__12575));
    InMux I__3194 (
            .O(N__12643),
            .I(N__12575));
    InMux I__3193 (
            .O(N__12642),
            .I(N__12570));
    InMux I__3192 (
            .O(N__12641),
            .I(N__12570));
    InMux I__3191 (
            .O(N__12640),
            .I(N__12567));
    Span4Mux_h I__3190 (
            .O(N__12637),
            .I(N__12562));
    LocalMux I__3189 (
            .O(N__12634),
            .I(N__12562));
    Span4Mux_v I__3188 (
            .O(N__12627),
            .I(N__12557));
    LocalMux I__3187 (
            .O(N__12624),
            .I(N__12557));
    LocalMux I__3186 (
            .O(N__12621),
            .I(N__12554));
    InMux I__3185 (
            .O(N__12620),
            .I(N__12551));
    InMux I__3184 (
            .O(N__12617),
            .I(N__12548));
    LocalMux I__3183 (
            .O(N__12614),
            .I(N__12541));
    Span4Mux_h I__3182 (
            .O(N__12611),
            .I(N__12534));
    LocalMux I__3181 (
            .O(N__12608),
            .I(N__12534));
    LocalMux I__3180 (
            .O(N__12605),
            .I(N__12534));
    InMux I__3179 (
            .O(N__12604),
            .I(N__12529));
    InMux I__3178 (
            .O(N__12603),
            .I(N__12529));
    Span4Mux_h I__3177 (
            .O(N__12600),
            .I(N__12521));
    LocalMux I__3176 (
            .O(N__12597),
            .I(N__12521));
    InMux I__3175 (
            .O(N__12596),
            .I(N__12516));
    InMux I__3174 (
            .O(N__12595),
            .I(N__12516));
    InMux I__3173 (
            .O(N__12594),
            .I(N__12509));
    InMux I__3172 (
            .O(N__12593),
            .I(N__12509));
    InMux I__3171 (
            .O(N__12592),
            .I(N__12509));
    InMux I__3170 (
            .O(N__12591),
            .I(N__12506));
    Span4Mux_v I__3169 (
            .O(N__12586),
            .I(N__12498));
    Span4Mux_v I__3168 (
            .O(N__12583),
            .I(N__12487));
    LocalMux I__3167 (
            .O(N__12580),
            .I(N__12487));
    LocalMux I__3166 (
            .O(N__12575),
            .I(N__12487));
    LocalMux I__3165 (
            .O(N__12570),
            .I(N__12487));
    LocalMux I__3164 (
            .O(N__12567),
            .I(N__12487));
    Span4Mux_v I__3163 (
            .O(N__12562),
            .I(N__12476));
    Span4Mux_v I__3162 (
            .O(N__12557),
            .I(N__12476));
    Span4Mux_v I__3161 (
            .O(N__12554),
            .I(N__12476));
    LocalMux I__3160 (
            .O(N__12551),
            .I(N__12476));
    LocalMux I__3159 (
            .O(N__12548),
            .I(N__12476));
    InMux I__3158 (
            .O(N__12547),
            .I(N__12469));
    InMux I__3157 (
            .O(N__12546),
            .I(N__12469));
    InMux I__3156 (
            .O(N__12545),
            .I(N__12469));
    CascadeMux I__3155 (
            .O(N__12544),
            .I(N__12464));
    Span4Mux_v I__3154 (
            .O(N__12541),
            .I(N__12459));
    Span4Mux_v I__3153 (
            .O(N__12534),
            .I(N__12459));
    LocalMux I__3152 (
            .O(N__12529),
            .I(N__12456));
    InMux I__3151 (
            .O(N__12528),
            .I(N__12453));
    InMux I__3150 (
            .O(N__12527),
            .I(N__12449));
    InMux I__3149 (
            .O(N__12526),
            .I(N__12446));
    Span4Mux_h I__3148 (
            .O(N__12521),
            .I(N__12434));
    LocalMux I__3147 (
            .O(N__12516),
            .I(N__12434));
    LocalMux I__3146 (
            .O(N__12509),
            .I(N__12434));
    LocalMux I__3145 (
            .O(N__12506),
            .I(N__12434));
    InMux I__3144 (
            .O(N__12505),
            .I(N__12431));
    CascadeMux I__3143 (
            .O(N__12504),
            .I(N__12427));
    CascadeMux I__3142 (
            .O(N__12503),
            .I(N__12423));
    CascadeMux I__3141 (
            .O(N__12502),
            .I(N__12420));
    CascadeMux I__3140 (
            .O(N__12501),
            .I(N__12416));
    Span4Mux_v I__3139 (
            .O(N__12498),
            .I(N__12407));
    Span4Mux_v I__3138 (
            .O(N__12487),
            .I(N__12402));
    Span4Mux_v I__3137 (
            .O(N__12476),
            .I(N__12402));
    LocalMux I__3136 (
            .O(N__12469),
            .I(N__12399));
    InMux I__3135 (
            .O(N__12468),
            .I(N__12392));
    InMux I__3134 (
            .O(N__12467),
            .I(N__12392));
    InMux I__3133 (
            .O(N__12464),
            .I(N__12392));
    Span4Mux_h I__3132 (
            .O(N__12459),
            .I(N__12385));
    Span4Mux_h I__3131 (
            .O(N__12456),
            .I(N__12385));
    LocalMux I__3130 (
            .O(N__12453),
            .I(N__12385));
    InMux I__3129 (
            .O(N__12452),
            .I(N__12382));
    LocalMux I__3128 (
            .O(N__12449),
            .I(N__12379));
    LocalMux I__3127 (
            .O(N__12446),
            .I(N__12376));
    InMux I__3126 (
            .O(N__12445),
            .I(N__12371));
    InMux I__3125 (
            .O(N__12444),
            .I(N__12371));
    InMux I__3124 (
            .O(N__12443),
            .I(N__12368));
    Span4Mux_v I__3123 (
            .O(N__12434),
            .I(N__12365));
    LocalMux I__3122 (
            .O(N__12431),
            .I(N__12362));
    InMux I__3121 (
            .O(N__12430),
            .I(N__12359));
    InMux I__3120 (
            .O(N__12427),
            .I(N__12356));
    InMux I__3119 (
            .O(N__12426),
            .I(N__12345));
    InMux I__3118 (
            .O(N__12423),
            .I(N__12345));
    InMux I__3117 (
            .O(N__12420),
            .I(N__12345));
    InMux I__3116 (
            .O(N__12419),
            .I(N__12345));
    InMux I__3115 (
            .O(N__12416),
            .I(N__12345));
    InMux I__3114 (
            .O(N__12415),
            .I(N__12342));
    InMux I__3113 (
            .O(N__12414),
            .I(N__12339));
    CascadeMux I__3112 (
            .O(N__12413),
            .I(N__12331));
    CascadeMux I__3111 (
            .O(N__12412),
            .I(N__12328));
    CascadeMux I__3110 (
            .O(N__12411),
            .I(N__12324));
    CascadeMux I__3109 (
            .O(N__12410),
            .I(N__12321));
    Sp12to4 I__3108 (
            .O(N__12407),
            .I(N__12316));
    Sp12to4 I__3107 (
            .O(N__12402),
            .I(N__12316));
    Span12Mux_s11_h I__3106 (
            .O(N__12399),
            .I(N__12313));
    LocalMux I__3105 (
            .O(N__12392),
            .I(N__12310));
    Sp12to4 I__3104 (
            .O(N__12385),
            .I(N__12305));
    LocalMux I__3103 (
            .O(N__12382),
            .I(N__12305));
    Span4Mux_v I__3102 (
            .O(N__12379),
            .I(N__12302));
    Span4Mux_h I__3101 (
            .O(N__12376),
            .I(N__12295));
    LocalMux I__3100 (
            .O(N__12371),
            .I(N__12295));
    LocalMux I__3099 (
            .O(N__12368),
            .I(N__12295));
    Span4Mux_v I__3098 (
            .O(N__12365),
            .I(N__12292));
    Span4Mux_h I__3097 (
            .O(N__12362),
            .I(N__12285));
    LocalMux I__3096 (
            .O(N__12359),
            .I(N__12285));
    LocalMux I__3095 (
            .O(N__12356),
            .I(N__12285));
    LocalMux I__3094 (
            .O(N__12345),
            .I(N__12280));
    LocalMux I__3093 (
            .O(N__12342),
            .I(N__12280));
    LocalMux I__3092 (
            .O(N__12339),
            .I(N__12277));
    InMux I__3091 (
            .O(N__12338),
            .I(N__12270));
    InMux I__3090 (
            .O(N__12337),
            .I(N__12270));
    InMux I__3089 (
            .O(N__12336),
            .I(N__12270));
    InMux I__3088 (
            .O(N__12335),
            .I(N__12263));
    InMux I__3087 (
            .O(N__12334),
            .I(N__12263));
    InMux I__3086 (
            .O(N__12331),
            .I(N__12263));
    InMux I__3085 (
            .O(N__12328),
            .I(N__12254));
    InMux I__3084 (
            .O(N__12327),
            .I(N__12254));
    InMux I__3083 (
            .O(N__12324),
            .I(N__12254));
    InMux I__3082 (
            .O(N__12321),
            .I(N__12254));
    Span12Mux_h I__3081 (
            .O(N__12316),
            .I(N__12251));
    Span12Mux_h I__3080 (
            .O(N__12313),
            .I(N__12248));
    Span12Mux_s11_h I__3079 (
            .O(N__12310),
            .I(N__12241));
    Span12Mux_s11_v I__3078 (
            .O(N__12305),
            .I(N__12241));
    Sp12to4 I__3077 (
            .O(N__12302),
            .I(N__12241));
    Span4Mux_v I__3076 (
            .O(N__12295),
            .I(N__12238));
    Span4Mux_v I__3075 (
            .O(N__12292),
            .I(N__12233));
    Span4Mux_v I__3074 (
            .O(N__12285),
            .I(N__12233));
    Span4Mux_v I__3073 (
            .O(N__12280),
            .I(N__12228));
    Span4Mux_v I__3072 (
            .O(N__12277),
            .I(N__12228));
    LocalMux I__3071 (
            .O(N__12270),
            .I(N__12225));
    LocalMux I__3070 (
            .O(N__12263),
            .I(N__12222));
    LocalMux I__3069 (
            .O(N__12254),
            .I(N__12219));
    Span12Mux_h I__3068 (
            .O(N__12251),
            .I(N__12216));
    Span12Mux_v I__3067 (
            .O(N__12248),
            .I(N__12211));
    Span12Mux_h I__3066 (
            .O(N__12241),
            .I(N__12211));
    Span4Mux_h I__3065 (
            .O(N__12238),
            .I(N__12208));
    Span4Mux_h I__3064 (
            .O(N__12233),
            .I(N__12205));
    Span4Mux_v I__3063 (
            .O(N__12228),
            .I(N__12196));
    Span4Mux_v I__3062 (
            .O(N__12225),
            .I(N__12196));
    Span4Mux_v I__3061 (
            .O(N__12222),
            .I(N__12196));
    Span4Mux_v I__3060 (
            .O(N__12219),
            .I(N__12196));
    Odrv12 I__3059 (
            .O(N__12216),
            .I(RnW_c));
    Odrv12 I__3058 (
            .O(N__12211),
            .I(RnW_c));
    Odrv4 I__3057 (
            .O(N__12208),
            .I(RnW_c));
    Odrv4 I__3056 (
            .O(N__12205),
            .I(RnW_c));
    Odrv4 I__3055 (
            .O(N__12196),
            .I(RnW_c));
    CascadeMux I__3054 (
            .O(N__12185),
            .I(N__12180));
    CascadeMux I__3053 (
            .O(N__12184),
            .I(N__12177));
    InMux I__3052 (
            .O(N__12183),
            .I(N__12172));
    InMux I__3051 (
            .O(N__12180),
            .I(N__12172));
    InMux I__3050 (
            .O(N__12177),
            .I(N__12169));
    LocalMux I__3049 (
            .O(N__12172),
            .I(N__12157));
    LocalMux I__3048 (
            .O(N__12169),
            .I(N__12157));
    InMux I__3047 (
            .O(N__12168),
            .I(N__12154));
    InMux I__3046 (
            .O(N__12167),
            .I(N__12151));
    InMux I__3045 (
            .O(N__12166),
            .I(N__12148));
    InMux I__3044 (
            .O(N__12165),
            .I(N__12145));
    CascadeMux I__3043 (
            .O(N__12164),
            .I(N__12141));
    CascadeMux I__3042 (
            .O(N__12163),
            .I(N__12138));
    CascadeMux I__3041 (
            .O(N__12162),
            .I(N__12128));
    Span4Mux_h I__3040 (
            .O(N__12157),
            .I(N__12119));
    LocalMux I__3039 (
            .O(N__12154),
            .I(N__12119));
    LocalMux I__3038 (
            .O(N__12151),
            .I(N__12119));
    LocalMux I__3037 (
            .O(N__12148),
            .I(N__12119));
    LocalMux I__3036 (
            .O(N__12145),
            .I(N__12116));
    InMux I__3035 (
            .O(N__12144),
            .I(N__12113));
    InMux I__3034 (
            .O(N__12141),
            .I(N__12110));
    InMux I__3033 (
            .O(N__12138),
            .I(N__12107));
    InMux I__3032 (
            .O(N__12137),
            .I(N__12103));
    CascadeMux I__3031 (
            .O(N__12136),
            .I(N__12100));
    InMux I__3030 (
            .O(N__12135),
            .I(N__12089));
    InMux I__3029 (
            .O(N__12134),
            .I(N__12089));
    InMux I__3028 (
            .O(N__12133),
            .I(N__12085));
    InMux I__3027 (
            .O(N__12132),
            .I(N__12082));
    InMux I__3026 (
            .O(N__12131),
            .I(N__12077));
    InMux I__3025 (
            .O(N__12128),
            .I(N__12077));
    Span4Mux_v I__3024 (
            .O(N__12119),
            .I(N__12058));
    Span4Mux_h I__3023 (
            .O(N__12116),
            .I(N__12058));
    LocalMux I__3022 (
            .O(N__12113),
            .I(N__12058));
    LocalMux I__3021 (
            .O(N__12110),
            .I(N__12058));
    LocalMux I__3020 (
            .O(N__12107),
            .I(N__12058));
    InMux I__3019 (
            .O(N__12106),
            .I(N__12055));
    LocalMux I__3018 (
            .O(N__12103),
            .I(N__12052));
    InMux I__3017 (
            .O(N__12100),
            .I(N__12049));
    InMux I__3016 (
            .O(N__12099),
            .I(N__12046));
    InMux I__3015 (
            .O(N__12098),
            .I(N__12039));
    InMux I__3014 (
            .O(N__12097),
            .I(N__12039));
    InMux I__3013 (
            .O(N__12096),
            .I(N__12039));
    CascadeMux I__3012 (
            .O(N__12095),
            .I(N__12036));
    CascadeMux I__3011 (
            .O(N__12094),
            .I(N__12026));
    LocalMux I__3010 (
            .O(N__12089),
            .I(N__12023));
    InMux I__3009 (
            .O(N__12088),
            .I(N__12020));
    LocalMux I__3008 (
            .O(N__12085),
            .I(N__12012));
    LocalMux I__3007 (
            .O(N__12082),
            .I(N__12012));
    LocalMux I__3006 (
            .O(N__12077),
            .I(N__12012));
    InMux I__3005 (
            .O(N__12076),
            .I(N__12009));
    InMux I__3004 (
            .O(N__12075),
            .I(N__11998));
    InMux I__3003 (
            .O(N__12074),
            .I(N__11998));
    InMux I__3002 (
            .O(N__12073),
            .I(N__11998));
    InMux I__3001 (
            .O(N__12072),
            .I(N__11998));
    InMux I__3000 (
            .O(N__12071),
            .I(N__11998));
    CascadeMux I__2999 (
            .O(N__12070),
            .I(N__11995));
    CascadeMux I__2998 (
            .O(N__12069),
            .I(N__11992));
    Span4Mux_v I__2997 (
            .O(N__12058),
            .I(N__11983));
    LocalMux I__2996 (
            .O(N__12055),
            .I(N__11983));
    Span4Mux_h I__2995 (
            .O(N__12052),
            .I(N__11976));
    LocalMux I__2994 (
            .O(N__12049),
            .I(N__11976));
    LocalMux I__2993 (
            .O(N__12046),
            .I(N__11976));
    LocalMux I__2992 (
            .O(N__12039),
            .I(N__11973));
    InMux I__2991 (
            .O(N__12036),
            .I(N__11970));
    InMux I__2990 (
            .O(N__12035),
            .I(N__11965));
    InMux I__2989 (
            .O(N__12034),
            .I(N__11965));
    InMux I__2988 (
            .O(N__12033),
            .I(N__11962));
    InMux I__2987 (
            .O(N__12032),
            .I(N__11959));
    CascadeMux I__2986 (
            .O(N__12031),
            .I(N__11954));
    CascadeMux I__2985 (
            .O(N__12030),
            .I(N__11949));
    CascadeMux I__2984 (
            .O(N__12029),
            .I(N__11946));
    InMux I__2983 (
            .O(N__12026),
            .I(N__11939));
    Span4Mux_h I__2982 (
            .O(N__12023),
            .I(N__11936));
    LocalMux I__2981 (
            .O(N__12020),
            .I(N__11933));
    CascadeMux I__2980 (
            .O(N__12019),
            .I(N__11929));
    Span4Mux_v I__2979 (
            .O(N__12012),
            .I(N__11924));
    LocalMux I__2978 (
            .O(N__12009),
            .I(N__11924));
    LocalMux I__2977 (
            .O(N__11998),
            .I(N__11921));
    InMux I__2976 (
            .O(N__11995),
            .I(N__11918));
    InMux I__2975 (
            .O(N__11992),
            .I(N__11915));
    CascadeMux I__2974 (
            .O(N__11991),
            .I(N__11909));
    CascadeMux I__2973 (
            .O(N__11990),
            .I(N__11906));
    CascadeMux I__2972 (
            .O(N__11989),
            .I(N__11902));
    CascadeMux I__2971 (
            .O(N__11988),
            .I(N__11899));
    Span4Mux_v I__2970 (
            .O(N__11983),
            .I(N__11884));
    Span4Mux_v I__2969 (
            .O(N__11976),
            .I(N__11884));
    Span4Mux_h I__2968 (
            .O(N__11973),
            .I(N__11884));
    LocalMux I__2967 (
            .O(N__11970),
            .I(N__11884));
    LocalMux I__2966 (
            .O(N__11965),
            .I(N__11884));
    LocalMux I__2965 (
            .O(N__11962),
            .I(N__11884));
    LocalMux I__2964 (
            .O(N__11959),
            .I(N__11884));
    InMux I__2963 (
            .O(N__11958),
            .I(N__11879));
    InMux I__2962 (
            .O(N__11957),
            .I(N__11879));
    InMux I__2961 (
            .O(N__11954),
            .I(N__11876));
    InMux I__2960 (
            .O(N__11953),
            .I(N__11872));
    InMux I__2959 (
            .O(N__11952),
            .I(N__11865));
    InMux I__2958 (
            .O(N__11949),
            .I(N__11865));
    InMux I__2957 (
            .O(N__11946),
            .I(N__11865));
    InMux I__2956 (
            .O(N__11945),
            .I(N__11862));
    CascadeMux I__2955 (
            .O(N__11944),
            .I(N__11859));
    CascadeMux I__2954 (
            .O(N__11943),
            .I(N__11856));
    CascadeMux I__2953 (
            .O(N__11942),
            .I(N__11853));
    LocalMux I__2952 (
            .O(N__11939),
            .I(N__11850));
    Span4Mux_v I__2951 (
            .O(N__11936),
            .I(N__11845));
    Span4Mux_h I__2950 (
            .O(N__11933),
            .I(N__11845));
    CascadeMux I__2949 (
            .O(N__11932),
            .I(N__11842));
    InMux I__2948 (
            .O(N__11929),
            .I(N__11839));
    Span4Mux_v I__2947 (
            .O(N__11924),
            .I(N__11830));
    Span4Mux_v I__2946 (
            .O(N__11921),
            .I(N__11830));
    LocalMux I__2945 (
            .O(N__11918),
            .I(N__11830));
    LocalMux I__2944 (
            .O(N__11915),
            .I(N__11830));
    CascadeMux I__2943 (
            .O(N__11914),
            .I(N__11826));
    CascadeMux I__2942 (
            .O(N__11913),
            .I(N__11821));
    CascadeMux I__2941 (
            .O(N__11912),
            .I(N__11818));
    InMux I__2940 (
            .O(N__11909),
            .I(N__11811));
    InMux I__2939 (
            .O(N__11906),
            .I(N__11811));
    InMux I__2938 (
            .O(N__11905),
            .I(N__11804));
    InMux I__2937 (
            .O(N__11902),
            .I(N__11804));
    InMux I__2936 (
            .O(N__11899),
            .I(N__11804));
    Span4Mux_v I__2935 (
            .O(N__11884),
            .I(N__11799));
    LocalMux I__2934 (
            .O(N__11879),
            .I(N__11799));
    LocalMux I__2933 (
            .O(N__11876),
            .I(N__11796));
    InMux I__2932 (
            .O(N__11875),
            .I(N__11793));
    LocalMux I__2931 (
            .O(N__11872),
            .I(N__11790));
    LocalMux I__2930 (
            .O(N__11865),
            .I(N__11785));
    LocalMux I__2929 (
            .O(N__11862),
            .I(N__11785));
    InMux I__2928 (
            .O(N__11859),
            .I(N__11780));
    InMux I__2927 (
            .O(N__11856),
            .I(N__11780));
    InMux I__2926 (
            .O(N__11853),
            .I(N__11777));
    Span4Mux_h I__2925 (
            .O(N__11850),
            .I(N__11772));
    Span4Mux_v I__2924 (
            .O(N__11845),
            .I(N__11772));
    InMux I__2923 (
            .O(N__11842),
            .I(N__11769));
    LocalMux I__2922 (
            .O(N__11839),
            .I(N__11766));
    Span4Mux_v I__2921 (
            .O(N__11830),
            .I(N__11763));
    InMux I__2920 (
            .O(N__11829),
            .I(N__11754));
    InMux I__2919 (
            .O(N__11826),
            .I(N__11754));
    InMux I__2918 (
            .O(N__11825),
            .I(N__11754));
    InMux I__2917 (
            .O(N__11824),
            .I(N__11754));
    InMux I__2916 (
            .O(N__11821),
            .I(N__11747));
    InMux I__2915 (
            .O(N__11818),
            .I(N__11747));
    InMux I__2914 (
            .O(N__11817),
            .I(N__11747));
    CascadeMux I__2913 (
            .O(N__11816),
            .I(N__11743));
    LocalMux I__2912 (
            .O(N__11811),
            .I(N__11737));
    LocalMux I__2911 (
            .O(N__11804),
            .I(N__11737));
    Span4Mux_h I__2910 (
            .O(N__11799),
            .I(N__11730));
    Span4Mux_v I__2909 (
            .O(N__11796),
            .I(N__11730));
    LocalMux I__2908 (
            .O(N__11793),
            .I(N__11730));
    Span4Mux_v I__2907 (
            .O(N__11790),
            .I(N__11721));
    Span4Mux_h I__2906 (
            .O(N__11785),
            .I(N__11721));
    LocalMux I__2905 (
            .O(N__11780),
            .I(N__11721));
    LocalMux I__2904 (
            .O(N__11777),
            .I(N__11721));
    Span4Mux_h I__2903 (
            .O(N__11772),
            .I(N__11716));
    LocalMux I__2902 (
            .O(N__11769),
            .I(N__11716));
    Span12Mux_h I__2901 (
            .O(N__11766),
            .I(N__11709));
    Sp12to4 I__2900 (
            .O(N__11763),
            .I(N__11709));
    LocalMux I__2899 (
            .O(N__11754),
            .I(N__11709));
    LocalMux I__2898 (
            .O(N__11747),
            .I(N__11706));
    InMux I__2897 (
            .O(N__11746),
            .I(N__11703));
    InMux I__2896 (
            .O(N__11743),
            .I(N__11698));
    InMux I__2895 (
            .O(N__11742),
            .I(N__11698));
    Span4Mux_v I__2894 (
            .O(N__11737),
            .I(N__11695));
    Span4Mux_h I__2893 (
            .O(N__11730),
            .I(N__11692));
    Span4Mux_h I__2892 (
            .O(N__11721),
            .I(N__11689));
    Span4Mux_v I__2891 (
            .O(N__11716),
            .I(N__11686));
    Span12Mux_h I__2890 (
            .O(N__11709),
            .I(N__11683));
    Span12Mux_h I__2889 (
            .O(N__11706),
            .I(N__11680));
    LocalMux I__2888 (
            .O(N__11703),
            .I(N__11675));
    LocalMux I__2887 (
            .O(N__11698),
            .I(N__11675));
    Sp12to4 I__2886 (
            .O(N__11695),
            .I(N__11672));
    Span4Mux_v I__2885 (
            .O(N__11692),
            .I(N__11669));
    Span4Mux_v I__2884 (
            .O(N__11689),
            .I(N__11666));
    Span4Mux_v I__2883 (
            .O(N__11686),
            .I(N__11663));
    Span12Mux_v I__2882 (
            .O(N__11683),
            .I(N__11660));
    Span12Mux_v I__2881 (
            .O(N__11680),
            .I(N__11655));
    Span12Mux_h I__2880 (
            .O(N__11675),
            .I(N__11655));
    Span12Mux_h I__2879 (
            .O(N__11672),
            .I(N__11652));
    Span4Mux_h I__2878 (
            .O(N__11669),
            .I(N__11647));
    Span4Mux_h I__2877 (
            .O(N__11666),
            .I(N__11647));
    IoSpan4Mux I__2876 (
            .O(N__11663),
            .I(N__11644));
    Odrv12 I__2875 (
            .O(N__11660),
            .I(TS_CPUn_c));
    Odrv12 I__2874 (
            .O(N__11655),
            .I(TS_CPUn_c));
    Odrv12 I__2873 (
            .O(N__11652),
            .I(TS_CPUn_c));
    Odrv4 I__2872 (
            .O(N__11647),
            .I(TS_CPUn_c));
    Odrv4 I__2871 (
            .O(N__11644),
            .I(TS_CPUn_c));
    InMux I__2870 (
            .O(N__11633),
            .I(N__11626));
    InMux I__2869 (
            .O(N__11632),
            .I(N__11621));
    InMux I__2868 (
            .O(N__11631),
            .I(N__11621));
    CascadeMux I__2867 (
            .O(N__11630),
            .I(N__11612));
    CascadeMux I__2866 (
            .O(N__11629),
            .I(N__11609));
    LocalMux I__2865 (
            .O(N__11626),
            .I(N__11601));
    LocalMux I__2864 (
            .O(N__11621),
            .I(N__11601));
    InMux I__2863 (
            .O(N__11620),
            .I(N__11596));
    InMux I__2862 (
            .O(N__11619),
            .I(N__11596));
    CascadeMux I__2861 (
            .O(N__11618),
            .I(N__11593));
    InMux I__2860 (
            .O(N__11617),
            .I(N__11590));
    InMux I__2859 (
            .O(N__11616),
            .I(N__11585));
    InMux I__2858 (
            .O(N__11615),
            .I(N__11585));
    InMux I__2857 (
            .O(N__11612),
            .I(N__11580));
    InMux I__2856 (
            .O(N__11609),
            .I(N__11580));
    InMux I__2855 (
            .O(N__11608),
            .I(N__11577));
    InMux I__2854 (
            .O(N__11607),
            .I(N__11574));
    CascadeMux I__2853 (
            .O(N__11606),
            .I(N__11567));
    Span4Mux_v I__2852 (
            .O(N__11601),
            .I(N__11558));
    LocalMux I__2851 (
            .O(N__11596),
            .I(N__11558));
    InMux I__2850 (
            .O(N__11593),
            .I(N__11555));
    LocalMux I__2849 (
            .O(N__11590),
            .I(N__11545));
    LocalMux I__2848 (
            .O(N__11585),
            .I(N__11536));
    LocalMux I__2847 (
            .O(N__11580),
            .I(N__11536));
    LocalMux I__2846 (
            .O(N__11577),
            .I(N__11536));
    LocalMux I__2845 (
            .O(N__11574),
            .I(N__11536));
    InMux I__2844 (
            .O(N__11573),
            .I(N__11529));
    InMux I__2843 (
            .O(N__11572),
            .I(N__11529));
    InMux I__2842 (
            .O(N__11571),
            .I(N__11529));
    InMux I__2841 (
            .O(N__11570),
            .I(N__11526));
    InMux I__2840 (
            .O(N__11567),
            .I(N__11523));
    InMux I__2839 (
            .O(N__11566),
            .I(N__11520));
    InMux I__2838 (
            .O(N__11565),
            .I(N__11517));
    CascadeMux I__2837 (
            .O(N__11564),
            .I(N__11511));
    InMux I__2836 (
            .O(N__11563),
            .I(N__11506));
    Span4Mux_h I__2835 (
            .O(N__11558),
            .I(N__11498));
    LocalMux I__2834 (
            .O(N__11555),
            .I(N__11498));
    InMux I__2833 (
            .O(N__11554),
            .I(N__11495));
    CascadeMux I__2832 (
            .O(N__11553),
            .I(N__11492));
    CascadeMux I__2831 (
            .O(N__11552),
            .I(N__11489));
    CascadeMux I__2830 (
            .O(N__11551),
            .I(N__11484));
    CascadeMux I__2829 (
            .O(N__11550),
            .I(N__11479));
    CascadeMux I__2828 (
            .O(N__11549),
            .I(N__11469));
    CascadeMux I__2827 (
            .O(N__11548),
            .I(N__11466));
    Span4Mux_v I__2826 (
            .O(N__11545),
            .I(N__11450));
    Span4Mux_v I__2825 (
            .O(N__11536),
            .I(N__11450));
    LocalMux I__2824 (
            .O(N__11529),
            .I(N__11450));
    LocalMux I__2823 (
            .O(N__11526),
            .I(N__11450));
    LocalMux I__2822 (
            .O(N__11523),
            .I(N__11450));
    LocalMux I__2821 (
            .O(N__11520),
            .I(N__11450));
    LocalMux I__2820 (
            .O(N__11517),
            .I(N__11450));
    InMux I__2819 (
            .O(N__11516),
            .I(N__11447));
    InMux I__2818 (
            .O(N__11515),
            .I(N__11444));
    InMux I__2817 (
            .O(N__11514),
            .I(N__11441));
    InMux I__2816 (
            .O(N__11511),
            .I(N__11438));
    CascadeMux I__2815 (
            .O(N__11510),
            .I(N__11435));
    CascadeMux I__2814 (
            .O(N__11509),
            .I(N__11431));
    LocalMux I__2813 (
            .O(N__11506),
            .I(N__11427));
    InMux I__2812 (
            .O(N__11505),
            .I(N__11424));
    InMux I__2811 (
            .O(N__11504),
            .I(N__11421));
    InMux I__2810 (
            .O(N__11503),
            .I(N__11418));
    Span4Mux_v I__2809 (
            .O(N__11498),
            .I(N__11415));
    LocalMux I__2808 (
            .O(N__11495),
            .I(N__11412));
    InMux I__2807 (
            .O(N__11492),
            .I(N__11409));
    InMux I__2806 (
            .O(N__11489),
            .I(N__11401));
    InMux I__2805 (
            .O(N__11488),
            .I(N__11401));
    InMux I__2804 (
            .O(N__11487),
            .I(N__11401));
    InMux I__2803 (
            .O(N__11484),
            .I(N__11398));
    InMux I__2802 (
            .O(N__11483),
            .I(N__11393));
    InMux I__2801 (
            .O(N__11482),
            .I(N__11393));
    InMux I__2800 (
            .O(N__11479),
            .I(N__11390));
    InMux I__2799 (
            .O(N__11478),
            .I(N__11385));
    InMux I__2798 (
            .O(N__11477),
            .I(N__11385));
    InMux I__2797 (
            .O(N__11476),
            .I(N__11382));
    InMux I__2796 (
            .O(N__11475),
            .I(N__11379));
    CascadeMux I__2795 (
            .O(N__11474),
            .I(N__11370));
    CascadeMux I__2794 (
            .O(N__11473),
            .I(N__11365));
    CascadeMux I__2793 (
            .O(N__11472),
            .I(N__11359));
    InMux I__2792 (
            .O(N__11469),
            .I(N__11355));
    InMux I__2791 (
            .O(N__11466),
            .I(N__11350));
    InMux I__2790 (
            .O(N__11465),
            .I(N__11350));
    Span4Mux_v I__2789 (
            .O(N__11450),
            .I(N__11338));
    LocalMux I__2788 (
            .O(N__11447),
            .I(N__11338));
    LocalMux I__2787 (
            .O(N__11444),
            .I(N__11338));
    LocalMux I__2786 (
            .O(N__11441),
            .I(N__11338));
    LocalMux I__2785 (
            .O(N__11438),
            .I(N__11338));
    InMux I__2784 (
            .O(N__11435),
            .I(N__11335));
    InMux I__2783 (
            .O(N__11434),
            .I(N__11332));
    InMux I__2782 (
            .O(N__11431),
            .I(N__11329));
    InMux I__2781 (
            .O(N__11430),
            .I(N__11326));
    Span4Mux_v I__2780 (
            .O(N__11427),
            .I(N__11321));
    LocalMux I__2779 (
            .O(N__11424),
            .I(N__11321));
    LocalMux I__2778 (
            .O(N__11421),
            .I(N__11316));
    LocalMux I__2777 (
            .O(N__11418),
            .I(N__11316));
    Span4Mux_h I__2776 (
            .O(N__11415),
            .I(N__11309));
    Span4Mux_v I__2775 (
            .O(N__11412),
            .I(N__11309));
    LocalMux I__2774 (
            .O(N__11409),
            .I(N__11309));
    CascadeMux I__2773 (
            .O(N__11408),
            .I(N__11305));
    LocalMux I__2772 (
            .O(N__11401),
            .I(N__11298));
    LocalMux I__2771 (
            .O(N__11398),
            .I(N__11298));
    LocalMux I__2770 (
            .O(N__11393),
            .I(N__11298));
    LocalMux I__2769 (
            .O(N__11390),
            .I(N__11289));
    LocalMux I__2768 (
            .O(N__11385),
            .I(N__11289));
    LocalMux I__2767 (
            .O(N__11382),
            .I(N__11289));
    LocalMux I__2766 (
            .O(N__11379),
            .I(N__11289));
    InMux I__2765 (
            .O(N__11378),
            .I(N__11280));
    InMux I__2764 (
            .O(N__11377),
            .I(N__11280));
    InMux I__2763 (
            .O(N__11376),
            .I(N__11280));
    InMux I__2762 (
            .O(N__11375),
            .I(N__11280));
    InMux I__2761 (
            .O(N__11374),
            .I(N__11275));
    InMux I__2760 (
            .O(N__11373),
            .I(N__11275));
    InMux I__2759 (
            .O(N__11370),
            .I(N__11264));
    InMux I__2758 (
            .O(N__11369),
            .I(N__11264));
    InMux I__2757 (
            .O(N__11368),
            .I(N__11264));
    InMux I__2756 (
            .O(N__11365),
            .I(N__11264));
    InMux I__2755 (
            .O(N__11364),
            .I(N__11264));
    InMux I__2754 (
            .O(N__11363),
            .I(N__11257));
    InMux I__2753 (
            .O(N__11362),
            .I(N__11257));
    InMux I__2752 (
            .O(N__11359),
            .I(N__11257));
    InMux I__2751 (
            .O(N__11358),
            .I(N__11254));
    LocalMux I__2750 (
            .O(N__11355),
            .I(N__11249));
    LocalMux I__2749 (
            .O(N__11350),
            .I(N__11249));
    CascadeMux I__2748 (
            .O(N__11349),
            .I(N__11246));
    Span4Mux_v I__2747 (
            .O(N__11338),
            .I(N__11241));
    LocalMux I__2746 (
            .O(N__11335),
            .I(N__11241));
    LocalMux I__2745 (
            .O(N__11332),
            .I(N__11234));
    LocalMux I__2744 (
            .O(N__11329),
            .I(N__11234));
    LocalMux I__2743 (
            .O(N__11326),
            .I(N__11234));
    Span4Mux_v I__2742 (
            .O(N__11321),
            .I(N__11228));
    Span4Mux_v I__2741 (
            .O(N__11316),
            .I(N__11225));
    Span4Mux_v I__2740 (
            .O(N__11309),
            .I(N__11222));
    InMux I__2739 (
            .O(N__11308),
            .I(N__11217));
    InMux I__2738 (
            .O(N__11305),
            .I(N__11217));
    Span12Mux_v I__2737 (
            .O(N__11298),
            .I(N__11213));
    Span12Mux_h I__2736 (
            .O(N__11289),
            .I(N__11210));
    LocalMux I__2735 (
            .O(N__11280),
            .I(N__11201));
    LocalMux I__2734 (
            .O(N__11275),
            .I(N__11201));
    LocalMux I__2733 (
            .O(N__11264),
            .I(N__11201));
    LocalMux I__2732 (
            .O(N__11257),
            .I(N__11201));
    LocalMux I__2731 (
            .O(N__11254),
            .I(N__11198));
    Span4Mux_v I__2730 (
            .O(N__11249),
            .I(N__11195));
    InMux I__2729 (
            .O(N__11246),
            .I(N__11192));
    Span4Mux_v I__2728 (
            .O(N__11241),
            .I(N__11187));
    Span4Mux_v I__2727 (
            .O(N__11234),
            .I(N__11187));
    InMux I__2726 (
            .O(N__11233),
            .I(N__11180));
    InMux I__2725 (
            .O(N__11232),
            .I(N__11180));
    InMux I__2724 (
            .O(N__11231),
            .I(N__11180));
    Span4Mux_h I__2723 (
            .O(N__11228),
            .I(N__11177));
    Sp12to4 I__2722 (
            .O(N__11225),
            .I(N__11172));
    Sp12to4 I__2721 (
            .O(N__11222),
            .I(N__11172));
    LocalMux I__2720 (
            .O(N__11217),
            .I(N__11169));
    InMux I__2719 (
            .O(N__11216),
            .I(N__11166));
    Span12Mux_h I__2718 (
            .O(N__11213),
            .I(N__11161));
    Span12Mux_v I__2717 (
            .O(N__11210),
            .I(N__11161));
    Span12Mux_v I__2716 (
            .O(N__11201),
            .I(N__11152));
    Span12Mux_s8_v I__2715 (
            .O(N__11198),
            .I(N__11152));
    Sp12to4 I__2714 (
            .O(N__11195),
            .I(N__11152));
    LocalMux I__2713 (
            .O(N__11192),
            .I(N__11152));
    Sp12to4 I__2712 (
            .O(N__11187),
            .I(N__11147));
    LocalMux I__2711 (
            .O(N__11180),
            .I(N__11147));
    Sp12to4 I__2710 (
            .O(N__11177),
            .I(N__11140));
    Span12Mux_h I__2709 (
            .O(N__11172),
            .I(N__11140));
    Sp12to4 I__2708 (
            .O(N__11169),
            .I(N__11140));
    LocalMux I__2707 (
            .O(N__11166),
            .I(N__11137));
    Span12Mux_v I__2706 (
            .O(N__11161),
            .I(N__11134));
    Span12Mux_h I__2705 (
            .O(N__11152),
            .I(N__11127));
    Span12Mux_h I__2704 (
            .O(N__11147),
            .I(N__11127));
    Span12Mux_v I__2703 (
            .O(N__11140),
            .I(N__11127));
    Span4Mux_v I__2702 (
            .O(N__11137),
            .I(N__11124));
    Odrv12 I__2701 (
            .O(N__11134),
            .I(LBENn_c));
    Odrv12 I__2700 (
            .O(N__11127),
            .I(LBENn_c));
    Odrv4 I__2699 (
            .O(N__11124),
            .I(LBENn_c));
    InMux I__2698 (
            .O(N__11117),
            .I(N__11103));
    InMux I__2697 (
            .O(N__11116),
            .I(N__11100));
    InMux I__2696 (
            .O(N__11115),
            .I(N__11097));
    InMux I__2695 (
            .O(N__11114),
            .I(N__11094));
    CascadeMux I__2694 (
            .O(N__11113),
            .I(N__11080));
    InMux I__2693 (
            .O(N__11112),
            .I(N__11076));
    InMux I__2692 (
            .O(N__11111),
            .I(N__11071));
    InMux I__2691 (
            .O(N__11110),
            .I(N__11071));
    InMux I__2690 (
            .O(N__11109),
            .I(N__11066));
    InMux I__2689 (
            .O(N__11108),
            .I(N__11066));
    CascadeMux I__2688 (
            .O(N__11107),
            .I(N__11061));
    CascadeMux I__2687 (
            .O(N__11106),
            .I(N__11058));
    LocalMux I__2686 (
            .O(N__11103),
            .I(N__11054));
    LocalMux I__2685 (
            .O(N__11100),
            .I(N__11049));
    LocalMux I__2684 (
            .O(N__11097),
            .I(N__11049));
    LocalMux I__2683 (
            .O(N__11094),
            .I(N__11046));
    InMux I__2682 (
            .O(N__11093),
            .I(N__11043));
    InMux I__2681 (
            .O(N__11092),
            .I(N__11040));
    InMux I__2680 (
            .O(N__11091),
            .I(N__11037));
    InMux I__2679 (
            .O(N__11090),
            .I(N__11034));
    InMux I__2678 (
            .O(N__11089),
            .I(N__11022));
    InMux I__2677 (
            .O(N__11088),
            .I(N__11022));
    InMux I__2676 (
            .O(N__11087),
            .I(N__11022));
    InMux I__2675 (
            .O(N__11086),
            .I(N__11017));
    InMux I__2674 (
            .O(N__11085),
            .I(N__11017));
    InMux I__2673 (
            .O(N__11084),
            .I(N__11008));
    InMux I__2672 (
            .O(N__11083),
            .I(N__11008));
    InMux I__2671 (
            .O(N__11080),
            .I(N__11003));
    InMux I__2670 (
            .O(N__11079),
            .I(N__11003));
    LocalMux I__2669 (
            .O(N__11076),
            .I(N__10996));
    LocalMux I__2668 (
            .O(N__11071),
            .I(N__10996));
    LocalMux I__2667 (
            .O(N__11066),
            .I(N__10993));
    InMux I__2666 (
            .O(N__11065),
            .I(N__10990));
    InMux I__2665 (
            .O(N__11064),
            .I(N__10987));
    InMux I__2664 (
            .O(N__11061),
            .I(N__10980));
    InMux I__2663 (
            .O(N__11058),
            .I(N__10980));
    InMux I__2662 (
            .O(N__11057),
            .I(N__10980));
    Span4Mux_v I__2661 (
            .O(N__11054),
            .I(N__10967));
    Span4Mux_v I__2660 (
            .O(N__11049),
            .I(N__10967));
    Span4Mux_h I__2659 (
            .O(N__11046),
            .I(N__10967));
    LocalMux I__2658 (
            .O(N__11043),
            .I(N__10967));
    LocalMux I__2657 (
            .O(N__11040),
            .I(N__10967));
    LocalMux I__2656 (
            .O(N__11037),
            .I(N__10967));
    LocalMux I__2655 (
            .O(N__11034),
            .I(N__10964));
    InMux I__2654 (
            .O(N__11033),
            .I(N__10961));
    InMux I__2653 (
            .O(N__11032),
            .I(N__10958));
    InMux I__2652 (
            .O(N__11031),
            .I(N__10955));
    InMux I__2651 (
            .O(N__11030),
            .I(N__10952));
    InMux I__2650 (
            .O(N__11029),
            .I(N__10949));
    LocalMux I__2649 (
            .O(N__11022),
            .I(N__10944));
    LocalMux I__2648 (
            .O(N__11017),
            .I(N__10944));
    InMux I__2647 (
            .O(N__11016),
            .I(N__10941));
    InMux I__2646 (
            .O(N__11015),
            .I(N__10938));
    InMux I__2645 (
            .O(N__11014),
            .I(N__10935));
    InMux I__2644 (
            .O(N__11013),
            .I(N__10932));
    LocalMux I__2643 (
            .O(N__11008),
            .I(N__10922));
    LocalMux I__2642 (
            .O(N__11003),
            .I(N__10919));
    InMux I__2641 (
            .O(N__11002),
            .I(N__10914));
    InMux I__2640 (
            .O(N__11001),
            .I(N__10914));
    Span4Mux_v I__2639 (
            .O(N__10996),
            .I(N__10903));
    Span4Mux_h I__2638 (
            .O(N__10993),
            .I(N__10903));
    LocalMux I__2637 (
            .O(N__10990),
            .I(N__10903));
    LocalMux I__2636 (
            .O(N__10987),
            .I(N__10903));
    LocalMux I__2635 (
            .O(N__10980),
            .I(N__10903));
    Span4Mux_v I__2634 (
            .O(N__10967),
            .I(N__10888));
    Span4Mux_h I__2633 (
            .O(N__10964),
            .I(N__10888));
    LocalMux I__2632 (
            .O(N__10961),
            .I(N__10888));
    LocalMux I__2631 (
            .O(N__10958),
            .I(N__10888));
    LocalMux I__2630 (
            .O(N__10955),
            .I(N__10888));
    LocalMux I__2629 (
            .O(N__10952),
            .I(N__10888));
    LocalMux I__2628 (
            .O(N__10949),
            .I(N__10888));
    Span4Mux_v I__2627 (
            .O(N__10944),
            .I(N__10883));
    LocalMux I__2626 (
            .O(N__10941),
            .I(N__10883));
    LocalMux I__2625 (
            .O(N__10938),
            .I(N__10880));
    LocalMux I__2624 (
            .O(N__10935),
            .I(N__10877));
    LocalMux I__2623 (
            .O(N__10932),
            .I(N__10874));
    InMux I__2622 (
            .O(N__10931),
            .I(N__10871));
    InMux I__2621 (
            .O(N__10930),
            .I(N__10868));
    InMux I__2620 (
            .O(N__10929),
            .I(N__10860));
    InMux I__2619 (
            .O(N__10928),
            .I(N__10853));
    InMux I__2618 (
            .O(N__10927),
            .I(N__10853));
    InMux I__2617 (
            .O(N__10926),
            .I(N__10853));
    InMux I__2616 (
            .O(N__10925),
            .I(N__10850));
    Span4Mux_h I__2615 (
            .O(N__10922),
            .I(N__10842));
    Span12Mux_v I__2614 (
            .O(N__10919),
            .I(N__10837));
    LocalMux I__2613 (
            .O(N__10914),
            .I(N__10834));
    Span4Mux_v I__2612 (
            .O(N__10903),
            .I(N__10829));
    Span4Mux_v I__2611 (
            .O(N__10888),
            .I(N__10829));
    Span4Mux_h I__2610 (
            .O(N__10883),
            .I(N__10824));
    Span4Mux_v I__2609 (
            .O(N__10880),
            .I(N__10824));
    Span4Mux_v I__2608 (
            .O(N__10877),
            .I(N__10818));
    Span4Mux_v I__2607 (
            .O(N__10874),
            .I(N__10815));
    LocalMux I__2606 (
            .O(N__10871),
            .I(N__10812));
    LocalMux I__2605 (
            .O(N__10868),
            .I(N__10809));
    InMux I__2604 (
            .O(N__10867),
            .I(N__10806));
    InMux I__2603 (
            .O(N__10866),
            .I(N__10803));
    InMux I__2602 (
            .O(N__10865),
            .I(N__10796));
    InMux I__2601 (
            .O(N__10864),
            .I(N__10796));
    InMux I__2600 (
            .O(N__10863),
            .I(N__10796));
    LocalMux I__2599 (
            .O(N__10860),
            .I(N__10788));
    LocalMux I__2598 (
            .O(N__10853),
            .I(N__10788));
    LocalMux I__2597 (
            .O(N__10850),
            .I(N__10785));
    InMux I__2596 (
            .O(N__10849),
            .I(N__10774));
    InMux I__2595 (
            .O(N__10848),
            .I(N__10774));
    InMux I__2594 (
            .O(N__10847),
            .I(N__10774));
    InMux I__2593 (
            .O(N__10846),
            .I(N__10774));
    InMux I__2592 (
            .O(N__10845),
            .I(N__10774));
    Span4Mux_h I__2591 (
            .O(N__10842),
            .I(N__10771));
    InMux I__2590 (
            .O(N__10841),
            .I(N__10766));
    InMux I__2589 (
            .O(N__10840),
            .I(N__10766));
    Span12Mux_h I__2588 (
            .O(N__10837),
            .I(N__10759));
    Span4Mux_h I__2587 (
            .O(N__10834),
            .I(N__10756));
    Sp12to4 I__2586 (
            .O(N__10829),
            .I(N__10753));
    Span4Mux_v I__2585 (
            .O(N__10824),
            .I(N__10750));
    InMux I__2584 (
            .O(N__10823),
            .I(N__10747));
    InMux I__2583 (
            .O(N__10822),
            .I(N__10742));
    InMux I__2582 (
            .O(N__10821),
            .I(N__10742));
    Span4Mux_v I__2581 (
            .O(N__10818),
            .I(N__10739));
    Span4Mux_h I__2580 (
            .O(N__10815),
            .I(N__10734));
    Span4Mux_v I__2579 (
            .O(N__10812),
            .I(N__10734));
    Span4Mux_v I__2578 (
            .O(N__10809),
            .I(N__10727));
    LocalMux I__2577 (
            .O(N__10806),
            .I(N__10727));
    LocalMux I__2576 (
            .O(N__10803),
            .I(N__10727));
    LocalMux I__2575 (
            .O(N__10796),
            .I(N__10724));
    InMux I__2574 (
            .O(N__10795),
            .I(N__10717));
    InMux I__2573 (
            .O(N__10794),
            .I(N__10717));
    InMux I__2572 (
            .O(N__10793),
            .I(N__10717));
    Span4Mux_v I__2571 (
            .O(N__10788),
            .I(N__10710));
    Span4Mux_h I__2570 (
            .O(N__10785),
            .I(N__10710));
    LocalMux I__2569 (
            .O(N__10774),
            .I(N__10710));
    Span4Mux_h I__2568 (
            .O(N__10771),
            .I(N__10705));
    LocalMux I__2567 (
            .O(N__10766),
            .I(N__10705));
    InMux I__2566 (
            .O(N__10765),
            .I(N__10696));
    InMux I__2565 (
            .O(N__10764),
            .I(N__10696));
    InMux I__2564 (
            .O(N__10763),
            .I(N__10696));
    InMux I__2563 (
            .O(N__10762),
            .I(N__10696));
    Span12Mux_h I__2562 (
            .O(N__10759),
            .I(N__10693));
    Sp12to4 I__2561 (
            .O(N__10756),
            .I(N__10690));
    Span12Mux_h I__2560 (
            .O(N__10753),
            .I(N__10683));
    Sp12to4 I__2559 (
            .O(N__10750),
            .I(N__10683));
    LocalMux I__2558 (
            .O(N__10747),
            .I(N__10683));
    LocalMux I__2557 (
            .O(N__10742),
            .I(N__10680));
    Span4Mux_v I__2556 (
            .O(N__10739),
            .I(N__10677));
    Span4Mux_h I__2555 (
            .O(N__10734),
            .I(N__10674));
    Span4Mux_h I__2554 (
            .O(N__10727),
            .I(N__10667));
    Span4Mux_v I__2553 (
            .O(N__10724),
            .I(N__10667));
    LocalMux I__2552 (
            .O(N__10717),
            .I(N__10667));
    Span4Mux_v I__2551 (
            .O(N__10710),
            .I(N__10660));
    Span4Mux_h I__2550 (
            .O(N__10705),
            .I(N__10660));
    LocalMux I__2549 (
            .O(N__10696),
            .I(N__10660));
    Span12Mux_v I__2548 (
            .O(N__10693),
            .I(N__10657));
    Span12Mux_v I__2547 (
            .O(N__10690),
            .I(N__10650));
    Span12Mux_h I__2546 (
            .O(N__10683),
            .I(N__10650));
    Span12Mux_v I__2545 (
            .O(N__10680),
            .I(N__10650));
    Span4Mux_h I__2544 (
            .O(N__10677),
            .I(N__10645));
    Span4Mux_v I__2543 (
            .O(N__10674),
            .I(N__10645));
    Span4Mux_v I__2542 (
            .O(N__10667),
            .I(N__10640));
    Span4Mux_v I__2541 (
            .O(N__10660),
            .I(N__10640));
    Odrv12 I__2540 (
            .O(N__10657),
            .I(BGn_c));
    Odrv12 I__2539 (
            .O(N__10650),
            .I(BGn_c));
    Odrv4 I__2538 (
            .O(N__10645),
            .I(BGn_c));
    Odrv4 I__2537 (
            .O(N__10640),
            .I(BGn_c));
    InMux I__2536 (
            .O(N__10631),
            .I(N__10628));
    LocalMux I__2535 (
            .O(N__10628),
            .I(N__10611));
    ClkMux I__2534 (
            .O(N__10627),
            .I(N__10448));
    ClkMux I__2533 (
            .O(N__10626),
            .I(N__10448));
    ClkMux I__2532 (
            .O(N__10625),
            .I(N__10448));
    ClkMux I__2531 (
            .O(N__10624),
            .I(N__10448));
    ClkMux I__2530 (
            .O(N__10623),
            .I(N__10448));
    ClkMux I__2529 (
            .O(N__10622),
            .I(N__10448));
    ClkMux I__2528 (
            .O(N__10621),
            .I(N__10448));
    ClkMux I__2527 (
            .O(N__10620),
            .I(N__10448));
    ClkMux I__2526 (
            .O(N__10619),
            .I(N__10448));
    ClkMux I__2525 (
            .O(N__10618),
            .I(N__10448));
    ClkMux I__2524 (
            .O(N__10617),
            .I(N__10448));
    ClkMux I__2523 (
            .O(N__10616),
            .I(N__10448));
    ClkMux I__2522 (
            .O(N__10615),
            .I(N__10448));
    ClkMux I__2521 (
            .O(N__10614),
            .I(N__10448));
    Glb2LocalMux I__2520 (
            .O(N__10611),
            .I(N__10448));
    ClkMux I__2519 (
            .O(N__10610),
            .I(N__10448));
    ClkMux I__2518 (
            .O(N__10609),
            .I(N__10448));
    ClkMux I__2517 (
            .O(N__10608),
            .I(N__10448));
    ClkMux I__2516 (
            .O(N__10607),
            .I(N__10448));
    ClkMux I__2515 (
            .O(N__10606),
            .I(N__10448));
    ClkMux I__2514 (
            .O(N__10605),
            .I(N__10448));
    ClkMux I__2513 (
            .O(N__10604),
            .I(N__10448));
    ClkMux I__2512 (
            .O(N__10603),
            .I(N__10448));
    ClkMux I__2511 (
            .O(N__10602),
            .I(N__10448));
    ClkMux I__2510 (
            .O(N__10601),
            .I(N__10448));
    ClkMux I__2509 (
            .O(N__10600),
            .I(N__10448));
    ClkMux I__2508 (
            .O(N__10599),
            .I(N__10448));
    ClkMux I__2507 (
            .O(N__10598),
            .I(N__10448));
    ClkMux I__2506 (
            .O(N__10597),
            .I(N__10448));
    ClkMux I__2505 (
            .O(N__10596),
            .I(N__10448));
    ClkMux I__2504 (
            .O(N__10595),
            .I(N__10448));
    ClkMux I__2503 (
            .O(N__10594),
            .I(N__10448));
    ClkMux I__2502 (
            .O(N__10593),
            .I(N__10448));
    ClkMux I__2501 (
            .O(N__10592),
            .I(N__10448));
    ClkMux I__2500 (
            .O(N__10591),
            .I(N__10448));
    ClkMux I__2499 (
            .O(N__10590),
            .I(N__10448));
    ClkMux I__2498 (
            .O(N__10589),
            .I(N__10448));
    ClkMux I__2497 (
            .O(N__10588),
            .I(N__10448));
    ClkMux I__2496 (
            .O(N__10587),
            .I(N__10448));
    ClkMux I__2495 (
            .O(N__10586),
            .I(N__10448));
    ClkMux I__2494 (
            .O(N__10585),
            .I(N__10448));
    ClkMux I__2493 (
            .O(N__10584),
            .I(N__10448));
    ClkMux I__2492 (
            .O(N__10583),
            .I(N__10448));
    ClkMux I__2491 (
            .O(N__10582),
            .I(N__10448));
    ClkMux I__2490 (
            .O(N__10581),
            .I(N__10448));
    ClkMux I__2489 (
            .O(N__10580),
            .I(N__10448));
    ClkMux I__2488 (
            .O(N__10579),
            .I(N__10448));
    ClkMux I__2487 (
            .O(N__10578),
            .I(N__10448));
    ClkMux I__2486 (
            .O(N__10577),
            .I(N__10448));
    ClkMux I__2485 (
            .O(N__10576),
            .I(N__10448));
    ClkMux I__2484 (
            .O(N__10575),
            .I(N__10448));
    ClkMux I__2483 (
            .O(N__10574),
            .I(N__10448));
    ClkMux I__2482 (
            .O(N__10573),
            .I(N__10448));
    ClkMux I__2481 (
            .O(N__10572),
            .I(N__10448));
    ClkMux I__2480 (
            .O(N__10571),
            .I(N__10448));
    ClkMux I__2479 (
            .O(N__10570),
            .I(N__10448));
    ClkMux I__2478 (
            .O(N__10569),
            .I(N__10448));
    ClkMux I__2477 (
            .O(N__10568),
            .I(N__10448));
    ClkMux I__2476 (
            .O(N__10567),
            .I(N__10448));
    GlobalMux I__2475 (
            .O(N__10448),
            .I(CLK40));
    CEMux I__2474 (
            .O(N__10445),
            .I(N__10325));
    CEMux I__2473 (
            .O(N__10444),
            .I(N__10325));
    CEMux I__2472 (
            .O(N__10443),
            .I(N__10325));
    CEMux I__2471 (
            .O(N__10442),
            .I(N__10325));
    CEMux I__2470 (
            .O(N__10441),
            .I(N__10325));
    CEMux I__2469 (
            .O(N__10440),
            .I(N__10325));
    CEMux I__2468 (
            .O(N__10439),
            .I(N__10325));
    CEMux I__2467 (
            .O(N__10438),
            .I(N__10325));
    CEMux I__2466 (
            .O(N__10437),
            .I(N__10325));
    CEMux I__2465 (
            .O(N__10436),
            .I(N__10325));
    CEMux I__2464 (
            .O(N__10435),
            .I(N__10325));
    CEMux I__2463 (
            .O(N__10434),
            .I(N__10325));
    CEMux I__2462 (
            .O(N__10433),
            .I(N__10325));
    CEMux I__2461 (
            .O(N__10432),
            .I(N__10325));
    CEMux I__2460 (
            .O(N__10431),
            .I(N__10325));
    CEMux I__2459 (
            .O(N__10430),
            .I(N__10325));
    CEMux I__2458 (
            .O(N__10429),
            .I(N__10325));
    CEMux I__2457 (
            .O(N__10428),
            .I(N__10325));
    CEMux I__2456 (
            .O(N__10427),
            .I(N__10325));
    CEMux I__2455 (
            .O(N__10426),
            .I(N__10325));
    CEMux I__2454 (
            .O(N__10425),
            .I(N__10325));
    CEMux I__2453 (
            .O(N__10424),
            .I(N__10325));
    CEMux I__2452 (
            .O(N__10423),
            .I(N__10325));
    CEMux I__2451 (
            .O(N__10422),
            .I(N__10325));
    CEMux I__2450 (
            .O(N__10421),
            .I(N__10325));
    CEMux I__2449 (
            .O(N__10420),
            .I(N__10325));
    CEMux I__2448 (
            .O(N__10419),
            .I(N__10325));
    CEMux I__2447 (
            .O(N__10418),
            .I(N__10325));
    CEMux I__2446 (
            .O(N__10417),
            .I(N__10325));
    CEMux I__2445 (
            .O(N__10416),
            .I(N__10325));
    CEMux I__2444 (
            .O(N__10415),
            .I(N__10325));
    CEMux I__2443 (
            .O(N__10414),
            .I(N__10325));
    CEMux I__2442 (
            .O(N__10413),
            .I(N__10325));
    CEMux I__2441 (
            .O(N__10412),
            .I(N__10325));
    CEMux I__2440 (
            .O(N__10411),
            .I(N__10325));
    CEMux I__2439 (
            .O(N__10410),
            .I(N__10325));
    CEMux I__2438 (
            .O(N__10409),
            .I(N__10325));
    CEMux I__2437 (
            .O(N__10408),
            .I(N__10325));
    CEMux I__2436 (
            .O(N__10407),
            .I(N__10325));
    CEMux I__2435 (
            .O(N__10406),
            .I(N__10325));
    GlobalMux I__2434 (
            .O(N__10325),
            .I(N__10322));
    gio2CtrlBuf I__2433 (
            .O(N__10322),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    InMux I__2432 (
            .O(N__10319),
            .I(N__10316));
    LocalMux I__2431 (
            .O(N__10316),
            .I(N__10266));
    SRMux I__2430 (
            .O(N__10315),
            .I(N__10169));
    SRMux I__2429 (
            .O(N__10314),
            .I(N__10169));
    SRMux I__2428 (
            .O(N__10313),
            .I(N__10169));
    SRMux I__2427 (
            .O(N__10312),
            .I(N__10169));
    SRMux I__2426 (
            .O(N__10311),
            .I(N__10169));
    SRMux I__2425 (
            .O(N__10310),
            .I(N__10169));
    SRMux I__2424 (
            .O(N__10309),
            .I(N__10169));
    SRMux I__2423 (
            .O(N__10308),
            .I(N__10169));
    SRMux I__2422 (
            .O(N__10307),
            .I(N__10169));
    SRMux I__2421 (
            .O(N__10306),
            .I(N__10169));
    SRMux I__2420 (
            .O(N__10305),
            .I(N__10169));
    SRMux I__2419 (
            .O(N__10304),
            .I(N__10169));
    SRMux I__2418 (
            .O(N__10303),
            .I(N__10169));
    SRMux I__2417 (
            .O(N__10302),
            .I(N__10169));
    SRMux I__2416 (
            .O(N__10301),
            .I(N__10169));
    SRMux I__2415 (
            .O(N__10300),
            .I(N__10169));
    SRMux I__2414 (
            .O(N__10299),
            .I(N__10169));
    SRMux I__2413 (
            .O(N__10298),
            .I(N__10169));
    SRMux I__2412 (
            .O(N__10297),
            .I(N__10169));
    SRMux I__2411 (
            .O(N__10296),
            .I(N__10169));
    SRMux I__2410 (
            .O(N__10295),
            .I(N__10169));
    SRMux I__2409 (
            .O(N__10294),
            .I(N__10169));
    SRMux I__2408 (
            .O(N__10293),
            .I(N__10169));
    SRMux I__2407 (
            .O(N__10292),
            .I(N__10169));
    SRMux I__2406 (
            .O(N__10291),
            .I(N__10169));
    SRMux I__2405 (
            .O(N__10290),
            .I(N__10169));
    SRMux I__2404 (
            .O(N__10289),
            .I(N__10169));
    SRMux I__2403 (
            .O(N__10288),
            .I(N__10169));
    SRMux I__2402 (
            .O(N__10287),
            .I(N__10169));
    SRMux I__2401 (
            .O(N__10286),
            .I(N__10169));
    SRMux I__2400 (
            .O(N__10285),
            .I(N__10169));
    SRMux I__2399 (
            .O(N__10284),
            .I(N__10169));
    SRMux I__2398 (
            .O(N__10283),
            .I(N__10169));
    SRMux I__2397 (
            .O(N__10282),
            .I(N__10169));
    SRMux I__2396 (
            .O(N__10281),
            .I(N__10169));
    SRMux I__2395 (
            .O(N__10280),
            .I(N__10169));
    SRMux I__2394 (
            .O(N__10279),
            .I(N__10169));
    SRMux I__2393 (
            .O(N__10278),
            .I(N__10169));
    SRMux I__2392 (
            .O(N__10277),
            .I(N__10169));
    SRMux I__2391 (
            .O(N__10276),
            .I(N__10169));
    SRMux I__2390 (
            .O(N__10275),
            .I(N__10169));
    SRMux I__2389 (
            .O(N__10274),
            .I(N__10169));
    SRMux I__2388 (
            .O(N__10273),
            .I(N__10169));
    SRMux I__2387 (
            .O(N__10272),
            .I(N__10169));
    SRMux I__2386 (
            .O(N__10271),
            .I(N__10169));
    SRMux I__2385 (
            .O(N__10270),
            .I(N__10169));
    SRMux I__2384 (
            .O(N__10269),
            .I(N__10169));
    Glb2LocalMux I__2383 (
            .O(N__10266),
            .I(N__10169));
    GlobalMux I__2382 (
            .O(N__10169),
            .I(N__10166));
    gio2CtrlBuf I__2381 (
            .O(N__10166),
            .I(RESETn_c_i_g));
    InMux I__2380 (
            .O(N__10163),
            .I(N__10160));
    LocalMux I__2379 (
            .O(N__10160),
            .I(READ_CYCLE_ACTIVE_rep1_i_ess));
    IoInMux I__2378 (
            .O(N__10157),
            .I(N__10154));
    LocalMux I__2377 (
            .O(N__10154),
            .I(N__10151));
    IoSpan4Mux I__2376 (
            .O(N__10151),
            .I(N__10148));
    Span4Mux_s3_h I__2375 (
            .O(N__10148),
            .I(N__10145));
    Odrv4 I__2374 (
            .O(N__10145),
            .I(N_181_i));
    InMux I__2373 (
            .O(N__10142),
            .I(N__10139));
    LocalMux I__2372 (
            .O(N__10139),
            .I(READ_CYCLE_ACTIVE_rep12_i_ess));
    IoInMux I__2371 (
            .O(N__10136),
            .I(N__10133));
    LocalMux I__2370 (
            .O(N__10133),
            .I(N__10130));
    Span4Mux_s2_v I__2369 (
            .O(N__10130),
            .I(N__10127));
    Span4Mux_v I__2368 (
            .O(N__10127),
            .I(N__10124));
    Odrv4 I__2367 (
            .O(N__10124),
            .I(N_192_i));
    InMux I__2366 (
            .O(N__10121),
            .I(N__10118));
    LocalMux I__2365 (
            .O(N__10118),
            .I(READ_CYCLE_ACTIVE_rep14_i_ess));
    InMux I__2364 (
            .O(N__10115),
            .I(N__10112));
    LocalMux I__2363 (
            .O(N__10112),
            .I(READ_CYCLE_ACTIVE_rep10_i_ess));
    InMux I__2362 (
            .O(N__10109),
            .I(N__10106));
    LocalMux I__2361 (
            .O(N__10106),
            .I(READ_CYCLE_ACTIVE_rep22_i_ess));
    IoInMux I__2360 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__2359 (
            .O(N__10100),
            .I(N__10097));
    Span4Mux_s3_h I__2358 (
            .O(N__10097),
            .I(N__10094));
    Odrv4 I__2357 (
            .O(N__10094),
            .I(N_202_i));
    InMux I__2356 (
            .O(N__10091),
            .I(N__10088));
    LocalMux I__2355 (
            .O(N__10088),
            .I(N__10085));
    Odrv4 I__2354 (
            .O(N__10085),
            .I(READ_CYCLE_ACTIVE_rep23_i_ess));
    IoInMux I__2353 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__2352 (
            .O(N__10079),
            .I(N__10076));
    Span4Mux_s3_h I__2351 (
            .O(N__10076),
            .I(N__10073));
    Odrv4 I__2350 (
            .O(N__10073),
            .I(N_203_i));
    InMux I__2349 (
            .O(N__10070),
            .I(N__10067));
    LocalMux I__2348 (
            .O(N__10067),
            .I(READ_CYCLE_ACTIVE_rep18_i_ess));
    InMux I__2347 (
            .O(N__10064),
            .I(N__10061));
    LocalMux I__2346 (
            .O(N__10061),
            .I(N__10058));
    Odrv4 I__2345 (
            .O(N__10058),
            .I(READ_CYCLE_ACTIVE_rep17_i_ess));
    IoInMux I__2344 (
            .O(N__10055),
            .I(N__10052));
    LocalMux I__2343 (
            .O(N__10052),
            .I(N__10049));
    IoSpan4Mux I__2342 (
            .O(N__10049),
            .I(N__10046));
    Span4Mux_s2_h I__2341 (
            .O(N__10046),
            .I(N__10043));
    Odrv4 I__2340 (
            .O(N__10043),
            .I(N_200_i));
    IoInMux I__2339 (
            .O(N__10040),
            .I(N__10037));
    LocalMux I__2338 (
            .O(N__10037),
            .I(N__10034));
    Odrv12 I__2337 (
            .O(N__10034),
            .I(N_188_i));
    InMux I__2336 (
            .O(N__10031),
            .I(N__10028));
    LocalMux I__2335 (
            .O(N__10028),
            .I(READ_CYCLE_ACTIVE_rep21_i_ess));
    IoInMux I__2334 (
            .O(N__10025),
            .I(N__10022));
    LocalMux I__2333 (
            .O(N__10022),
            .I(N__10019));
    Odrv12 I__2332 (
            .O(N__10019),
            .I(N_201_i));
    InMux I__2331 (
            .O(N__10016),
            .I(N__10013));
    LocalMux I__2330 (
            .O(N__10013),
            .I(READ_CYCLE_ACTIVE_rep20_i_ess));
    InMux I__2329 (
            .O(N__10010),
            .I(N__10007));
    LocalMux I__2328 (
            .O(N__10007),
            .I(READ_CYCLE_ACTIVE_rep8_i_ess));
    IoInMux I__2327 (
            .O(N__10004),
            .I(N__10001));
    LocalMux I__2326 (
            .O(N__10001),
            .I(N__9998));
    Span4Mux_s3_h I__2325 (
            .O(N__9998),
            .I(N__9995));
    Odrv4 I__2324 (
            .O(N__9995),
            .I(N_190_i));
    IoInMux I__2323 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__2322 (
            .O(N__9989),
            .I(N__9986));
    Span4Mux_s3_h I__2321 (
            .O(N__9986),
            .I(N__9983));
    Odrv4 I__2320 (
            .O(N__9983),
            .I(N_194_i));
    InMux I__2319 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__2318 (
            .O(N__9977),
            .I(READ_CYCLE_ACTIVE_rep29_i_ess));
    InMux I__2317 (
            .O(N__9974),
            .I(N__9971));
    LocalMux I__2316 (
            .O(N__9971),
            .I(READ_CYCLE_ACTIVE_rep24_i_ess));
    InMux I__2315 (
            .O(N__9968),
            .I(N__9965));
    LocalMux I__2314 (
            .O(N__9965),
            .I(READ_CYCLE_ACTIVE_rep26_i_ess));
    IoInMux I__2313 (
            .O(N__9962),
            .I(N__9959));
    LocalMux I__2312 (
            .O(N__9959),
            .I(N__9956));
    Span4Mux_s3_h I__2311 (
            .O(N__9956),
            .I(N__9953));
    Span4Mux_v I__2310 (
            .O(N__9953),
            .I(N__9950));
    Odrv4 I__2309 (
            .O(N__9950),
            .I(N_197_i));
    IoInMux I__2308 (
            .O(N__9947),
            .I(N__9944));
    LocalMux I__2307 (
            .O(N__9944),
            .I(N__9941));
    IoSpan4Mux I__2306 (
            .O(N__9941),
            .I(N__9938));
    Span4Mux_s0_h I__2305 (
            .O(N__9938),
            .I(N__9935));
    Span4Mux_v I__2304 (
            .O(N__9935),
            .I(N__9932));
    Odrv4 I__2303 (
            .O(N__9932),
            .I(N_211_i));
    IoInMux I__2302 (
            .O(N__9929),
            .I(N__9926));
    LocalMux I__2301 (
            .O(N__9926),
            .I(N__9923));
    Span4Mux_s3_h I__2300 (
            .O(N__9923),
            .I(N__9920));
    Span4Mux_v I__2299 (
            .O(N__9920),
            .I(N__9917));
    Odrv4 I__2298 (
            .O(N__9917),
            .I(N_198_i));
    IoInMux I__2297 (
            .O(N__9914),
            .I(N__9911));
    LocalMux I__2296 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_s3_h I__2295 (
            .O(N__9908),
            .I(N__9905));
    Odrv4 I__2294 (
            .O(N__9905),
            .I(N_199_i));
    InMux I__2293 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__2292 (
            .O(N__9899),
            .I(N__9896));
    Odrv4 I__2291 (
            .O(N__9896),
            .I(READ_CYCLE_ACTIVE_rep31_i_ess));
    InMux I__2290 (
            .O(N__9893),
            .I(N__9890));
    LocalMux I__2289 (
            .O(N__9890),
            .I(READ_CYCLE_ACTIVE_rep19_i_ess));
    InMux I__2288 (
            .O(N__9887),
            .I(N__9884));
    LocalMux I__2287 (
            .O(N__9884),
            .I(N__9881));
    Odrv12 I__2286 (
            .O(N__9881),
            .I(READ_CYCLE_ACTIVE_rep5_i_ess));
    IoInMux I__2285 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__2284 (
            .O(N__9875),
            .I(N__9872));
    Span4Mux_s2_v I__2283 (
            .O(N__9872),
            .I(N__9869));
    Span4Mux_v I__2282 (
            .O(N__9869),
            .I(N__9866));
    Odrv4 I__2281 (
            .O(N__9866),
            .I(N_185_i));
    InMux I__2280 (
            .O(N__9863),
            .I(N__9860));
    LocalMux I__2279 (
            .O(N__9860),
            .I(READ_CYCLE_ACTIVE_rep13_i_ess));
    IoInMux I__2278 (
            .O(N__9857),
            .I(N__9854));
    LocalMux I__2277 (
            .O(N__9854),
            .I(N__9851));
    Span4Mux_s2_v I__2276 (
            .O(N__9851),
            .I(N__9848));
    Span4Mux_v I__2275 (
            .O(N__9848),
            .I(N__9845));
    Odrv4 I__2274 (
            .O(N__9845),
            .I(N_193_i));
    IoInMux I__2273 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__2272 (
            .O(N__9839),
            .I(N__9836));
    Span4Mux_s3_h I__2271 (
            .O(N__9836),
            .I(N__9833));
    Span4Mux_v I__2270 (
            .O(N__9833),
            .I(N__9830));
    Odrv4 I__2269 (
            .O(N__9830),
            .I(N_208_i));
    InMux I__2268 (
            .O(N__9827),
            .I(N__9824));
    LocalMux I__2267 (
            .O(N__9824),
            .I(READ_CYCLE_ACTIVE_rep28_i_ess));
    IoInMux I__2266 (
            .O(N__9821),
            .I(N__9818));
    LocalMux I__2265 (
            .O(N__9818),
            .I(N__9815));
    IoSpan4Mux I__2264 (
            .O(N__9815),
            .I(N__9812));
    Span4Mux_s3_h I__2263 (
            .O(N__9812),
            .I(N__9809));
    Span4Mux_v I__2262 (
            .O(N__9809),
            .I(N__9806));
    Odrv4 I__2261 (
            .O(N__9806),
            .I(N_204_i));
    InMux I__2260 (
            .O(N__9803),
            .I(N__9800));
    LocalMux I__2259 (
            .O(N__9800),
            .I(READ_CYCLE_ACTIVE_rep30_i_ess));
    IoInMux I__2258 (
            .O(N__9797),
            .I(N__9794));
    LocalMux I__2257 (
            .O(N__9794),
            .I(N__9791));
    IoSpan4Mux I__2256 (
            .O(N__9791),
            .I(N__9788));
    IoSpan4Mux I__2255 (
            .O(N__9788),
            .I(N__9785));
    Span4Mux_s1_h I__2254 (
            .O(N__9785),
            .I(N__9782));
    Odrv4 I__2253 (
            .O(N__9782),
            .I(N_210_i));
    IoInMux I__2252 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__2251 (
            .O(N__9776),
            .I(N__9773));
    Span4Mux_s3_h I__2250 (
            .O(N__9773),
            .I(N__9770));
    Span4Mux_v I__2249 (
            .O(N__9770),
            .I(N__9767));
    Odrv4 I__2248 (
            .O(N__9767),
            .I(N_206_i));
    IoInMux I__2247 (
            .O(N__9764),
            .I(N__9761));
    LocalMux I__2246 (
            .O(N__9761),
            .I(N__9758));
    Span4Mux_s3_h I__2245 (
            .O(N__9758),
            .I(N__9755));
    Span4Mux_v I__2244 (
            .O(N__9755),
            .I(N__9752));
    Odrv4 I__2243 (
            .O(N__9752),
            .I(N_209_i));
    IoInMux I__2242 (
            .O(N__9749),
            .I(N__9746));
    LocalMux I__2241 (
            .O(N__9746),
            .I(N__9743));
    IoSpan4Mux I__2240 (
            .O(N__9743),
            .I(N__9740));
    Span4Mux_s3_v I__2239 (
            .O(N__9740),
            .I(N__9737));
    Span4Mux_v I__2238 (
            .O(N__9737),
            .I(N__9734));
    Odrv4 I__2237 (
            .O(N__9734),
            .I(N_207_i));
    IoInMux I__2236 (
            .O(N__9731),
            .I(N__9728));
    LocalMux I__2235 (
            .O(N__9728),
            .I(N__9725));
    IoSpan4Mux I__2234 (
            .O(N__9725),
            .I(N__9722));
    Span4Mux_s3_v I__2233 (
            .O(N__9722),
            .I(N__9719));
    Span4Mux_v I__2232 (
            .O(N__9719),
            .I(N__9716));
    Odrv4 I__2231 (
            .O(N__9716),
            .I(N_205_i));
    InMux I__2230 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__2229 (
            .O(N__9710),
            .I(READ_CYCLE_ACTIVE_rep27_i_ess));
    InMux I__2228 (
            .O(N__9707),
            .I(N__9704));
    LocalMux I__2227 (
            .O(N__9704),
            .I(N__9701));
    Odrv4 I__2226 (
            .O(N__9701),
            .I(READ_CYCLE_ACTIVE_rep25_i_ess));
    IoInMux I__2225 (
            .O(N__9698),
            .I(N__9695));
    LocalMux I__2224 (
            .O(N__9695),
            .I(N__9692));
    IoSpan4Mux I__2223 (
            .O(N__9692),
            .I(N__9689));
    IoSpan4Mux I__2222 (
            .O(N__9689),
            .I(N__9686));
    Span4Mux_s1_h I__2221 (
            .O(N__9686),
            .I(N__9683));
    Odrv4 I__2220 (
            .O(N__9683),
            .I(N_196_i));
    InMux I__2219 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__2218 (
            .O(N__9677),
            .I(READ_CYCLE_ACTIVE_rep16_i_ess));
    IoInMux I__2217 (
            .O(N__9674),
            .I(N__9671));
    LocalMux I__2216 (
            .O(N__9671),
            .I(N__9668));
    IoSpan4Mux I__2215 (
            .O(N__9668),
            .I(N__9663));
    IoInMux I__2214 (
            .O(N__9667),
            .I(N__9660));
    IoInMux I__2213 (
            .O(N__9666),
            .I(N__9657));
    IoSpan4Mux I__2212 (
            .O(N__9663),
            .I(N__9652));
    LocalMux I__2211 (
            .O(N__9660),
            .I(N__9652));
    LocalMux I__2210 (
            .O(N__9657),
            .I(N__9649));
    IoSpan4Mux I__2209 (
            .O(N__9652),
            .I(N__9646));
    Span12Mux_s0_h I__2208 (
            .O(N__9649),
            .I(N__9643));
    Sp12to4 I__2207 (
            .O(N__9646),
            .I(N__9639));
    Span12Mux_h I__2206 (
            .O(N__9643),
            .I(N__9636));
    IoInMux I__2205 (
            .O(N__9642),
            .I(N__9633));
    Span12Mux_s9_v I__2204 (
            .O(N__9639),
            .I(N__9630));
    Span12Mux_h I__2203 (
            .O(N__9636),
            .I(N__9625));
    LocalMux I__2202 (
            .O(N__9633),
            .I(N__9625));
    Odrv12 I__2201 (
            .O(N__9630),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__2200 (
            .O(N__9625),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__2199 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__2198 (
            .O(N__9617),
            .I(READ_CYCLE_ACTIVE_rep4_i_ess));
    IoInMux I__2197 (
            .O(N__9614),
            .I(N__9611));
    LocalMux I__2196 (
            .O(N__9611),
            .I(N__9608));
    Span4Mux_s2_v I__2195 (
            .O(N__9608),
            .I(N__9605));
    Span4Mux_v I__2194 (
            .O(N__9605),
            .I(N__9602));
    Odrv4 I__2193 (
            .O(N__9602),
            .I(N_184_i));
    InMux I__2192 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__2191 (
            .O(N__9596),
            .I(READ_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__2190 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__2189 (
            .O(N__9590),
            .I(N__9587));
    Span4Mux_s2_v I__2188 (
            .O(N__9587),
            .I(N__9584));
    Span4Mux_v I__2187 (
            .O(N__9584),
            .I(N__9581));
    Odrv4 I__2186 (
            .O(N__9581),
            .I(N_182_i));
    InMux I__2185 (
            .O(N__9578),
            .I(N__9575));
    LocalMux I__2184 (
            .O(N__9575),
            .I(READ_CYCLE_ACTIVE_rep0_i_ess));
    IoInMux I__2183 (
            .O(N__9572),
            .I(N__9569));
    LocalMux I__2182 (
            .O(N__9569),
            .I(N__9566));
    IoSpan4Mux I__2181 (
            .O(N__9566),
            .I(N__9563));
    Span4Mux_s2_v I__2180 (
            .O(N__9563),
            .I(N__9560));
    Span4Mux_v I__2179 (
            .O(N__9560),
            .I(N__9557));
    Odrv4 I__2178 (
            .O(N__9557),
            .I(N_180_i));
    InMux I__2177 (
            .O(N__9554),
            .I(N__9551));
    LocalMux I__2176 (
            .O(N__9551),
            .I(N__9548));
    Odrv4 I__2175 (
            .O(N__9548),
            .I(READ_CYCLE_ACTIVE_rep7_i_ess));
    IoInMux I__2174 (
            .O(N__9545),
            .I(N__9542));
    LocalMux I__2173 (
            .O(N__9542),
            .I(N__9539));
    Span12Mux_s6_v I__2172 (
            .O(N__9539),
            .I(N__9536));
    Odrv12 I__2171 (
            .O(N__9536),
            .I(N_187_i));
    InMux I__2170 (
            .O(N__9533),
            .I(N__9530));
    LocalMux I__2169 (
            .O(N__9530),
            .I(READ_CYCLE_ACTIVE_rep6_i_ess));
    IoInMux I__2168 (
            .O(N__9527),
            .I(N__9524));
    LocalMux I__2167 (
            .O(N__9524),
            .I(N__9521));
    Span4Mux_s2_v I__2166 (
            .O(N__9521),
            .I(N__9518));
    Span4Mux_v I__2165 (
            .O(N__9518),
            .I(N__9515));
    Odrv4 I__2164 (
            .O(N__9515),
            .I(N_186_i));
    InMux I__2163 (
            .O(N__9512),
            .I(N__9508));
    IoInMux I__2162 (
            .O(N__9511),
            .I(N__9505));
    LocalMux I__2161 (
            .O(N__9508),
            .I(N__9502));
    LocalMux I__2160 (
            .O(N__9505),
            .I(N__9499));
    Span4Mux_h I__2159 (
            .O(N__9502),
            .I(N__9496));
    Span12Mux_s9_h I__2158 (
            .O(N__9499),
            .I(N__9493));
    Sp12to4 I__2157 (
            .O(N__9496),
            .I(N__9490));
    Span12Mux_v I__2156 (
            .O(N__9493),
            .I(N__9487));
    Span12Mux_v I__2155 (
            .O(N__9490),
            .I(N__9484));
    Span12Mux_h I__2154 (
            .O(N__9487),
            .I(N__9479));
    Span12Mux_v I__2153 (
            .O(N__9484),
            .I(N__9479));
    Odrv12 I__2152 (
            .O(N__9479),
            .I(D_LM_040_in_2));
    InMux I__2151 (
            .O(N__9476),
            .I(N__9473));
    LocalMux I__2150 (
            .O(N__9473),
            .I(N__9470));
    Span4Mux_v I__2149 (
            .O(N__9470),
            .I(N__9467));
    Span4Mux_h I__2148 (
            .O(N__9467),
            .I(N__9464));
    IoSpan4Mux I__2147 (
            .O(N__9464),
            .I(N__9461));
    Odrv4 I__2146 (
            .O(N__9461),
            .I(D_UU_040_in_2));
    IoInMux I__2145 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__2144 (
            .O(N__9455),
            .I(N__9452));
    IoSpan4Mux I__2143 (
            .O(N__9452),
            .I(N__9449));
    IoSpan4Mux I__2142 (
            .O(N__9449),
            .I(N__9446));
    IoSpan4Mux I__2141 (
            .O(N__9446),
            .I(N__9443));
    Span4Mux_s2_v I__2140 (
            .O(N__9443),
            .I(N__9440));
    Span4Mux_v I__2139 (
            .O(N__9440),
            .I(N__9437));
    Odrv4 I__2138 (
            .O(N__9437),
            .I(un1_D_UU_040_2));
    InMux I__2137 (
            .O(N__9434),
            .I(N__9431));
    LocalMux I__2136 (
            .O(N__9431),
            .I(N__9428));
    Span4Mux_h I__2135 (
            .O(N__9428),
            .I(N__9425));
    Span4Mux_v I__2134 (
            .O(N__9425),
            .I(N__9422));
    Span4Mux_h I__2133 (
            .O(N__9422),
            .I(N__9419));
    Odrv4 I__2132 (
            .O(N__9419),
            .I(D_UU_040_in_0));
    IoInMux I__2131 (
            .O(N__9416),
            .I(N__9413));
    LocalMux I__2130 (
            .O(N__9413),
            .I(N__9409));
    InMux I__2129 (
            .O(N__9412),
            .I(N__9406));
    IoSpan4Mux I__2128 (
            .O(N__9409),
            .I(N__9403));
    LocalMux I__2127 (
            .O(N__9406),
            .I(N__9400));
    IoSpan4Mux I__2126 (
            .O(N__9403),
            .I(N__9397));
    Span4Mux_v I__2125 (
            .O(N__9400),
            .I(N__9394));
    Span4Mux_s2_h I__2124 (
            .O(N__9397),
            .I(N__9391));
    Sp12to4 I__2123 (
            .O(N__9394),
            .I(N__9388));
    Sp12to4 I__2122 (
            .O(N__9391),
            .I(N__9385));
    Span12Mux_h I__2121 (
            .O(N__9388),
            .I(N__9382));
    Span12Mux_h I__2120 (
            .O(N__9385),
            .I(N__9379));
    Span12Mux_v I__2119 (
            .O(N__9382),
            .I(N__9376));
    Span12Mux_h I__2118 (
            .O(N__9379),
            .I(N__9373));
    Span12Mux_v I__2117 (
            .O(N__9376),
            .I(N__9370));
    Odrv12 I__2116 (
            .O(N__9373),
            .I(D_LM_040_in_0));
    Odrv12 I__2115 (
            .O(N__9370),
            .I(D_LM_040_in_0));
    IoInMux I__2114 (
            .O(N__9365),
            .I(N__9362));
    LocalMux I__2113 (
            .O(N__9362),
            .I(N__9359));
    IoSpan4Mux I__2112 (
            .O(N__9359),
            .I(N__9356));
    Sp12to4 I__2111 (
            .O(N__9356),
            .I(N__9353));
    Span12Mux_s6_v I__2110 (
            .O(N__9353),
            .I(N__9350));
    Odrv12 I__2109 (
            .O(N__9350),
            .I(un1_D_UU_040_0));
    IoInMux I__2108 (
            .O(N__9347),
            .I(N__9344));
    LocalMux I__2107 (
            .O(N__9344),
            .I(N__9341));
    IoSpan4Mux I__2106 (
            .O(N__9341),
            .I(N__9338));
    IoSpan4Mux I__2105 (
            .O(N__9338),
            .I(N__9334));
    InMux I__2104 (
            .O(N__9337),
            .I(N__9331));
    Span4Mux_s2_h I__2103 (
            .O(N__9334),
            .I(N__9328));
    LocalMux I__2102 (
            .O(N__9331),
            .I(N__9325));
    Sp12to4 I__2101 (
            .O(N__9328),
            .I(N__9322));
    Span4Mux_v I__2100 (
            .O(N__9325),
            .I(N__9319));
    Span12Mux_h I__2099 (
            .O(N__9322),
            .I(N__9316));
    Sp12to4 I__2098 (
            .O(N__9319),
            .I(N__9313));
    Span12Mux_h I__2097 (
            .O(N__9316),
            .I(N__9310));
    Span12Mux_v I__2096 (
            .O(N__9313),
            .I(N__9307));
    Odrv12 I__2095 (
            .O(N__9310),
            .I(D_LM_040_in_3));
    Odrv12 I__2094 (
            .O(N__9307),
            .I(D_LM_040_in_3));
    InMux I__2093 (
            .O(N__9302),
            .I(N__9299));
    LocalMux I__2092 (
            .O(N__9299),
            .I(N__9296));
    Span4Mux_v I__2091 (
            .O(N__9296),
            .I(N__9293));
    Sp12to4 I__2090 (
            .O(N__9293),
            .I(N__9290));
    Span12Mux_h I__2089 (
            .O(N__9290),
            .I(N__9287));
    Odrv12 I__2088 (
            .O(N__9287),
            .I(D_UU_040_in_3));
    IoInMux I__2087 (
            .O(N__9284),
            .I(N__9281));
    LocalMux I__2086 (
            .O(N__9281),
            .I(N__9278));
    IoSpan4Mux I__2085 (
            .O(N__9278),
            .I(N__9275));
    Span4Mux_s0_v I__2084 (
            .O(N__9275),
            .I(N__9272));
    Span4Mux_h I__2083 (
            .O(N__9272),
            .I(N__9269));
    Sp12to4 I__2082 (
            .O(N__9269),
            .I(N__9266));
    Span12Mux_h I__2081 (
            .O(N__9266),
            .I(N__9263));
    Odrv12 I__2080 (
            .O(N__9263),
            .I(un1_D_UU_040_3));
    InMux I__2079 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__2078 (
            .O(N__9257),
            .I(N__9254));
    Span4Mux_v I__2077 (
            .O(N__9254),
            .I(N__9251));
    Span4Mux_h I__2076 (
            .O(N__9251),
            .I(N__9248));
    Odrv4 I__2075 (
            .O(N__9248),
            .I(D_UU_040_in_4));
    IoInMux I__2074 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__2073 (
            .O(N__9242),
            .I(N__9239));
    Span4Mux_s1_h I__2072 (
            .O(N__9239),
            .I(N__9236));
    Sp12to4 I__2071 (
            .O(N__9236),
            .I(N__9232));
    InMux I__2070 (
            .O(N__9235),
            .I(N__9229));
    Span12Mux_v I__2069 (
            .O(N__9232),
            .I(N__9226));
    LocalMux I__2068 (
            .O(N__9229),
            .I(N__9223));
    Span12Mux_h I__2067 (
            .O(N__9226),
            .I(N__9220));
    Span12Mux_h I__2066 (
            .O(N__9223),
            .I(N__9217));
    Span12Mux_h I__2065 (
            .O(N__9220),
            .I(N__9214));
    Span12Mux_v I__2064 (
            .O(N__9217),
            .I(N__9211));
    Odrv12 I__2063 (
            .O(N__9214),
            .I(D_LM_040_in_4));
    Odrv12 I__2062 (
            .O(N__9211),
            .I(D_LM_040_in_4));
    IoInMux I__2061 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__2060 (
            .O(N__9203),
            .I(N__9200));
    IoSpan4Mux I__2059 (
            .O(N__9200),
            .I(N__9197));
    Span4Mux_s2_v I__2058 (
            .O(N__9197),
            .I(N__9194));
    Span4Mux_v I__2057 (
            .O(N__9194),
            .I(N__9191));
    Sp12to4 I__2056 (
            .O(N__9191),
            .I(N__9188));
    Odrv12 I__2055 (
            .O(N__9188),
            .I(un1_D_UU_040_4));
    InMux I__2054 (
            .O(N__9185),
            .I(N__9182));
    LocalMux I__2053 (
            .O(N__9182),
            .I(N__9179));
    Span12Mux_h I__2052 (
            .O(N__9179),
            .I(N__9176));
    Odrv12 I__2051 (
            .O(N__9176),
            .I(D_UM_040_in_0));
    IoInMux I__2050 (
            .O(N__9173),
            .I(N__9170));
    LocalMux I__2049 (
            .O(N__9170),
            .I(N__9167));
    IoSpan4Mux I__2048 (
            .O(N__9167),
            .I(N__9164));
    Span4Mux_s2_h I__2047 (
            .O(N__9164),
            .I(N__9160));
    InMux I__2046 (
            .O(N__9163),
            .I(N__9157));
    Sp12to4 I__2045 (
            .O(N__9160),
            .I(N__9154));
    LocalMux I__2044 (
            .O(N__9157),
            .I(N__9151));
    Span12Mux_h I__2043 (
            .O(N__9154),
            .I(N__9148));
    Span12Mux_v I__2042 (
            .O(N__9151),
            .I(N__9145));
    Span12Mux_h I__2041 (
            .O(N__9148),
            .I(N__9142));
    Span12Mux_v I__2040 (
            .O(N__9145),
            .I(N__9139));
    Odrv12 I__2039 (
            .O(N__9142),
            .I(D_LL_040_in_0));
    Odrv12 I__2038 (
            .O(N__9139),
            .I(D_LL_040_in_0));
    IoInMux I__2037 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__2036 (
            .O(N__9131),
            .I(N__9128));
    IoSpan4Mux I__2035 (
            .O(N__9128),
            .I(N__9125));
    Span4Mux_s2_h I__2034 (
            .O(N__9125),
            .I(N__9122));
    Span4Mux_h I__2033 (
            .O(N__9122),
            .I(N__9119));
    Span4Mux_h I__2032 (
            .O(N__9119),
            .I(N__9116));
    Sp12to4 I__2031 (
            .O(N__9116),
            .I(N__9113));
    Odrv12 I__2030 (
            .O(N__9113),
            .I(un1_D_UM_040_0));
    InMux I__2029 (
            .O(N__9110),
            .I(N__9107));
    LocalMux I__2028 (
            .O(N__9107),
            .I(N__9104));
    Span4Mux_h I__2027 (
            .O(N__9104),
            .I(N__9101));
    Sp12to4 I__2026 (
            .O(N__9101),
            .I(N__9098));
    Span12Mux_v I__2025 (
            .O(N__9098),
            .I(N__9095));
    Odrv12 I__2024 (
            .O(N__9095),
            .I(D_UM_040_in_3));
    IoInMux I__2023 (
            .O(N__9092),
            .I(N__9088));
    InMux I__2022 (
            .O(N__9091),
            .I(N__9085));
    LocalMux I__2021 (
            .O(N__9088),
            .I(N__9082));
    LocalMux I__2020 (
            .O(N__9085),
            .I(N__9079));
    Span4Mux_s3_h I__2019 (
            .O(N__9082),
            .I(N__9076));
    Span4Mux_v I__2018 (
            .O(N__9079),
            .I(N__9073));
    Sp12to4 I__2017 (
            .O(N__9076),
            .I(N__9070));
    Sp12to4 I__2016 (
            .O(N__9073),
            .I(N__9067));
    Span12Mux_v I__2015 (
            .O(N__9070),
            .I(N__9064));
    Span12Mux_h I__2014 (
            .O(N__9067),
            .I(N__9061));
    Span12Mux_h I__2013 (
            .O(N__9064),
            .I(N__9058));
    Span12Mux_v I__2012 (
            .O(N__9061),
            .I(N__9055));
    Span12Mux_h I__2011 (
            .O(N__9058),
            .I(N__9052));
    Span12Mux_v I__2010 (
            .O(N__9055),
            .I(N__9049));
    Odrv12 I__2009 (
            .O(N__9052),
            .I(D_LL_040_in_3));
    Odrv12 I__2008 (
            .O(N__9049),
            .I(D_LL_040_in_3));
    IoInMux I__2007 (
            .O(N__9044),
            .I(N__9041));
    LocalMux I__2006 (
            .O(N__9041),
            .I(N__9038));
    IoSpan4Mux I__2005 (
            .O(N__9038),
            .I(N__9035));
    Span4Mux_s0_h I__2004 (
            .O(N__9035),
            .I(N__9032));
    Span4Mux_h I__2003 (
            .O(N__9032),
            .I(N__9029));
    Sp12to4 I__2002 (
            .O(N__9029),
            .I(N__9026));
    Span12Mux_h I__2001 (
            .O(N__9026),
            .I(N__9023));
    Odrv12 I__2000 (
            .O(N__9023),
            .I(un1_D_UM_040_3));
    InMux I__1999 (
            .O(N__9020),
            .I(N__9015));
    InMux I__1998 (
            .O(N__9019),
            .I(N__9012));
    InMux I__1997 (
            .O(N__9018),
            .I(N__9009));
    LocalMux I__1996 (
            .O(N__9015),
            .I(N__8994));
    LocalMux I__1995 (
            .O(N__9012),
            .I(N__8988));
    LocalMux I__1994 (
            .O(N__9009),
            .I(N__8988));
    InMux I__1993 (
            .O(N__9008),
            .I(N__8985));
    InMux I__1992 (
            .O(N__9007),
            .I(N__8981));
    InMux I__1991 (
            .O(N__9006),
            .I(N__8976));
    InMux I__1990 (
            .O(N__9005),
            .I(N__8970));
    InMux I__1989 (
            .O(N__9004),
            .I(N__8966));
    InMux I__1988 (
            .O(N__9003),
            .I(N__8960));
    InMux I__1987 (
            .O(N__9002),
            .I(N__8953));
    InMux I__1986 (
            .O(N__9001),
            .I(N__8953));
    InMux I__1985 (
            .O(N__9000),
            .I(N__8948));
    InMux I__1984 (
            .O(N__8999),
            .I(N__8948));
    InMux I__1983 (
            .O(N__8998),
            .I(N__8945));
    InMux I__1982 (
            .O(N__8997),
            .I(N__8942));
    Span4Mux_v I__1981 (
            .O(N__8994),
            .I(N__8939));
    InMux I__1980 (
            .O(N__8993),
            .I(N__8936));
    Span4Mux_v I__1979 (
            .O(N__8988),
            .I(N__8932));
    LocalMux I__1978 (
            .O(N__8985),
            .I(N__8929));
    InMux I__1977 (
            .O(N__8984),
            .I(N__8926));
    LocalMux I__1976 (
            .O(N__8981),
            .I(N__8923));
    InMux I__1975 (
            .O(N__8980),
            .I(N__8920));
    InMux I__1974 (
            .O(N__8979),
            .I(N__8916));
    LocalMux I__1973 (
            .O(N__8976),
            .I(N__8912));
    InMux I__1972 (
            .O(N__8975),
            .I(N__8909));
    InMux I__1971 (
            .O(N__8974),
            .I(N__8906));
    InMux I__1970 (
            .O(N__8973),
            .I(N__8903));
    LocalMux I__1969 (
            .O(N__8970),
            .I(N__8900));
    InMux I__1968 (
            .O(N__8969),
            .I(N__8897));
    LocalMux I__1967 (
            .O(N__8966),
            .I(N__8894));
    InMux I__1966 (
            .O(N__8965),
            .I(N__8891));
    InMux I__1965 (
            .O(N__8964),
            .I(N__8887));
    InMux I__1964 (
            .O(N__8963),
            .I(N__8884));
    LocalMux I__1963 (
            .O(N__8960),
            .I(N__8881));
    InMux I__1962 (
            .O(N__8959),
            .I(N__8878));
    InMux I__1961 (
            .O(N__8958),
            .I(N__8875));
    LocalMux I__1960 (
            .O(N__8953),
            .I(N__8866));
    LocalMux I__1959 (
            .O(N__8948),
            .I(N__8866));
    LocalMux I__1958 (
            .O(N__8945),
            .I(N__8866));
    LocalMux I__1957 (
            .O(N__8942),
            .I(N__8866));
    Span4Mux_h I__1956 (
            .O(N__8939),
            .I(N__8861));
    LocalMux I__1955 (
            .O(N__8936),
            .I(N__8861));
    InMux I__1954 (
            .O(N__8935),
            .I(N__8858));
    Span4Mux_v I__1953 (
            .O(N__8932),
            .I(N__8851));
    Span4Mux_h I__1952 (
            .O(N__8929),
            .I(N__8851));
    LocalMux I__1951 (
            .O(N__8926),
            .I(N__8851));
    Span4Mux_v I__1950 (
            .O(N__8923),
            .I(N__8846));
    LocalMux I__1949 (
            .O(N__8920),
            .I(N__8846));
    InMux I__1948 (
            .O(N__8919),
            .I(N__8843));
    LocalMux I__1947 (
            .O(N__8916),
            .I(N__8840));
    InMux I__1946 (
            .O(N__8915),
            .I(N__8837));
    Span4Mux_h I__1945 (
            .O(N__8912),
            .I(N__8832));
    LocalMux I__1944 (
            .O(N__8909),
            .I(N__8832));
    LocalMux I__1943 (
            .O(N__8906),
            .I(N__8829));
    LocalMux I__1942 (
            .O(N__8903),
            .I(N__8826));
    Span4Mux_h I__1941 (
            .O(N__8900),
            .I(N__8821));
    LocalMux I__1940 (
            .O(N__8897),
            .I(N__8821));
    Span4Mux_v I__1939 (
            .O(N__8894),
            .I(N__8816));
    LocalMux I__1938 (
            .O(N__8891),
            .I(N__8816));
    InMux I__1937 (
            .O(N__8890),
            .I(N__8813));
    LocalMux I__1936 (
            .O(N__8887),
            .I(N__8804));
    LocalMux I__1935 (
            .O(N__8884),
            .I(N__8804));
    Span12Mux_h I__1934 (
            .O(N__8881),
            .I(N__8804));
    LocalMux I__1933 (
            .O(N__8878),
            .I(N__8804));
    LocalMux I__1932 (
            .O(N__8875),
            .I(N__8801));
    Span12Mux_h I__1931 (
            .O(N__8866),
            .I(N__8796));
    Sp12to4 I__1930 (
            .O(N__8861),
            .I(N__8796));
    LocalMux I__1929 (
            .O(N__8858),
            .I(N__8793));
    Span4Mux_v I__1928 (
            .O(N__8851),
            .I(N__8790));
    Span4Mux_h I__1927 (
            .O(N__8846),
            .I(N__8785));
    LocalMux I__1926 (
            .O(N__8843),
            .I(N__8785));
    Span4Mux_h I__1925 (
            .O(N__8840),
            .I(N__8780));
    LocalMux I__1924 (
            .O(N__8837),
            .I(N__8780));
    Span4Mux_v I__1923 (
            .O(N__8832),
            .I(N__8775));
    Span4Mux_h I__1922 (
            .O(N__8829),
            .I(N__8775));
    Span4Mux_h I__1921 (
            .O(N__8826),
            .I(N__8770));
    Span4Mux_v I__1920 (
            .O(N__8821),
            .I(N__8770));
    Span4Mux_h I__1919 (
            .O(N__8816),
            .I(N__8767));
    LocalMux I__1918 (
            .O(N__8813),
            .I(N__8764));
    Span12Mux_v I__1917 (
            .O(N__8804),
            .I(N__8758));
    Span12Mux_v I__1916 (
            .O(N__8801),
            .I(N__8758));
    Span12Mux_v I__1915 (
            .O(N__8796),
            .I(N__8751));
    Span12Mux_v I__1914 (
            .O(N__8793),
            .I(N__8751));
    Sp12to4 I__1913 (
            .O(N__8790),
            .I(N__8751));
    Span4Mux_h I__1912 (
            .O(N__8785),
            .I(N__8746));
    Span4Mux_v I__1911 (
            .O(N__8780),
            .I(N__8746));
    Span4Mux_v I__1910 (
            .O(N__8775),
            .I(N__8737));
    Span4Mux_h I__1909 (
            .O(N__8770),
            .I(N__8737));
    Span4Mux_v I__1908 (
            .O(N__8767),
            .I(N__8737));
    Span4Mux_h I__1907 (
            .O(N__8764),
            .I(N__8737));
    InMux I__1906 (
            .O(N__8763),
            .I(N__8734));
    Odrv12 I__1905 (
            .O(N__8758),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1904 (
            .O(N__8751),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1903 (
            .O(N__8746),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1902 (
            .O(N__8737),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1901 (
            .O(N__8734),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    IoInMux I__1900 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__1899 (
            .O(N__8720),
            .I(N__8717));
    IoSpan4Mux I__1898 (
            .O(N__8717),
            .I(N__8713));
    InMux I__1897 (
            .O(N__8716),
            .I(N__8710));
    Span4Mux_s3_h I__1896 (
            .O(N__8713),
            .I(N__8707));
    LocalMux I__1895 (
            .O(N__8710),
            .I(N__8704));
    Sp12to4 I__1894 (
            .O(N__8707),
            .I(N__8701));
    Span4Mux_h I__1893 (
            .O(N__8704),
            .I(N__8698));
    Span12Mux_v I__1892 (
            .O(N__8701),
            .I(N__8695));
    Sp12to4 I__1891 (
            .O(N__8698),
            .I(N__8692));
    Span12Mux_h I__1890 (
            .O(N__8695),
            .I(N__8689));
    Span12Mux_v I__1889 (
            .O(N__8692),
            .I(N__8686));
    Span12Mux_h I__1888 (
            .O(N__8689),
            .I(N__8683));
    Span12Mux_v I__1887 (
            .O(N__8686),
            .I(N__8680));
    Odrv12 I__1886 (
            .O(N__8683),
            .I(D_LL_040_in_7));
    Odrv12 I__1885 (
            .O(N__8680),
            .I(D_LL_040_in_7));
    InMux I__1884 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__1883 (
            .O(N__8672),
            .I(N__8669));
    Span4Mux_v I__1882 (
            .O(N__8669),
            .I(N__8666));
    Span4Mux_v I__1881 (
            .O(N__8666),
            .I(N__8663));
    Sp12to4 I__1880 (
            .O(N__8663),
            .I(N__8660));
    Odrv12 I__1879 (
            .O(N__8660),
            .I(D_UM_040_in_7));
    IoInMux I__1878 (
            .O(N__8657),
            .I(N__8654));
    LocalMux I__1877 (
            .O(N__8654),
            .I(N__8651));
    Span4Mux_s1_h I__1876 (
            .O(N__8651),
            .I(N__8648));
    Span4Mux_h I__1875 (
            .O(N__8648),
            .I(N__8645));
    Span4Mux_h I__1874 (
            .O(N__8645),
            .I(N__8642));
    Span4Mux_h I__1873 (
            .O(N__8642),
            .I(N__8639));
    Span4Mux_h I__1872 (
            .O(N__8639),
            .I(N__8636));
    Span4Mux_h I__1871 (
            .O(N__8636),
            .I(N__8633));
    Odrv4 I__1870 (
            .O(N__8633),
            .I(un1_D_UM_040_7));
    InMux I__1869 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__1868 (
            .O(N__8627),
            .I(N__8624));
    Span4Mux_v I__1867 (
            .O(N__8624),
            .I(N__8621));
    Odrv4 I__1866 (
            .O(N__8621),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1865 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__1864 (
            .O(N__8615),
            .I(N__8611));
    InMux I__1863 (
            .O(N__8614),
            .I(N__8608));
    Span4Mux_v I__1862 (
            .O(N__8611),
            .I(N__8603));
    LocalMux I__1861 (
            .O(N__8608),
            .I(N__8603));
    Sp12to4 I__1860 (
            .O(N__8603),
            .I(N__8599));
    InMux I__1859 (
            .O(N__8602),
            .I(N__8596));
    Span12Mux_v I__1858 (
            .O(N__8599),
            .I(N__8593));
    LocalMux I__1857 (
            .O(N__8596),
            .I(N__8590));
    Span12Mux_h I__1856 (
            .O(N__8593),
            .I(N__8587));
    Span12Mux_v I__1855 (
            .O(N__8590),
            .I(N__8584));
    Odrv12 I__1854 (
            .O(N__8587),
            .I(D_UU_AMIGA_in_5));
    Odrv12 I__1853 (
            .O(N__8584),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1852 (
            .O(N__8579),
            .I(N__8576));
    LocalMux I__1851 (
            .O(N__8576),
            .I(N__8573));
    Span4Mux_s3_v I__1850 (
            .O(N__8573),
            .I(N__8570));
    Span4Mux_v I__1849 (
            .O(N__8570),
            .I(N__8567));
    Sp12to4 I__1848 (
            .O(N__8567),
            .I(N__8564));
    Odrv12 I__1847 (
            .O(N__8564),
            .I(un1_D_UU_AMIGA_5));
    InMux I__1846 (
            .O(N__8561),
            .I(N__8558));
    LocalMux I__1845 (
            .O(N__8558),
            .I(N__8555));
    Odrv12 I__1844 (
            .O(N__8555),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    InMux I__1843 (
            .O(N__8552),
            .I(N__8548));
    InMux I__1842 (
            .O(N__8551),
            .I(N__8545));
    LocalMux I__1841 (
            .O(N__8548),
            .I(N__8541));
    LocalMux I__1840 (
            .O(N__8545),
            .I(N__8538));
    InMux I__1839 (
            .O(N__8544),
            .I(N__8535));
    Span4Mux_v I__1838 (
            .O(N__8541),
            .I(N__8532));
    Span4Mux_v I__1837 (
            .O(N__8538),
            .I(N__8529));
    LocalMux I__1836 (
            .O(N__8535),
            .I(N__8524));
    Sp12to4 I__1835 (
            .O(N__8532),
            .I(N__8524));
    Sp12to4 I__1834 (
            .O(N__8529),
            .I(N__8521));
    Span12Mux_h I__1833 (
            .O(N__8524),
            .I(N__8518));
    Span12Mux_h I__1832 (
            .O(N__8521),
            .I(N__8515));
    Odrv12 I__1831 (
            .O(N__8518),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__1830 (
            .O(N__8515),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1829 (
            .O(N__8510),
            .I(N__8507));
    LocalMux I__1828 (
            .O(N__8507),
            .I(N__8504));
    Span4Mux_s2_v I__1827 (
            .O(N__8504),
            .I(N__8501));
    Span4Mux_v I__1826 (
            .O(N__8501),
            .I(N__8498));
    Sp12to4 I__1825 (
            .O(N__8498),
            .I(N__8495));
    Odrv12 I__1824 (
            .O(N__8495),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1823 (
            .O(N__8492),
            .I(N__8488));
    InMux I__1822 (
            .O(N__8491),
            .I(N__8484));
    LocalMux I__1821 (
            .O(N__8488),
            .I(N__8481));
    InMux I__1820 (
            .O(N__8487),
            .I(N__8478));
    LocalMux I__1819 (
            .O(N__8484),
            .I(N__8475));
    Span4Mux_v I__1818 (
            .O(N__8481),
            .I(N__8470));
    LocalMux I__1817 (
            .O(N__8478),
            .I(N__8470));
    Span4Mux_v I__1816 (
            .O(N__8475),
            .I(N__8467));
    Sp12to4 I__1815 (
            .O(N__8470),
            .I(N__8464));
    Sp12to4 I__1814 (
            .O(N__8467),
            .I(N__8461));
    Span12Mux_h I__1813 (
            .O(N__8464),
            .I(N__8458));
    Span12Mux_h I__1812 (
            .O(N__8461),
            .I(N__8455));
    Odrv12 I__1811 (
            .O(N__8458),
            .I(D_UU_AMIGA_in_6));
    Odrv12 I__1810 (
            .O(N__8455),
            .I(D_UU_AMIGA_in_6));
    InMux I__1809 (
            .O(N__8450),
            .I(N__8447));
    LocalMux I__1808 (
            .O(N__8447),
            .I(N__8434));
    InMux I__1807 (
            .O(N__8446),
            .I(N__8427));
    InMux I__1806 (
            .O(N__8445),
            .I(N__8427));
    InMux I__1805 (
            .O(N__8444),
            .I(N__8427));
    InMux I__1804 (
            .O(N__8443),
            .I(N__8422));
    InMux I__1803 (
            .O(N__8442),
            .I(N__8422));
    InMux I__1802 (
            .O(N__8441),
            .I(N__8417));
    InMux I__1801 (
            .O(N__8440),
            .I(N__8417));
    InMux I__1800 (
            .O(N__8439),
            .I(N__8412));
    InMux I__1799 (
            .O(N__8438),
            .I(N__8412));
    InMux I__1798 (
            .O(N__8437),
            .I(N__8409));
    Span4Mux_v I__1797 (
            .O(N__8434),
            .I(N__8404));
    LocalMux I__1796 (
            .O(N__8427),
            .I(N__8393));
    LocalMux I__1795 (
            .O(N__8422),
            .I(N__8393));
    LocalMux I__1794 (
            .O(N__8417),
            .I(N__8393));
    LocalMux I__1793 (
            .O(N__8412),
            .I(N__8393));
    LocalMux I__1792 (
            .O(N__8409),
            .I(N__8393));
    InMux I__1791 (
            .O(N__8408),
            .I(N__8390));
    InMux I__1790 (
            .O(N__8407),
            .I(N__8387));
    Sp12to4 I__1789 (
            .O(N__8404),
            .I(N__8381));
    Span4Mux_v I__1788 (
            .O(N__8393),
            .I(N__8374));
    LocalMux I__1787 (
            .O(N__8390),
            .I(N__8374));
    LocalMux I__1786 (
            .O(N__8387),
            .I(N__8374));
    InMux I__1785 (
            .O(N__8386),
            .I(N__8369));
    InMux I__1784 (
            .O(N__8385),
            .I(N__8369));
    CascadeMux I__1783 (
            .O(N__8384),
            .I(N__8365));
    Span12Mux_h I__1782 (
            .O(N__8381),
            .I(N__8360));
    Sp12to4 I__1781 (
            .O(N__8374),
            .I(N__8360));
    LocalMux I__1780 (
            .O(N__8369),
            .I(N__8357));
    InMux I__1779 (
            .O(N__8368),
            .I(N__8354));
    InMux I__1778 (
            .O(N__8365),
            .I(N__8351));
    Odrv12 I__1777 (
            .O(N__8360),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__1776 (
            .O(N__8357),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1775 (
            .O(N__8354),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1774 (
            .O(N__8351),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    InMux I__1773 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1772 (
            .O(N__8339),
            .I(N__8336));
    Odrv12 I__1771 (
            .O(N__8336),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    IoInMux I__1770 (
            .O(N__8333),
            .I(N__8330));
    LocalMux I__1769 (
            .O(N__8330),
            .I(N__8327));
    Span12Mux_s8_v I__1768 (
            .O(N__8327),
            .I(N__8324));
    Span12Mux_h I__1767 (
            .O(N__8324),
            .I(N__8321));
    Odrv12 I__1766 (
            .O(N__8321),
            .I(un1_D_UU_AMIGA_6));
    IoInMux I__1765 (
            .O(N__8318),
            .I(N__8315));
    LocalMux I__1764 (
            .O(N__8315),
            .I(N__8312));
    Span4Mux_s2_h I__1763 (
            .O(N__8312),
            .I(N__8309));
    Span4Mux_v I__1762 (
            .O(N__8309),
            .I(N__8305));
    InMux I__1761 (
            .O(N__8308),
            .I(N__8302));
    Sp12to4 I__1760 (
            .O(N__8305),
            .I(N__8299));
    LocalMux I__1759 (
            .O(N__8302),
            .I(N__8296));
    Span12Mux_h I__1758 (
            .O(N__8299),
            .I(N__8293));
    Span12Mux_s11_v I__1757 (
            .O(N__8296),
            .I(N__8290));
    Span12Mux_h I__1756 (
            .O(N__8293),
            .I(N__8287));
    Span12Mux_h I__1755 (
            .O(N__8290),
            .I(N__8284));
    Odrv12 I__1754 (
            .O(N__8287),
            .I(D_LM_040_in_6));
    Odrv12 I__1753 (
            .O(N__8284),
            .I(D_LM_040_in_6));
    InMux I__1752 (
            .O(N__8279),
            .I(N__8276));
    LocalMux I__1751 (
            .O(N__8276),
            .I(N__8273));
    Span4Mux_v I__1750 (
            .O(N__8273),
            .I(N__8270));
    Sp12to4 I__1749 (
            .O(N__8270),
            .I(N__8267));
    Span12Mux_h I__1748 (
            .O(N__8267),
            .I(N__8264));
    Odrv12 I__1747 (
            .O(N__8264),
            .I(D_UU_040_in_6));
    IoInMux I__1746 (
            .O(N__8261),
            .I(N__8258));
    LocalMux I__1745 (
            .O(N__8258),
            .I(N__8255));
    Span4Mux_s3_v I__1744 (
            .O(N__8255),
            .I(N__8252));
    Span4Mux_h I__1743 (
            .O(N__8252),
            .I(N__8249));
    Sp12to4 I__1742 (
            .O(N__8249),
            .I(N__8246));
    Span12Mux_h I__1741 (
            .O(N__8246),
            .I(N__8243));
    Odrv12 I__1740 (
            .O(N__8243),
            .I(un1_D_UU_040_6));
    InMux I__1739 (
            .O(N__8240),
            .I(N__8237));
    LocalMux I__1738 (
            .O(N__8237),
            .I(N__8234));
    Span4Mux_v I__1737 (
            .O(N__8234),
            .I(N__8231));
    Sp12to4 I__1736 (
            .O(N__8231),
            .I(N__8228));
    Span12Mux_h I__1735 (
            .O(N__8228),
            .I(N__8225));
    Odrv12 I__1734 (
            .O(N__8225),
            .I(D_UM_040_in_6));
    IoInMux I__1733 (
            .O(N__8222),
            .I(N__8219));
    LocalMux I__1732 (
            .O(N__8219),
            .I(N__8216));
    IoSpan4Mux I__1731 (
            .O(N__8216),
            .I(N__8212));
    InMux I__1730 (
            .O(N__8215),
            .I(N__8209));
    IoSpan4Mux I__1729 (
            .O(N__8212),
            .I(N__8206));
    LocalMux I__1728 (
            .O(N__8209),
            .I(N__8203));
    Span4Mux_s2_h I__1727 (
            .O(N__8206),
            .I(N__8200));
    Span4Mux_v I__1726 (
            .O(N__8203),
            .I(N__8197));
    Sp12to4 I__1725 (
            .O(N__8200),
            .I(N__8194));
    Sp12to4 I__1724 (
            .O(N__8197),
            .I(N__8191));
    Span12Mux_h I__1723 (
            .O(N__8194),
            .I(N__8188));
    Span12Mux_h I__1722 (
            .O(N__8191),
            .I(N__8185));
    Span12Mux_h I__1721 (
            .O(N__8188),
            .I(N__8182));
    Span12Mux_v I__1720 (
            .O(N__8185),
            .I(N__8179));
    Odrv12 I__1719 (
            .O(N__8182),
            .I(D_LL_040_in_6));
    Odrv12 I__1718 (
            .O(N__8179),
            .I(D_LL_040_in_6));
    IoInMux I__1717 (
            .O(N__8174),
            .I(N__8171));
    LocalMux I__1716 (
            .O(N__8171),
            .I(N__8168));
    Span12Mux_s2_h I__1715 (
            .O(N__8168),
            .I(N__8165));
    Span12Mux_v I__1714 (
            .O(N__8165),
            .I(N__8162));
    Span12Mux_h I__1713 (
            .O(N__8162),
            .I(N__8159));
    Odrv12 I__1712 (
            .O(N__8159),
            .I(un1_D_UM_040_6));
    InMux I__1711 (
            .O(N__8156),
            .I(N__8152));
    IoInMux I__1710 (
            .O(N__8155),
            .I(N__8149));
    LocalMux I__1709 (
            .O(N__8152),
            .I(N__8146));
    LocalMux I__1708 (
            .O(N__8149),
            .I(N__8143));
    Span4Mux_v I__1707 (
            .O(N__8146),
            .I(N__8140));
    Span4Mux_s2_h I__1706 (
            .O(N__8143),
            .I(N__8137));
    Sp12to4 I__1705 (
            .O(N__8140),
            .I(N__8134));
    Span4Mux_v I__1704 (
            .O(N__8137),
            .I(N__8131));
    Span12Mux_h I__1703 (
            .O(N__8134),
            .I(N__8128));
    Sp12to4 I__1702 (
            .O(N__8131),
            .I(N__8125));
    Span12Mux_v I__1701 (
            .O(N__8128),
            .I(N__8122));
    Span12Mux_h I__1700 (
            .O(N__8125),
            .I(N__8119));
    Span12Mux_v I__1699 (
            .O(N__8122),
            .I(N__8114));
    Span12Mux_h I__1698 (
            .O(N__8119),
            .I(N__8114));
    Odrv12 I__1697 (
            .O(N__8114),
            .I(D_LL_040_in_4));
    InMux I__1696 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__1695 (
            .O(N__8108),
            .I(N__8105));
    Span12Mux_v I__1694 (
            .O(N__8105),
            .I(N__8102));
    Span12Mux_h I__1693 (
            .O(N__8102),
            .I(N__8099));
    Odrv12 I__1692 (
            .O(N__8099),
            .I(D_UM_040_in_4));
    IoInMux I__1691 (
            .O(N__8096),
            .I(N__8093));
    LocalMux I__1690 (
            .O(N__8093),
            .I(N__8090));
    Span4Mux_s3_h I__1689 (
            .O(N__8090),
            .I(N__8087));
    Span4Mux_h I__1688 (
            .O(N__8087),
            .I(N__8084));
    Sp12to4 I__1687 (
            .O(N__8084),
            .I(N__8081));
    Span12Mux_s7_v I__1686 (
            .O(N__8081),
            .I(N__8078));
    Odrv12 I__1685 (
            .O(N__8078),
            .I(un1_D_UM_040_4));
    InMux I__1684 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__1683 (
            .O(N__8072),
            .I(N__8069));
    Span4Mux_v I__1682 (
            .O(N__8069),
            .I(N__8066));
    Sp12to4 I__1681 (
            .O(N__8066),
            .I(N__8063));
    Span12Mux_h I__1680 (
            .O(N__8063),
            .I(N__8060));
    Odrv12 I__1679 (
            .O(N__8060),
            .I(D_UM_040_in_5));
    IoInMux I__1678 (
            .O(N__8057),
            .I(N__8054));
    LocalMux I__1677 (
            .O(N__8054),
            .I(N__8051));
    IoSpan4Mux I__1676 (
            .O(N__8051),
            .I(N__8048));
    Span4Mux_s2_h I__1675 (
            .O(N__8048),
            .I(N__8044));
    InMux I__1674 (
            .O(N__8047),
            .I(N__8041));
    Span4Mux_h I__1673 (
            .O(N__8044),
            .I(N__8038));
    LocalMux I__1672 (
            .O(N__8041),
            .I(N__8035));
    Span4Mux_v I__1671 (
            .O(N__8038),
            .I(N__8032));
    Sp12to4 I__1670 (
            .O(N__8035),
            .I(N__8029));
    Sp12to4 I__1669 (
            .O(N__8032),
            .I(N__8026));
    Span12Mux_v I__1668 (
            .O(N__8029),
            .I(N__8023));
    Span12Mux_h I__1667 (
            .O(N__8026),
            .I(N__8018));
    Span12Mux_v I__1666 (
            .O(N__8023),
            .I(N__8018));
    Span12Mux_h I__1665 (
            .O(N__8018),
            .I(N__8015));
    Odrv12 I__1664 (
            .O(N__8015),
            .I(D_LL_040_in_5));
    IoInMux I__1663 (
            .O(N__8012),
            .I(N__8009));
    LocalMux I__1662 (
            .O(N__8009),
            .I(N__8006));
    IoSpan4Mux I__1661 (
            .O(N__8006),
            .I(N__8003));
    IoSpan4Mux I__1660 (
            .O(N__8003),
            .I(N__8000));
    IoSpan4Mux I__1659 (
            .O(N__8000),
            .I(N__7997));
    IoSpan4Mux I__1658 (
            .O(N__7997),
            .I(N__7994));
    Span4Mux_s3_v I__1657 (
            .O(N__7994),
            .I(N__7991));
    Odrv4 I__1656 (
            .O(N__7991),
            .I(un1_D_UM_040_5));
    IoInMux I__1655 (
            .O(N__7988),
            .I(N__7985));
    LocalMux I__1654 (
            .O(N__7985),
            .I(N__7982));
    Span4Mux_s3_h I__1653 (
            .O(N__7982),
            .I(N__7978));
    InMux I__1652 (
            .O(N__7981),
            .I(N__7975));
    Sp12to4 I__1651 (
            .O(N__7978),
            .I(N__7972));
    LocalMux I__1650 (
            .O(N__7975),
            .I(N__7969));
    Span12Mux_v I__1649 (
            .O(N__7972),
            .I(N__7966));
    Span12Mux_v I__1648 (
            .O(N__7969),
            .I(N__7963));
    Span12Mux_h I__1647 (
            .O(N__7966),
            .I(N__7960));
    Span12Mux_v I__1646 (
            .O(N__7963),
            .I(N__7957));
    Span12Mux_h I__1645 (
            .O(N__7960),
            .I(N__7954));
    Span12Mux_h I__1644 (
            .O(N__7957),
            .I(N__7951));
    Odrv12 I__1643 (
            .O(N__7954),
            .I(D_LL_040_in_1));
    Odrv12 I__1642 (
            .O(N__7951),
            .I(D_LL_040_in_1));
    InMux I__1641 (
            .O(N__7946),
            .I(N__7943));
    LocalMux I__1640 (
            .O(N__7943),
            .I(N__7940));
    Span4Mux_h I__1639 (
            .O(N__7940),
            .I(N__7937));
    Sp12to4 I__1638 (
            .O(N__7937),
            .I(N__7934));
    Span12Mux_v I__1637 (
            .O(N__7934),
            .I(N__7931));
    Odrv12 I__1636 (
            .O(N__7931),
            .I(D_UM_040_in_1));
    IoInMux I__1635 (
            .O(N__7928),
            .I(N__7925));
    LocalMux I__1634 (
            .O(N__7925),
            .I(N__7922));
    IoSpan4Mux I__1633 (
            .O(N__7922),
            .I(N__7919));
    Span4Mux_s0_h I__1632 (
            .O(N__7919),
            .I(N__7916));
    Sp12to4 I__1631 (
            .O(N__7916),
            .I(N__7913));
    Span12Mux_s8_h I__1630 (
            .O(N__7913),
            .I(N__7910));
    Odrv12 I__1629 (
            .O(N__7910),
            .I(un1_D_UM_040_1));
    CEMux I__1628 (
            .O(N__7907),
            .I(N__7900));
    CEMux I__1627 (
            .O(N__7906),
            .I(N__7897));
    CEMux I__1626 (
            .O(N__7905),
            .I(N__7894));
    CEMux I__1625 (
            .O(N__7904),
            .I(N__7891));
    CEMux I__1624 (
            .O(N__7903),
            .I(N__7888));
    LocalMux I__1623 (
            .O(N__7900),
            .I(\U111_CYCLE_SM.N_159_0 ));
    LocalMux I__1622 (
            .O(N__7897),
            .I(\U111_CYCLE_SM.N_159_0 ));
    LocalMux I__1621 (
            .O(N__7894),
            .I(\U111_CYCLE_SM.N_159_0 ));
    LocalMux I__1620 (
            .O(N__7891),
            .I(\U111_CYCLE_SM.N_159_0 ));
    LocalMux I__1619 (
            .O(N__7888),
            .I(\U111_CYCLE_SM.N_159_0 ));
    SRMux I__1618 (
            .O(N__7877),
            .I(N__7873));
    SRMux I__1617 (
            .O(N__7876),
            .I(N__7868));
    LocalMux I__1616 (
            .O(N__7873),
            .I(N__7865));
    SRMux I__1615 (
            .O(N__7872),
            .I(N__7862));
    SRMux I__1614 (
            .O(N__7871),
            .I(N__7858));
    LocalMux I__1613 (
            .O(N__7868),
            .I(N__7851));
    Span4Mux_h I__1612 (
            .O(N__7865),
            .I(N__7851));
    LocalMux I__1611 (
            .O(N__7862),
            .I(N__7851));
    SRMux I__1610 (
            .O(N__7861),
            .I(N__7848));
    LocalMux I__1609 (
            .O(N__7858),
            .I(N__7845));
    Span4Mux_v I__1608 (
            .O(N__7851),
            .I(N__7840));
    LocalMux I__1607 (
            .O(N__7848),
            .I(N__7840));
    Span4Mux_h I__1606 (
            .O(N__7845),
            .I(N__7837));
    Span4Mux_h I__1605 (
            .O(N__7840),
            .I(N__7834));
    Odrv4 I__1604 (
            .O(N__7837),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    Odrv4 I__1603 (
            .O(N__7834),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    InMux I__1602 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__1601 (
            .O(N__7826),
            .I(N__7823));
    Span4Mux_v I__1600 (
            .O(N__7823),
            .I(N__7819));
    InMux I__1599 (
            .O(N__7822),
            .I(N__7816));
    Odrv4 I__1598 (
            .O(N__7819),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1597 (
            .O(N__7816),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    IoInMux I__1596 (
            .O(N__7811),
            .I(N__7808));
    LocalMux I__1595 (
            .O(N__7808),
            .I(N__7805));
    Span4Mux_s2_v I__1594 (
            .O(N__7805),
            .I(N__7802));
    Span4Mux_v I__1593 (
            .O(N__7802),
            .I(N__7799));
    Span4Mux_v I__1592 (
            .O(N__7799),
            .I(N__7796));
    Odrv4 I__1591 (
            .O(N__7796),
            .I(TAn_1_i));
    InMux I__1590 (
            .O(N__7793),
            .I(N__7790));
    LocalMux I__1589 (
            .O(N__7790),
            .I(N__7787));
    Odrv4 I__1588 (
            .O(N__7787),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    InMux I__1587 (
            .O(N__7784),
            .I(N__7780));
    InMux I__1586 (
            .O(N__7783),
            .I(N__7777));
    LocalMux I__1585 (
            .O(N__7780),
            .I(N__7774));
    LocalMux I__1584 (
            .O(N__7777),
            .I(N__7770));
    Span4Mux_v I__1583 (
            .O(N__7774),
            .I(N__7767));
    InMux I__1582 (
            .O(N__7773),
            .I(N__7764));
    Span4Mux_v I__1581 (
            .O(N__7770),
            .I(N__7761));
    Span4Mux_h I__1580 (
            .O(N__7767),
            .I(N__7758));
    LocalMux I__1579 (
            .O(N__7764),
            .I(N__7755));
    Sp12to4 I__1578 (
            .O(N__7761),
            .I(N__7752));
    Sp12to4 I__1577 (
            .O(N__7758),
            .I(N__7747));
    Span12Mux_h I__1576 (
            .O(N__7755),
            .I(N__7747));
    Span12Mux_h I__1575 (
            .O(N__7752),
            .I(N__7744));
    Span12Mux_h I__1574 (
            .O(N__7747),
            .I(N__7741));
    Span12Mux_v I__1573 (
            .O(N__7744),
            .I(N__7738));
    Odrv12 I__1572 (
            .O(N__7741),
            .I(D_UU_AMIGA_in_3));
    Odrv12 I__1571 (
            .O(N__7738),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1570 (
            .O(N__7733),
            .I(N__7730));
    LocalMux I__1569 (
            .O(N__7730),
            .I(N__7727));
    Span4Mux_s0_v I__1568 (
            .O(N__7727),
            .I(N__7724));
    Span4Mux_v I__1567 (
            .O(N__7724),
            .I(N__7721));
    Sp12to4 I__1566 (
            .O(N__7721),
            .I(N__7718));
    Span12Mux_h I__1565 (
            .O(N__7718),
            .I(N__7715));
    Odrv12 I__1564 (
            .O(N__7715),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1563 (
            .O(N__7712),
            .I(N__7709));
    LocalMux I__1562 (
            .O(N__7709),
            .I(N__7706));
    Odrv4 I__1561 (
            .O(N__7706),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    InMux I__1560 (
            .O(N__7703),
            .I(N__7699));
    InMux I__1559 (
            .O(N__7702),
            .I(N__7695));
    LocalMux I__1558 (
            .O(N__7699),
            .I(N__7692));
    InMux I__1557 (
            .O(N__7698),
            .I(N__7689));
    LocalMux I__1556 (
            .O(N__7695),
            .I(N__7686));
    Span4Mux_v I__1555 (
            .O(N__7692),
            .I(N__7681));
    LocalMux I__1554 (
            .O(N__7689),
            .I(N__7681));
    Span12Mux_v I__1553 (
            .O(N__7686),
            .I(N__7678));
    Span4Mux_v I__1552 (
            .O(N__7681),
            .I(N__7675));
    Span12Mux_v I__1551 (
            .O(N__7678),
            .I(N__7672));
    Sp12to4 I__1550 (
            .O(N__7675),
            .I(N__7669));
    Span12Mux_h I__1549 (
            .O(N__7672),
            .I(N__7666));
    Span12Mux_h I__1548 (
            .O(N__7669),
            .I(N__7663));
    Odrv12 I__1547 (
            .O(N__7666),
            .I(D_UM_AMIGA_in_3));
    Odrv12 I__1546 (
            .O(N__7663),
            .I(D_UM_AMIGA_in_3));
    IoInMux I__1545 (
            .O(N__7658),
            .I(N__7655));
    LocalMux I__1544 (
            .O(N__7655),
            .I(N__7652));
    IoSpan4Mux I__1543 (
            .O(N__7652),
            .I(N__7649));
    Span4Mux_s1_h I__1542 (
            .O(N__7649),
            .I(N__7646));
    Sp12to4 I__1541 (
            .O(N__7646),
            .I(N__7643));
    Span12Mux_h I__1540 (
            .O(N__7643),
            .I(N__7640));
    Odrv12 I__1539 (
            .O(N__7640),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1538 (
            .O(N__7637),
            .I(N__7633));
    InMux I__1537 (
            .O(N__7636),
            .I(N__7629));
    LocalMux I__1536 (
            .O(N__7633),
            .I(N__7626));
    InMux I__1535 (
            .O(N__7632),
            .I(N__7623));
    LocalMux I__1534 (
            .O(N__7629),
            .I(N__7620));
    Span4Mux_v I__1533 (
            .O(N__7626),
            .I(N__7615));
    LocalMux I__1532 (
            .O(N__7623),
            .I(N__7615));
    Span12Mux_v I__1531 (
            .O(N__7620),
            .I(N__7612));
    Span4Mux_v I__1530 (
            .O(N__7615),
            .I(N__7609));
    Span12Mux_h I__1529 (
            .O(N__7612),
            .I(N__7606));
    Sp12to4 I__1528 (
            .O(N__7609),
            .I(N__7603));
    Span12Mux_v I__1527 (
            .O(N__7606),
            .I(N__7600));
    Span12Mux_h I__1526 (
            .O(N__7603),
            .I(N__7597));
    Odrv12 I__1525 (
            .O(N__7600),
            .I(D_UM_AMIGA_in_4));
    Odrv12 I__1524 (
            .O(N__7597),
            .I(D_UM_AMIGA_in_4));
    InMux I__1523 (
            .O(N__7592),
            .I(N__7589));
    LocalMux I__1522 (
            .O(N__7589),
            .I(N__7586));
    Odrv12 I__1521 (
            .O(N__7586),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    IoInMux I__1520 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__1519 (
            .O(N__7580),
            .I(N__7577));
    IoSpan4Mux I__1518 (
            .O(N__7577),
            .I(N__7574));
    IoSpan4Mux I__1517 (
            .O(N__7574),
            .I(N__7571));
    Span4Mux_s3_v I__1516 (
            .O(N__7571),
            .I(N__7568));
    Span4Mux_h I__1515 (
            .O(N__7568),
            .I(N__7565));
    Span4Mux_v I__1514 (
            .O(N__7565),
            .I(N__7562));
    Odrv4 I__1513 (
            .O(N__7562),
            .I(un1_D_UM_AMIGA_4));
    IoInMux I__1512 (
            .O(N__7559),
            .I(N__7556));
    LocalMux I__1511 (
            .O(N__7556),
            .I(N__7553));
    IoSpan4Mux I__1510 (
            .O(N__7553),
            .I(N__7550));
    Span4Mux_s1_h I__1509 (
            .O(N__7550),
            .I(N__7547));
    Sp12to4 I__1508 (
            .O(N__7547),
            .I(N__7544));
    Span12Mux_h I__1507 (
            .O(N__7544),
            .I(N__7541));
    Odrv12 I__1506 (
            .O(N__7541),
            .I(un1_D_UM_AMIGA_0));
    CascadeMux I__1505 (
            .O(N__7538),
            .I(N__7534));
    InMux I__1504 (
            .O(N__7537),
            .I(N__7530));
    InMux I__1503 (
            .O(N__7534),
            .I(N__7525));
    InMux I__1502 (
            .O(N__7533),
            .I(N__7525));
    LocalMux I__1501 (
            .O(N__7530),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__1500 (
            .O(N__7525),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    CascadeMux I__1499 (
            .O(N__7520),
            .I(N__7517));
    InMux I__1498 (
            .O(N__7517),
            .I(N__7513));
    InMux I__1497 (
            .O(N__7516),
            .I(N__7510));
    LocalMux I__1496 (
            .O(N__7513),
            .I(N__7505));
    LocalMux I__1495 (
            .O(N__7510),
            .I(N__7505));
    Span4Mux_v I__1494 (
            .O(N__7505),
            .I(N__7501));
    InMux I__1493 (
            .O(N__7504),
            .I(N__7498));
    Sp12to4 I__1492 (
            .O(N__7501),
            .I(N__7493));
    LocalMux I__1491 (
            .O(N__7498),
            .I(N__7493));
    Span12Mux_h I__1490 (
            .O(N__7493),
            .I(N__7490));
    Span12Mux_v I__1489 (
            .O(N__7490),
            .I(N__7487));
    Odrv12 I__1488 (
            .O(N__7487),
            .I(PORTSIZE_c));
    InMux I__1487 (
            .O(N__7484),
            .I(N__7481));
    LocalMux I__1486 (
            .O(N__7481),
            .I(N__7477));
    InMux I__1485 (
            .O(N__7480),
            .I(N__7474));
    Span4Mux_v I__1484 (
            .O(N__7477),
            .I(N__7466));
    LocalMux I__1483 (
            .O(N__7474),
            .I(N__7466));
    InMux I__1482 (
            .O(N__7473),
            .I(N__7463));
    InMux I__1481 (
            .O(N__7472),
            .I(N__7460));
    InMux I__1480 (
            .O(N__7471),
            .I(N__7457));
    Odrv4 I__1479 (
            .O(N__7466),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1478 (
            .O(N__7463),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1477 (
            .O(N__7460),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1476 (
            .O(N__7457),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    InMux I__1475 (
            .O(N__7448),
            .I(N__7444));
    InMux I__1474 (
            .O(N__7447),
            .I(N__7440));
    LocalMux I__1473 (
            .O(N__7444),
            .I(N__7436));
    InMux I__1472 (
            .O(N__7443),
            .I(N__7433));
    LocalMux I__1471 (
            .O(N__7440),
            .I(N__7430));
    InMux I__1470 (
            .O(N__7439),
            .I(N__7427));
    Odrv4 I__1469 (
            .O(N__7436),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1468 (
            .O(N__7433),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    Odrv4 I__1467 (
            .O(N__7430),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1466 (
            .O(N__7427),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    IoInMux I__1465 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__1464 (
            .O(N__7415),
            .I(N__7412));
    Span12Mux_s3_h I__1463 (
            .O(N__7412),
            .I(N__7409));
    Span12Mux_h I__1462 (
            .O(N__7409),
            .I(N__7406));
    Odrv12 I__1461 (
            .O(N__7406),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1460 (
            .O(N__7403),
            .I(N__7400));
    LocalMux I__1459 (
            .O(N__7400),
            .I(N__7397));
    Span4Mux_v I__1458 (
            .O(N__7397),
            .I(N__7394));
    Span4Mux_v I__1457 (
            .O(N__7394),
            .I(N__7389));
    InMux I__1456 (
            .O(N__7393),
            .I(N__7386));
    InMux I__1455 (
            .O(N__7392),
            .I(N__7383));
    Sp12to4 I__1454 (
            .O(N__7389),
            .I(N__7378));
    LocalMux I__1453 (
            .O(N__7386),
            .I(N__7378));
    LocalMux I__1452 (
            .O(N__7383),
            .I(N__7375));
    Span12Mux_h I__1451 (
            .O(N__7378),
            .I(N__7372));
    Span12Mux_v I__1450 (
            .O(N__7375),
            .I(N__7369));
    Span12Mux_v I__1449 (
            .O(N__7372),
            .I(N__7366));
    Span12Mux_h I__1448 (
            .O(N__7369),
            .I(N__7363));
    Odrv12 I__1447 (
            .O(N__7366),
            .I(D_UM_AMIGA_in_6));
    Odrv12 I__1446 (
            .O(N__7363),
            .I(D_UM_AMIGA_in_6));
    InMux I__1445 (
            .O(N__7358),
            .I(N__7355));
    LocalMux I__1444 (
            .O(N__7355),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    IoInMux I__1443 (
            .O(N__7352),
            .I(N__7349));
    LocalMux I__1442 (
            .O(N__7349),
            .I(N__7346));
    IoSpan4Mux I__1441 (
            .O(N__7346),
            .I(N__7343));
    Span4Mux_s2_h I__1440 (
            .O(N__7343),
            .I(N__7340));
    Span4Mux_h I__1439 (
            .O(N__7340),
            .I(N__7337));
    Sp12to4 I__1438 (
            .O(N__7337),
            .I(N__7334));
    Odrv12 I__1437 (
            .O(N__7334),
            .I(un1_D_UM_AMIGA_6));
    InMux I__1436 (
            .O(N__7331),
            .I(N__7328));
    LocalMux I__1435 (
            .O(N__7328),
            .I(N__7325));
    Span4Mux_v I__1434 (
            .O(N__7325),
            .I(N__7320));
    InMux I__1433 (
            .O(N__7324),
            .I(N__7317));
    InMux I__1432 (
            .O(N__7323),
            .I(N__7314));
    Span4Mux_v I__1431 (
            .O(N__7320),
            .I(N__7307));
    LocalMux I__1430 (
            .O(N__7317),
            .I(N__7307));
    LocalMux I__1429 (
            .O(N__7314),
            .I(N__7307));
    Span4Mux_v I__1428 (
            .O(N__7307),
            .I(N__7304));
    Sp12to4 I__1427 (
            .O(N__7304),
            .I(N__7301));
    Span12Mux_h I__1426 (
            .O(N__7301),
            .I(N__7298));
    Odrv12 I__1425 (
            .O(N__7298),
            .I(D_UM_AMIGA_in_2));
    InMux I__1424 (
            .O(N__7295),
            .I(N__7292));
    LocalMux I__1423 (
            .O(N__7292),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    InMux I__1422 (
            .O(N__7289),
            .I(N__7286));
    LocalMux I__1421 (
            .O(N__7286),
            .I(N__7283));
    Span4Mux_v I__1420 (
            .O(N__7283),
            .I(N__7278));
    InMux I__1419 (
            .O(N__7282),
            .I(N__7275));
    InMux I__1418 (
            .O(N__7281),
            .I(N__7272));
    Span4Mux_v I__1417 (
            .O(N__7278),
            .I(N__7269));
    LocalMux I__1416 (
            .O(N__7275),
            .I(N__7266));
    LocalMux I__1415 (
            .O(N__7272),
            .I(N__7263));
    Span4Mux_v I__1414 (
            .O(N__7269),
            .I(N__7256));
    Span4Mux_v I__1413 (
            .O(N__7266),
            .I(N__7256));
    Span4Mux_v I__1412 (
            .O(N__7263),
            .I(N__7256));
    Sp12to4 I__1411 (
            .O(N__7256),
            .I(N__7253));
    Span12Mux_h I__1410 (
            .O(N__7253),
            .I(N__7250));
    Odrv12 I__1409 (
            .O(N__7250),
            .I(D_UM_AMIGA_in_0));
    InMux I__1408 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__1407 (
            .O(N__7244),
            .I(N__7241));
    Odrv4 I__1406 (
            .O(N__7241),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__1405 (
            .O(N__7238),
            .I(N__7235));
    LocalMux I__1404 (
            .O(N__7235),
            .I(N__7231));
    InMux I__1403 (
            .O(N__7234),
            .I(N__7228));
    Odrv12 I__1402 (
            .O(N__7231),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1401 (
            .O(N__7228),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    InMux I__1400 (
            .O(N__7223),
            .I(N__7220));
    LocalMux I__1399 (
            .O(N__7220),
            .I(N__7217));
    Odrv12 I__1398 (
            .O(N__7217),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    InMux I__1397 (
            .O(N__7214),
            .I(N__7211));
    LocalMux I__1396 (
            .O(N__7211),
            .I(N__7207));
    InMux I__1395 (
            .O(N__7210),
            .I(N__7204));
    Span4Mux_v I__1394 (
            .O(N__7207),
            .I(N__7201));
    LocalMux I__1393 (
            .O(N__7204),
            .I(N__7197));
    Span4Mux_h I__1392 (
            .O(N__7201),
            .I(N__7194));
    InMux I__1391 (
            .O(N__7200),
            .I(N__7191));
    Sp12to4 I__1390 (
            .O(N__7197),
            .I(N__7188));
    Sp12to4 I__1389 (
            .O(N__7194),
            .I(N__7185));
    LocalMux I__1388 (
            .O(N__7191),
            .I(N__7180));
    Span12Mux_s11_v I__1387 (
            .O(N__7188),
            .I(N__7180));
    Span12Mux_v I__1386 (
            .O(N__7185),
            .I(N__7177));
    Span12Mux_h I__1385 (
            .O(N__7180),
            .I(N__7174));
    Odrv12 I__1384 (
            .O(N__7177),
            .I(D_UM_AMIGA_in_5));
    Odrv12 I__1383 (
            .O(N__7174),
            .I(D_UM_AMIGA_in_5));
    IoInMux I__1382 (
            .O(N__7169),
            .I(N__7166));
    LocalMux I__1381 (
            .O(N__7166),
            .I(N__7163));
    IoSpan4Mux I__1380 (
            .O(N__7163),
            .I(N__7160));
    Span4Mux_s3_v I__1379 (
            .O(N__7160),
            .I(N__7157));
    Span4Mux_h I__1378 (
            .O(N__7157),
            .I(N__7154));
    Span4Mux_h I__1377 (
            .O(N__7154),
            .I(N__7151));
    Span4Mux_v I__1376 (
            .O(N__7151),
            .I(N__7148));
    Odrv4 I__1375 (
            .O(N__7148),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1374 (
            .O(N__7145),
            .I(N__7142));
    LocalMux I__1373 (
            .O(N__7142),
            .I(N__7137));
    InMux I__1372 (
            .O(N__7141),
            .I(N__7134));
    InMux I__1371 (
            .O(N__7140),
            .I(N__7131));
    Span4Mux_v I__1370 (
            .O(N__7137),
            .I(N__7128));
    LocalMux I__1369 (
            .O(N__7134),
            .I(N__7123));
    LocalMux I__1368 (
            .O(N__7131),
            .I(N__7123));
    Sp12to4 I__1367 (
            .O(N__7128),
            .I(N__7120));
    Span12Mux_v I__1366 (
            .O(N__7123),
            .I(N__7117));
    Span12Mux_v I__1365 (
            .O(N__7120),
            .I(N__7114));
    Span12Mux_h I__1364 (
            .O(N__7117),
            .I(N__7111));
    Odrv12 I__1363 (
            .O(N__7114),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1362 (
            .O(N__7111),
            .I(D_UM_AMIGA_in_7));
    InMux I__1361 (
            .O(N__7106),
            .I(N__7103));
    LocalMux I__1360 (
            .O(N__7103),
            .I(N__7100));
    Odrv12 I__1359 (
            .O(N__7100),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1358 (
            .O(N__7097),
            .I(N__7094));
    LocalMux I__1357 (
            .O(N__7094),
            .I(N__7091));
    IoSpan4Mux I__1356 (
            .O(N__7091),
            .I(N__7088));
    Span4Mux_s2_h I__1355 (
            .O(N__7088),
            .I(N__7085));
    Span4Mux_h I__1354 (
            .O(N__7085),
            .I(N__7082));
    Sp12to4 I__1353 (
            .O(N__7082),
            .I(N__7079));
    Span12Mux_s7_v I__1352 (
            .O(N__7079),
            .I(N__7076));
    Odrv12 I__1351 (
            .O(N__7076),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1350 (
            .O(N__7073),
            .I(N__7070));
    LocalMux I__1349 (
            .O(N__7070),
            .I(N__7067));
    Span4Mux_v I__1348 (
            .O(N__7067),
            .I(N__7062));
    InMux I__1347 (
            .O(N__7066),
            .I(N__7059));
    InMux I__1346 (
            .O(N__7065),
            .I(N__7056));
    Span4Mux_v I__1345 (
            .O(N__7062),
            .I(N__7053));
    LocalMux I__1344 (
            .O(N__7059),
            .I(N__7050));
    LocalMux I__1343 (
            .O(N__7056),
            .I(N__7047));
    Span4Mux_v I__1342 (
            .O(N__7053),
            .I(N__7040));
    Span4Mux_v I__1341 (
            .O(N__7050),
            .I(N__7040));
    Span4Mux_v I__1340 (
            .O(N__7047),
            .I(N__7040));
    Sp12to4 I__1339 (
            .O(N__7040),
            .I(N__7037));
    Span12Mux_h I__1338 (
            .O(N__7037),
            .I(N__7034));
    Odrv12 I__1337 (
            .O(N__7034),
            .I(D_UU_AMIGA_in_0));
    InMux I__1336 (
            .O(N__7031),
            .I(N__7028));
    LocalMux I__1335 (
            .O(N__7028),
            .I(N__7025));
    Odrv12 I__1334 (
            .O(N__7025),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    IoInMux I__1333 (
            .O(N__7022),
            .I(N__7019));
    LocalMux I__1332 (
            .O(N__7019),
            .I(N__7016));
    Span12Mux_s9_v I__1331 (
            .O(N__7016),
            .I(N__7013));
    Span12Mux_h I__1330 (
            .O(N__7013),
            .I(N__7010));
    Odrv12 I__1329 (
            .O(N__7010),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1328 (
            .O(N__7007),
            .I(N__7004));
    LocalMux I__1327 (
            .O(N__7004),
            .I(N__7001));
    Span4Mux_v I__1326 (
            .O(N__7001),
            .I(N__6998));
    Odrv4 I__1325 (
            .O(N__6998),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__1324 (
            .O(N__6995),
            .I(N__6990));
    InMux I__1323 (
            .O(N__6994),
            .I(N__6987));
    InMux I__1322 (
            .O(N__6993),
            .I(N__6984));
    LocalMux I__1321 (
            .O(N__6990),
            .I(N__6981));
    LocalMux I__1320 (
            .O(N__6987),
            .I(N__6978));
    LocalMux I__1319 (
            .O(N__6984),
            .I(N__6975));
    Span12Mux_v I__1318 (
            .O(N__6981),
            .I(N__6972));
    Span12Mux_s7_v I__1317 (
            .O(N__6978),
            .I(N__6969));
    Span4Mux_h I__1316 (
            .O(N__6975),
            .I(N__6966));
    Span12Mux_h I__1315 (
            .O(N__6972),
            .I(N__6963));
    Span12Mux_h I__1314 (
            .O(N__6969),
            .I(N__6958));
    Sp12to4 I__1313 (
            .O(N__6966),
            .I(N__6958));
    Odrv12 I__1312 (
            .O(N__6963),
            .I(D_UU_AMIGA_in_7));
    Odrv12 I__1311 (
            .O(N__6958),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1310 (
            .O(N__6953),
            .I(N__6950));
    LocalMux I__1309 (
            .O(N__6950),
            .I(N__6947));
    Span4Mux_s2_v I__1308 (
            .O(N__6947),
            .I(N__6944));
    Span4Mux_v I__1307 (
            .O(N__6944),
            .I(N__6941));
    Sp12to4 I__1306 (
            .O(N__6941),
            .I(N__6938));
    Odrv12 I__1305 (
            .O(N__6938),
            .I(un1_D_UU_AMIGA_7));
    InMux I__1304 (
            .O(N__6935),
            .I(N__6932));
    LocalMux I__1303 (
            .O(N__6932),
            .I(N__6929));
    Odrv12 I__1302 (
            .O(N__6929),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    InMux I__1301 (
            .O(N__6926),
            .I(N__6922));
    InMux I__1300 (
            .O(N__6925),
            .I(N__6919));
    LocalMux I__1299 (
            .O(N__6922),
            .I(N__6915));
    LocalMux I__1298 (
            .O(N__6919),
            .I(N__6912));
    InMux I__1297 (
            .O(N__6918),
            .I(N__6909));
    Span4Mux_v I__1296 (
            .O(N__6915),
            .I(N__6906));
    Span4Mux_v I__1295 (
            .O(N__6912),
            .I(N__6903));
    LocalMux I__1294 (
            .O(N__6909),
            .I(N__6898));
    Sp12to4 I__1293 (
            .O(N__6906),
            .I(N__6898));
    Sp12to4 I__1292 (
            .O(N__6903),
            .I(N__6895));
    Span12Mux_h I__1291 (
            .O(N__6898),
            .I(N__6892));
    Span12Mux_h I__1290 (
            .O(N__6895),
            .I(N__6889));
    Odrv12 I__1289 (
            .O(N__6892),
            .I(D_UU_AMIGA_in_2));
    Odrv12 I__1288 (
            .O(N__6889),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1287 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1286 (
            .O(N__6881),
            .I(N__6878));
    Span4Mux_s0_v I__1285 (
            .O(N__6878),
            .I(N__6875));
    Sp12to4 I__1284 (
            .O(N__6875),
            .I(N__6872));
    Span12Mux_h I__1283 (
            .O(N__6872),
            .I(N__6869));
    Odrv12 I__1282 (
            .O(N__6869),
            .I(un1_D_UU_AMIGA_2));
    CascadeMux I__1281 (
            .O(N__6866),
            .I(N__6863));
    InMux I__1280 (
            .O(N__6863),
            .I(N__6860));
    LocalMux I__1279 (
            .O(N__6860),
            .I(N__6857));
    Span4Mux_v I__1278 (
            .O(N__6857),
            .I(N__6854));
    Odrv4 I__1277 (
            .O(N__6854),
            .I(\U111_CYCLE_SM.FLIP_WORD_2 ));
    InMux I__1276 (
            .O(N__6851),
            .I(N__6843));
    InMux I__1275 (
            .O(N__6850),
            .I(N__6840));
    InMux I__1274 (
            .O(N__6849),
            .I(N__6837));
    InMux I__1273 (
            .O(N__6848),
            .I(N__6834));
    InMux I__1272 (
            .O(N__6847),
            .I(N__6829));
    InMux I__1271 (
            .O(N__6846),
            .I(N__6829));
    LocalMux I__1270 (
            .O(N__6843),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1269 (
            .O(N__6840),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1268 (
            .O(N__6837),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1267 (
            .O(N__6834),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1266 (
            .O(N__6829),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    InMux I__1265 (
            .O(N__6818),
            .I(N__6815));
    LocalMux I__1264 (
            .O(N__6815),
            .I(\U111_CYCLE_SM.N_160 ));
    InMux I__1263 (
            .O(N__6812),
            .I(N__6806));
    InMux I__1262 (
            .O(N__6811),
            .I(N__6806));
    LocalMux I__1261 (
            .O(N__6806),
            .I(N__6803));
    Span12Mux_v I__1260 (
            .O(N__6803),
            .I(N__6799));
    InMux I__1259 (
            .O(N__6802),
            .I(N__6796));
    Odrv12 I__1258 (
            .O(N__6799),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__1257 (
            .O(N__6796),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    InMux I__1256 (
            .O(N__6791),
            .I(N__6787));
    InMux I__1255 (
            .O(N__6790),
            .I(N__6784));
    LocalMux I__1254 (
            .O(N__6787),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ));
    LocalMux I__1253 (
            .O(N__6784),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ));
    InMux I__1252 (
            .O(N__6779),
            .I(N__6775));
    InMux I__1251 (
            .O(N__6778),
            .I(N__6772));
    LocalMux I__1250 (
            .O(N__6775),
            .I(N__6768));
    LocalMux I__1249 (
            .O(N__6772),
            .I(N__6765));
    InMux I__1248 (
            .O(N__6771),
            .I(N__6762));
    Span4Mux_h I__1247 (
            .O(N__6768),
            .I(N__6759));
    Span4Mux_h I__1246 (
            .O(N__6765),
            .I(N__6754));
    LocalMux I__1245 (
            .O(N__6762),
            .I(N__6751));
    Span4Mux_h I__1244 (
            .O(N__6759),
            .I(N__6748));
    InMux I__1243 (
            .O(N__6758),
            .I(N__6743));
    InMux I__1242 (
            .O(N__6757),
            .I(N__6743));
    Odrv4 I__1241 (
            .O(N__6754),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv4 I__1240 (
            .O(N__6751),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv4 I__1239 (
            .O(N__6748),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1238 (
            .O(N__6743),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1237 (
            .O(N__6734),
            .I(N__6727));
    InMux I__1236 (
            .O(N__6733),
            .I(N__6727));
    InMux I__1235 (
            .O(N__6732),
            .I(N__6724));
    LocalMux I__1234 (
            .O(N__6727),
            .I(N__6720));
    LocalMux I__1233 (
            .O(N__6724),
            .I(N__6714));
    InMux I__1232 (
            .O(N__6723),
            .I(N__6711));
    Span4Mux_v I__1231 (
            .O(N__6720),
            .I(N__6706));
    InMux I__1230 (
            .O(N__6719),
            .I(N__6703));
    InMux I__1229 (
            .O(N__6718),
            .I(N__6700));
    InMux I__1228 (
            .O(N__6717),
            .I(N__6697));
    Span4Mux_v I__1227 (
            .O(N__6714),
            .I(N__6692));
    LocalMux I__1226 (
            .O(N__6711),
            .I(N__6692));
    InMux I__1225 (
            .O(N__6710),
            .I(N__6689));
    InMux I__1224 (
            .O(N__6709),
            .I(N__6686));
    Sp12to4 I__1223 (
            .O(N__6706),
            .I(N__6675));
    LocalMux I__1222 (
            .O(N__6703),
            .I(N__6675));
    LocalMux I__1221 (
            .O(N__6700),
            .I(N__6675));
    LocalMux I__1220 (
            .O(N__6697),
            .I(N__6675));
    Sp12to4 I__1219 (
            .O(N__6692),
            .I(N__6675));
    LocalMux I__1218 (
            .O(N__6689),
            .I(N__6672));
    LocalMux I__1217 (
            .O(N__6686),
            .I(N__6669));
    Span12Mux_v I__1216 (
            .O(N__6675),
            .I(N__6666));
    Span12Mux_h I__1215 (
            .O(N__6672),
            .I(N__6661));
    Span12Mux_s7_h I__1214 (
            .O(N__6669),
            .I(N__6661));
    Span12Mux_h I__1213 (
            .O(N__6666),
            .I(N__6658));
    Span12Mux_v I__1212 (
            .O(N__6661),
            .I(N__6655));
    Odrv12 I__1211 (
            .O(N__6658),
            .I(RESETn_c));
    Odrv12 I__1210 (
            .O(N__6655),
            .I(RESETn_c));
    CascadeMux I__1209 (
            .O(N__6650),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ));
    InMux I__1208 (
            .O(N__6647),
            .I(N__6640));
    InMux I__1207 (
            .O(N__6646),
            .I(N__6640));
    InMux I__1206 (
            .O(N__6645),
            .I(N__6637));
    LocalMux I__1205 (
            .O(N__6640),
            .I(N__6632));
    LocalMux I__1204 (
            .O(N__6637),
            .I(N__6629));
    InMux I__1203 (
            .O(N__6636),
            .I(N__6624));
    InMux I__1202 (
            .O(N__6635),
            .I(N__6624));
    Odrv4 I__1201 (
            .O(N__6632),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    Odrv12 I__1200 (
            .O(N__6629),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1199 (
            .O(N__6624),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    InMux I__1198 (
            .O(N__6617),
            .I(N__6614));
    LocalMux I__1197 (
            .O(N__6614),
            .I(N__6610));
    InMux I__1196 (
            .O(N__6613),
            .I(N__6607));
    Span4Mux_v I__1195 (
            .O(N__6610),
            .I(N__6604));
    LocalMux I__1194 (
            .O(N__6607),
            .I(N__6601));
    Sp12to4 I__1193 (
            .O(N__6604),
            .I(N__6597));
    Span4Mux_v I__1192 (
            .O(N__6601),
            .I(N__6594));
    InMux I__1191 (
            .O(N__6600),
            .I(N__6591));
    Span12Mux_h I__1190 (
            .O(N__6597),
            .I(N__6588));
    Sp12to4 I__1189 (
            .O(N__6594),
            .I(N__6583));
    LocalMux I__1188 (
            .O(N__6591),
            .I(N__6583));
    Span12Mux_v I__1187 (
            .O(N__6588),
            .I(N__6578));
    Span12Mux_h I__1186 (
            .O(N__6583),
            .I(N__6578));
    Odrv12 I__1185 (
            .O(N__6578),
            .I(D_UM_AMIGA_in_1));
    InMux I__1184 (
            .O(N__6575),
            .I(N__6572));
    LocalMux I__1183 (
            .O(N__6572),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1182 (
            .O(N__6569),
            .I(N__6566));
    LocalMux I__1181 (
            .O(N__6566),
            .I(N__6563));
    IoSpan4Mux I__1180 (
            .O(N__6563),
            .I(N__6560));
    Span4Mux_s2_h I__1179 (
            .O(N__6560),
            .I(N__6557));
    Sp12to4 I__1178 (
            .O(N__6557),
            .I(N__6554));
    Span12Mux_h I__1177 (
            .O(N__6554),
            .I(N__6551));
    Odrv12 I__1176 (
            .O(N__6551),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1175 (
            .O(N__6548),
            .I(N__6545));
    LocalMux I__1174 (
            .O(N__6545),
            .I(N__6542));
    Glb2LocalMux I__1173 (
            .O(N__6542),
            .I(N__6539));
    GlobalMux I__1172 (
            .O(N__6539),
            .I(CLK80));
    IoInMux I__1171 (
            .O(N__6536),
            .I(N__6533));
    LocalMux I__1170 (
            .O(N__6533),
            .I(N__6530));
    IoSpan4Mux I__1169 (
            .O(N__6530),
            .I(N__6526));
    IoInMux I__1168 (
            .O(N__6529),
            .I(N__6523));
    Span4Mux_s3_v I__1167 (
            .O(N__6526),
            .I(N__6520));
    LocalMux I__1166 (
            .O(N__6523),
            .I(N__6517));
    Span4Mux_v I__1165 (
            .O(N__6520),
            .I(N__6514));
    IoSpan4Mux I__1164 (
            .O(N__6517),
            .I(N__6511));
    Span4Mux_v I__1163 (
            .O(N__6514),
            .I(N__6508));
    IoSpan4Mux I__1162 (
            .O(N__6511),
            .I(N__6505));
    Sp12to4 I__1161 (
            .O(N__6508),
            .I(N__6502));
    Span4Mux_s3_h I__1160 (
            .O(N__6505),
            .I(N__6499));
    Span12Mux_v I__1159 (
            .O(N__6502),
            .I(N__6494));
    Sp12to4 I__1158 (
            .O(N__6499),
            .I(N__6494));
    Odrv12 I__1157 (
            .O(N__6494),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1156 (
            .O(N__6491),
            .I(N__6488));
    LocalMux I__1155 (
            .O(N__6488),
            .I(N__6485));
    Span4Mux_v I__1154 (
            .O(N__6485),
            .I(N__6482));
    Sp12to4 I__1153 (
            .O(N__6482),
            .I(N__6479));
    Span12Mux_h I__1152 (
            .O(N__6479),
            .I(N__6476));
    Odrv12 I__1151 (
            .O(N__6476),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__1150 (
            .O(N__6473),
            .I(N__6470));
    LocalMux I__1149 (
            .O(N__6470),
            .I(N__6467));
    IoSpan4Mux I__1148 (
            .O(N__6467),
            .I(N__6464));
    Span4Mux_s3_h I__1147 (
            .O(N__6464),
            .I(N__6461));
    Span4Mux_h I__1146 (
            .O(N__6461),
            .I(N__6458));
    Sp12to4 I__1145 (
            .O(N__6458),
            .I(N__6455));
    Odrv12 I__1144 (
            .O(N__6455),
            .I(un2_D_LM_AMIGA_6));
    CascadeMux I__1143 (
            .O(N__6452),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ));
    InMux I__1142 (
            .O(N__6449),
            .I(N__6446));
    LocalMux I__1141 (
            .O(N__6446),
            .I(\U111_CYCLE_SM.N_149 ));
    InMux I__1140 (
            .O(N__6443),
            .I(N__6436));
    InMux I__1139 (
            .O(N__6442),
            .I(N__6433));
    InMux I__1138 (
            .O(N__6441),
            .I(N__6430));
    InMux I__1137 (
            .O(N__6440),
            .I(N__6425));
    InMux I__1136 (
            .O(N__6439),
            .I(N__6422));
    LocalMux I__1135 (
            .O(N__6436),
            .I(N__6417));
    LocalMux I__1134 (
            .O(N__6433),
            .I(N__6417));
    LocalMux I__1133 (
            .O(N__6430),
            .I(N__6414));
    InMux I__1132 (
            .O(N__6429),
            .I(N__6411));
    InMux I__1131 (
            .O(N__6428),
            .I(N__6408));
    LocalMux I__1130 (
            .O(N__6425),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1129 (
            .O(N__6422),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    Odrv4 I__1128 (
            .O(N__6417),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    Odrv4 I__1127 (
            .O(N__6414),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1126 (
            .O(N__6411),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1125 (
            .O(N__6408),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    InMux I__1124 (
            .O(N__6395),
            .I(N__6387));
    InMux I__1123 (
            .O(N__6394),
            .I(N__6384));
    InMux I__1122 (
            .O(N__6393),
            .I(N__6379));
    InMux I__1121 (
            .O(N__6392),
            .I(N__6379));
    InMux I__1120 (
            .O(N__6391),
            .I(N__6374));
    InMux I__1119 (
            .O(N__6390),
            .I(N__6374));
    LocalMux I__1118 (
            .O(N__6387),
            .I(N__6369));
    LocalMux I__1117 (
            .O(N__6384),
            .I(N__6369));
    LocalMux I__1116 (
            .O(N__6379),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1115 (
            .O(N__6374),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    Odrv4 I__1114 (
            .O(N__6369),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    CascadeMux I__1113 (
            .O(N__6362),
            .I(N__6359));
    InMux I__1112 (
            .O(N__6359),
            .I(N__6354));
    InMux I__1111 (
            .O(N__6358),
            .I(N__6351));
    InMux I__1110 (
            .O(N__6357),
            .I(N__6348));
    LocalMux I__1109 (
            .O(N__6354),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1108 (
            .O(N__6351),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1107 (
            .O(N__6348),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    CascadeMux I__1106 (
            .O(N__6341),
            .I(\U111_CYCLE_SM.N_132_0_cascade_ ));
    InMux I__1105 (
            .O(N__6338),
            .I(N__6334));
    InMux I__1104 (
            .O(N__6337),
            .I(N__6331));
    LocalMux I__1103 (
            .O(N__6334),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    LocalMux I__1102 (
            .O(N__6331),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    CascadeMux I__1101 (
            .O(N__6326),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_ ));
    CascadeMux I__1100 (
            .O(N__6323),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ));
    InMux I__1099 (
            .O(N__6320),
            .I(N__6317));
    LocalMux I__1098 (
            .O(N__6317),
            .I(N__6310));
    InMux I__1097 (
            .O(N__6316),
            .I(N__6307));
    InMux I__1096 (
            .O(N__6315),
            .I(N__6302));
    InMux I__1095 (
            .O(N__6314),
            .I(N__6302));
    InMux I__1094 (
            .O(N__6313),
            .I(N__6299));
    Span4Mux_v I__1093 (
            .O(N__6310),
            .I(N__6292));
    LocalMux I__1092 (
            .O(N__6307),
            .I(N__6292));
    LocalMux I__1091 (
            .O(N__6302),
            .I(N__6292));
    LocalMux I__1090 (
            .O(N__6299),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2 ));
    Odrv4 I__1089 (
            .O(N__6292),
            .I(\U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2 ));
    IoInMux I__1088 (
            .O(N__6287),
            .I(N__6282));
    InMux I__1087 (
            .O(N__6286),
            .I(N__6277));
    InMux I__1086 (
            .O(N__6285),
            .I(N__6277));
    LocalMux I__1085 (
            .O(N__6282),
            .I(N__6273));
    LocalMux I__1084 (
            .O(N__6277),
            .I(N__6270));
    InMux I__1083 (
            .O(N__6276),
            .I(N__6267));
    Span4Mux_s1_v I__1082 (
            .O(N__6273),
            .I(N__6262));
    Span4Mux_v I__1081 (
            .O(N__6270),
            .I(N__6257));
    LocalMux I__1080 (
            .O(N__6267),
            .I(N__6257));
    InMux I__1079 (
            .O(N__6266),
            .I(N__6254));
    InMux I__1078 (
            .O(N__6265),
            .I(N__6251));
    Span4Mux_v I__1077 (
            .O(N__6262),
            .I(N__6248));
    Span4Mux_v I__1076 (
            .O(N__6257),
            .I(N__6240));
    LocalMux I__1075 (
            .O(N__6254),
            .I(N__6240));
    LocalMux I__1074 (
            .O(N__6251),
            .I(N__6240));
    Sp12to4 I__1073 (
            .O(N__6248),
            .I(N__6237));
    InMux I__1072 (
            .O(N__6247),
            .I(N__6234));
    Span4Mux_v I__1071 (
            .O(N__6240),
            .I(N__6231));
    Span12Mux_h I__1070 (
            .O(N__6237),
            .I(N__6225));
    LocalMux I__1069 (
            .O(N__6234),
            .I(N__6225));
    Sp12to4 I__1068 (
            .O(N__6231),
            .I(N__6222));
    InMux I__1067 (
            .O(N__6230),
            .I(N__6219));
    Span12Mux_v I__1066 (
            .O(N__6225),
            .I(N__6212));
    Span12Mux_h I__1065 (
            .O(N__6222),
            .I(N__6212));
    LocalMux I__1064 (
            .O(N__6219),
            .I(N__6212));
    Span12Mux_v I__1063 (
            .O(N__6212),
            .I(N__6209));
    Odrv12 I__1062 (
            .O(N__6209),
            .I(TACKn_in));
    CascadeMux I__1061 (
            .O(N__6206),
            .I(N__6202));
    IoInMux I__1060 (
            .O(N__6205),
            .I(N__6198));
    InMux I__1059 (
            .O(N__6202),
            .I(N__6193));
    InMux I__1058 (
            .O(N__6201),
            .I(N__6193));
    LocalMux I__1057 (
            .O(N__6198),
            .I(N__6189));
    LocalMux I__1056 (
            .O(N__6193),
            .I(N__6186));
    InMux I__1055 (
            .O(N__6192),
            .I(N__6183));
    Span4Mux_s1_v I__1054 (
            .O(N__6189),
            .I(N__6179));
    Span4Mux_v I__1053 (
            .O(N__6186),
            .I(N__6174));
    LocalMux I__1052 (
            .O(N__6183),
            .I(N__6174));
    InMux I__1051 (
            .O(N__6182),
            .I(N__6171));
    Span4Mux_v I__1050 (
            .O(N__6179),
            .I(N__6168));
    Span4Mux_v I__1049 (
            .O(N__6174),
            .I(N__6162));
    LocalMux I__1048 (
            .O(N__6171),
            .I(N__6162));
    Sp12to4 I__1047 (
            .O(N__6168),
            .I(N__6158));
    InMux I__1046 (
            .O(N__6167),
            .I(N__6155));
    Span4Mux_v I__1045 (
            .O(N__6162),
            .I(N__6152));
    InMux I__1044 (
            .O(N__6161),
            .I(N__6149));
    Span12Mux_h I__1043 (
            .O(N__6158),
            .I(N__6146));
    LocalMux I__1042 (
            .O(N__6155),
            .I(N__6139));
    Sp12to4 I__1041 (
            .O(N__6152),
            .I(N__6139));
    LocalMux I__1040 (
            .O(N__6149),
            .I(N__6139));
    Span12Mux_v I__1039 (
            .O(N__6146),
            .I(N__6134));
    Span12Mux_h I__1038 (
            .O(N__6139),
            .I(N__6134));
    Span12Mux_v I__1037 (
            .O(N__6134),
            .I(N__6131));
    Odrv12 I__1036 (
            .O(N__6131),
            .I(TEAn_c));
    InMux I__1035 (
            .O(N__6128),
            .I(N__6125));
    LocalMux I__1034 (
            .O(N__6125),
            .I(N__6122));
    Odrv4 I__1033 (
            .O(N__6122),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ));
    CascadeMux I__1032 (
            .O(N__6119),
            .I(\U111_CYCLE_SM.N_160_cascade_ ));
    InMux I__1031 (
            .O(N__6116),
            .I(N__6110));
    InMux I__1030 (
            .O(N__6115),
            .I(N__6110));
    LocalMux I__1029 (
            .O(N__6110),
            .I(N__6107));
    Span4Mux_v I__1028 (
            .O(N__6107),
            .I(N__6104));
    Sp12to4 I__1027 (
            .O(N__6104),
            .I(N__6101));
    Span12Mux_h I__1026 (
            .O(N__6101),
            .I(N__6098));
    Span12Mux_v I__1025 (
            .O(N__6098),
            .I(N__6095));
    Odrv12 I__1024 (
            .O(N__6095),
            .I(SIZ_c_1));
    CascadeMux I__1023 (
            .O(N__6092),
            .I(N__6088));
    InMux I__1022 (
            .O(N__6091),
            .I(N__6083));
    InMux I__1021 (
            .O(N__6088),
            .I(N__6083));
    LocalMux I__1020 (
            .O(N__6083),
            .I(N__6080));
    Span4Mux_v I__1019 (
            .O(N__6080),
            .I(N__6077));
    Sp12to4 I__1018 (
            .O(N__6077),
            .I(N__6074));
    Span12Mux_h I__1017 (
            .O(N__6074),
            .I(N__6071));
    Span12Mux_v I__1016 (
            .O(N__6071),
            .I(N__6068));
    Odrv12 I__1015 (
            .O(N__6068),
            .I(SIZ_c_0));
    CascadeMux I__1014 (
            .O(N__6065),
            .I(\U111_CYCLE_SM.PORT_MISMATCH_2_cascade_ ));
    InMux I__1013 (
            .O(N__6062),
            .I(N__6057));
    InMux I__1012 (
            .O(N__6061),
            .I(N__6052));
    InMux I__1011 (
            .O(N__6060),
            .I(N__6049));
    LocalMux I__1010 (
            .O(N__6057),
            .I(N__6046));
    InMux I__1009 (
            .O(N__6056),
            .I(N__6043));
    InMux I__1008 (
            .O(N__6055),
            .I(N__6040));
    LocalMux I__1007 (
            .O(N__6052),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1006 (
            .O(N__6049),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    Odrv4 I__1005 (
            .O(N__6046),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1004 (
            .O(N__6043),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1003 (
            .O(N__6040),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    InMux I__1002 (
            .O(N__6029),
            .I(N__6026));
    LocalMux I__1001 (
            .O(N__6026),
            .I(\U111_CYCLE_SM.N_142_0 ));
    CascadeMux I__1000 (
            .O(N__6023),
            .I(N__6020));
    InMux I__999 (
            .O(N__6020),
            .I(N__6017));
    LocalMux I__998 (
            .O(N__6017),
            .I(N__6014));
    Span4Mux_h I__997 (
            .O(N__6014),
            .I(N__6011));
    Span4Mux_h I__996 (
            .O(N__6011),
            .I(N__6007));
    IoInMux I__995 (
            .O(N__6010),
            .I(N__6004));
    Sp12to4 I__994 (
            .O(N__6007),
            .I(N__6001));
    LocalMux I__993 (
            .O(N__6004),
            .I(N__5998));
    Span12Mux_v I__992 (
            .O(N__6001),
            .I(N__5995));
    IoSpan4Mux I__991 (
            .O(N__5998),
            .I(N__5992));
    Odrv12 I__990 (
            .O(N__5995),
            .I(TBIn_c));
    Odrv4 I__989 (
            .O(N__5992),
            .I(TBIn_c));
    InMux I__988 (
            .O(N__5987),
            .I(N__5983));
    InMux I__987 (
            .O(N__5986),
            .I(N__5980));
    LocalMux I__986 (
            .O(N__5983),
            .I(N__5976));
    LocalMux I__985 (
            .O(N__5980),
            .I(N__5973));
    InMux I__984 (
            .O(N__5979),
            .I(N__5970));
    Span4Mux_v I__983 (
            .O(N__5976),
            .I(N__5967));
    Span4Mux_v I__982 (
            .O(N__5973),
            .I(N__5962));
    LocalMux I__981 (
            .O(N__5970),
            .I(N__5962));
    Span4Mux_v I__980 (
            .O(N__5967),
            .I(N__5959));
    Span4Mux_v I__979 (
            .O(N__5962),
            .I(N__5956));
    Span4Mux_v I__978 (
            .O(N__5959),
            .I(N__5953));
    Span4Mux_h I__977 (
            .O(N__5956),
            .I(N__5950));
    Sp12to4 I__976 (
            .O(N__5953),
            .I(N__5945));
    Sp12to4 I__975 (
            .O(N__5950),
            .I(N__5945));
    Odrv12 I__974 (
            .O(N__5945),
            .I(D_UU_AMIGA_in_1));
    InMux I__973 (
            .O(N__5942),
            .I(N__5939));
    LocalMux I__972 (
            .O(N__5939),
            .I(N__5936));
    Odrv4 I__971 (
            .O(N__5936),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    IoInMux I__970 (
            .O(N__5933),
            .I(N__5930));
    LocalMux I__969 (
            .O(N__5930),
            .I(N__5927));
    Span4Mux_s2_h I__968 (
            .O(N__5927),
            .I(N__5924));
    Span4Mux_h I__967 (
            .O(N__5924),
            .I(N__5921));
    Sp12to4 I__966 (
            .O(N__5921),
            .I(N__5918));
    Span12Mux_s8_v I__965 (
            .O(N__5918),
            .I(N__5915));
    Odrv12 I__964 (
            .O(N__5915),
            .I(un1_D_UU_AMIGA_1));
    InMux I__963 (
            .O(N__5912),
            .I(N__5909));
    LocalMux I__962 (
            .O(N__5909),
            .I(N__5906));
    Span4Mux_v I__961 (
            .O(N__5906),
            .I(N__5903));
    Sp12to4 I__960 (
            .O(N__5903),
            .I(N__5900));
    Span12Mux_h I__959 (
            .O(N__5900),
            .I(N__5897));
    Odrv12 I__958 (
            .O(N__5897),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__957 (
            .O(N__5894),
            .I(N__5891));
    LocalMux I__956 (
            .O(N__5891),
            .I(N__5888));
    IoSpan4Mux I__955 (
            .O(N__5888),
            .I(N__5885));
    IoSpan4Mux I__954 (
            .O(N__5885),
            .I(N__5882));
    Span4Mux_s3_h I__953 (
            .O(N__5882),
            .I(N__5879));
    Sp12to4 I__952 (
            .O(N__5879),
            .I(N__5876));
    Odrv12 I__951 (
            .O(N__5876),
            .I(un2_D_LL_AMIGA_2));
    InMux I__950 (
            .O(N__5873),
            .I(N__5870));
    LocalMux I__949 (
            .O(N__5870),
            .I(N__5866));
    InMux I__948 (
            .O(N__5869),
            .I(N__5863));
    Odrv4 I__947 (
            .O(N__5866),
            .I(\U111_CYCLE_SM.TS_ENZ0Z6 ));
    LocalMux I__946 (
            .O(N__5863),
            .I(\U111_CYCLE_SM.TS_ENZ0Z6 ));
    CascadeMux I__945 (
            .O(N__5858),
            .I(\U111_CYCLE_SM.N_158_cascade_ ));
    InMux I__944 (
            .O(N__5855),
            .I(N__5852));
    LocalMux I__943 (
            .O(N__5852),
            .I(\U111_CYCLE_SM.N_130_0 ));
    CascadeMux I__942 (
            .O(N__5849),
            .I(N__5845));
    InMux I__941 (
            .O(N__5848),
            .I(N__5842));
    InMux I__940 (
            .O(N__5845),
            .I(N__5839));
    LocalMux I__939 (
            .O(N__5842),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    LocalMux I__938 (
            .O(N__5839),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    CascadeMux I__937 (
            .O(N__5834),
            .I(N__5831));
    InMux I__936 (
            .O(N__5831),
            .I(N__5828));
    LocalMux I__935 (
            .O(N__5828),
            .I(\U111_CYCLE_SM.TS_EN_6 ));
    InMux I__934 (
            .O(N__5825),
            .I(N__5822));
    LocalMux I__933 (
            .O(N__5822),
            .I(N__5819));
    Sp12to4 I__932 (
            .O(N__5819),
            .I(N__5815));
    InMux I__931 (
            .O(N__5818),
            .I(N__5812));
    Span12Mux_v I__930 (
            .O(N__5815),
            .I(N__5807));
    LocalMux I__929 (
            .O(N__5812),
            .I(N__5807));
    Span12Mux_h I__928 (
            .O(N__5807),
            .I(N__5804));
    Odrv12 I__927 (
            .O(N__5804),
            .I(A_040_c_1));
    IoInMux I__926 (
            .O(N__5801),
            .I(N__5798));
    LocalMux I__925 (
            .O(N__5798),
            .I(N__5795));
    Sp12to4 I__924 (
            .O(N__5795),
            .I(N__5792));
    Span12Mux_v I__923 (
            .O(N__5792),
            .I(N__5789));
    Odrv12 I__922 (
            .O(N__5789),
            .I(TSn_c));
    InMux I__921 (
            .O(N__5786),
            .I(N__5782));
    InMux I__920 (
            .O(N__5785),
            .I(N__5779));
    LocalMux I__919 (
            .O(N__5782),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__918 (
            .O(N__5779),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    CascadeMux I__917 (
            .O(N__5774),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ));
    CascadeMux I__916 (
            .O(N__5771),
            .I(\U111_CYCLE_SM.N_148_cascade_ ));
    CascadeMux I__915 (
            .O(N__5768),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ));
    InMux I__914 (
            .O(N__5765),
            .I(N__5762));
    LocalMux I__913 (
            .O(N__5762),
            .I(N__5759));
    Span4Mux_v I__912 (
            .O(N__5759),
            .I(N__5756));
    Span4Mux_h I__911 (
            .O(N__5756),
            .I(N__5753));
    Sp12to4 I__910 (
            .O(N__5753),
            .I(N__5750));
    Span12Mux_h I__909 (
            .O(N__5750),
            .I(N__5747));
    Odrv12 I__908 (
            .O(N__5747),
            .I(D_UU_040_in_5));
    IoInMux I__907 (
            .O(N__5744),
            .I(N__5741));
    LocalMux I__906 (
            .O(N__5741),
            .I(N__5738));
    IoSpan4Mux I__905 (
            .O(N__5738),
            .I(N__5734));
    InMux I__904 (
            .O(N__5737),
            .I(N__5731));
    IoSpan4Mux I__903 (
            .O(N__5734),
            .I(N__5728));
    LocalMux I__902 (
            .O(N__5731),
            .I(N__5725));
    Span4Mux_s2_h I__901 (
            .O(N__5728),
            .I(N__5722));
    Span4Mux_v I__900 (
            .O(N__5725),
            .I(N__5719));
    Sp12to4 I__899 (
            .O(N__5722),
            .I(N__5716));
    Sp12to4 I__898 (
            .O(N__5719),
            .I(N__5713));
    Span12Mux_h I__897 (
            .O(N__5716),
            .I(N__5710));
    Span12Mux_h I__896 (
            .O(N__5713),
            .I(N__5707));
    Span12Mux_h I__895 (
            .O(N__5710),
            .I(N__5702));
    Span12Mux_v I__894 (
            .O(N__5707),
            .I(N__5702));
    Odrv12 I__893 (
            .O(N__5702),
            .I(D_LM_040_in_5));
    IoInMux I__892 (
            .O(N__5699),
            .I(N__5696));
    LocalMux I__891 (
            .O(N__5696),
            .I(N__5693));
    Span4Mux_s2_h I__890 (
            .O(N__5693),
            .I(N__5690));
    Span4Mux_v I__889 (
            .O(N__5690),
            .I(N__5687));
    Sp12to4 I__888 (
            .O(N__5687),
            .I(N__5684));
    Odrv12 I__887 (
            .O(N__5684),
            .I(un1_D_UU_040_5));
    InMux I__886 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__885 (
            .O(N__5678),
            .I(N__5675));
    Span4Mux_v I__884 (
            .O(N__5675),
            .I(N__5672));
    Sp12to4 I__883 (
            .O(N__5672),
            .I(N__5669));
    Odrv12 I__882 (
            .O(N__5669),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__881 (
            .O(N__5666),
            .I(N__5663));
    LocalMux I__880 (
            .O(N__5663),
            .I(N__5660));
    Span4Mux_s2_h I__879 (
            .O(N__5660),
            .I(N__5657));
    Span4Mux_v I__878 (
            .O(N__5657),
            .I(N__5654));
    Span4Mux_v I__877 (
            .O(N__5654),
            .I(N__5651));
    Sp12to4 I__876 (
            .O(N__5651),
            .I(N__5648));
    Span12Mux_s11_h I__875 (
            .O(N__5648),
            .I(N__5645));
    Odrv12 I__874 (
            .O(N__5645),
            .I(un2_D_LL_AMIGA_6));
    InMux I__873 (
            .O(N__5642),
            .I(N__5639));
    LocalMux I__872 (
            .O(N__5639),
            .I(N__5636));
    Span4Mux_v I__871 (
            .O(N__5636),
            .I(N__5633));
    Sp12to4 I__870 (
            .O(N__5633),
            .I(N__5630));
    Span12Mux_h I__869 (
            .O(N__5630),
            .I(N__5627));
    Odrv12 I__868 (
            .O(N__5627),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__867 (
            .O(N__5624),
            .I(N__5621));
    LocalMux I__866 (
            .O(N__5621),
            .I(N__5618));
    IoSpan4Mux I__865 (
            .O(N__5618),
            .I(N__5615));
    Sp12to4 I__864 (
            .O(N__5615),
            .I(N__5612));
    Span12Mux_s7_h I__863 (
            .O(N__5612),
            .I(N__5609));
    Span12Mux_h I__862 (
            .O(N__5609),
            .I(N__5606));
    Odrv12 I__861 (
            .O(N__5606),
            .I(un2_D_LM_AMIGA_0));
    InMux I__860 (
            .O(N__5603),
            .I(N__5600));
    LocalMux I__859 (
            .O(N__5600),
            .I(N__5597));
    Span4Mux_v I__858 (
            .O(N__5597),
            .I(N__5594));
    Sp12to4 I__857 (
            .O(N__5594),
            .I(N__5591));
    Span12Mux_h I__856 (
            .O(N__5591),
            .I(N__5588));
    Odrv12 I__855 (
            .O(N__5588),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__854 (
            .O(N__5585),
            .I(N__5582));
    LocalMux I__853 (
            .O(N__5582),
            .I(N__5579));
    Span4Mux_s2_h I__852 (
            .O(N__5579),
            .I(N__5576));
    Span4Mux_v I__851 (
            .O(N__5576),
            .I(N__5573));
    Span4Mux_h I__850 (
            .O(N__5573),
            .I(N__5570));
    Sp12to4 I__849 (
            .O(N__5570),
            .I(N__5567));
    Span12Mux_h I__848 (
            .O(N__5567),
            .I(N__5564));
    Odrv12 I__847 (
            .O(N__5564),
            .I(un2_D_LL_AMIGA_3));
    InMux I__846 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__845 (
            .O(N__5558),
            .I(N__5555));
    Span4Mux_v I__844 (
            .O(N__5555),
            .I(N__5552));
    Sp12to4 I__843 (
            .O(N__5552),
            .I(N__5549));
    Span12Mux_h I__842 (
            .O(N__5549),
            .I(N__5546));
    Odrv12 I__841 (
            .O(N__5546),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__840 (
            .O(N__5543),
            .I(N__5540));
    LocalMux I__839 (
            .O(N__5540),
            .I(N__5537));
    Span12Mux_s6_h I__838 (
            .O(N__5537),
            .I(N__5534));
    Span12Mux_h I__837 (
            .O(N__5534),
            .I(N__5531));
    Odrv12 I__836 (
            .O(N__5531),
            .I(un2_D_LL_AMIGA_4));
    InMux I__835 (
            .O(N__5528),
            .I(N__5525));
    LocalMux I__834 (
            .O(N__5525),
            .I(N__5522));
    Span4Mux_v I__833 (
            .O(N__5522),
            .I(N__5519));
    Sp12to4 I__832 (
            .O(N__5519),
            .I(N__5516));
    Span12Mux_h I__831 (
            .O(N__5516),
            .I(N__5513));
    Odrv12 I__830 (
            .O(N__5513),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__829 (
            .O(N__5510),
            .I(N__5507));
    LocalMux I__828 (
            .O(N__5507),
            .I(N__5504));
    IoSpan4Mux I__827 (
            .O(N__5504),
            .I(N__5501));
    Span4Mux_s2_h I__826 (
            .O(N__5501),
            .I(N__5498));
    Span4Mux_h I__825 (
            .O(N__5498),
            .I(N__5495));
    Sp12to4 I__824 (
            .O(N__5495),
            .I(N__5492));
    Span12Mux_h I__823 (
            .O(N__5492),
            .I(N__5489));
    Odrv12 I__822 (
            .O(N__5489),
            .I(un2_D_LM_AMIGA_4));
    IoInMux I__821 (
            .O(N__5486),
            .I(N__5482));
    IoInMux I__820 (
            .O(N__5485),
            .I(N__5479));
    LocalMux I__819 (
            .O(N__5482),
            .I(N__5476));
    LocalMux I__818 (
            .O(N__5479),
            .I(N__5473));
    Span4Mux_s2_v I__817 (
            .O(N__5476),
            .I(N__5470));
    IoSpan4Mux I__816 (
            .O(N__5473),
            .I(N__5467));
    Span4Mux_h I__815 (
            .O(N__5470),
            .I(N__5464));
    Span4Mux_s2_v I__814 (
            .O(N__5467),
            .I(N__5461));
    Span4Mux_v I__813 (
            .O(N__5464),
            .I(N__5458));
    Span4Mux_v I__812 (
            .O(N__5461),
            .I(N__5455));
    Odrv4 I__811 (
            .O(N__5458),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__810 (
            .O(N__5455),
            .I(CONSTANT_ONE_NET));
    IoInMux I__809 (
            .O(N__5450),
            .I(N__5447));
    LocalMux I__808 (
            .O(N__5447),
            .I(N__5444));
    Odrv12 I__807 (
            .O(N__5444),
            .I(LBENn_c_i_0));
    InMux I__806 (
            .O(N__5441),
            .I(N__5438));
    LocalMux I__805 (
            .O(N__5438),
            .I(N__5435));
    Span4Mux_v I__804 (
            .O(N__5435),
            .I(N__5432));
    Sp12to4 I__803 (
            .O(N__5432),
            .I(N__5429));
    Span12Mux_h I__802 (
            .O(N__5429),
            .I(N__5426));
    Odrv12 I__801 (
            .O(N__5426),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__800 (
            .O(N__5423),
            .I(N__5420));
    LocalMux I__799 (
            .O(N__5420),
            .I(N__5417));
    IoSpan4Mux I__798 (
            .O(N__5417),
            .I(N__5414));
    IoSpan4Mux I__797 (
            .O(N__5414),
            .I(N__5411));
    Span4Mux_s2_h I__796 (
            .O(N__5411),
            .I(N__5408));
    Sp12to4 I__795 (
            .O(N__5408),
            .I(N__5405));
    Span12Mux_s9_h I__794 (
            .O(N__5405),
            .I(N__5402));
    Odrv12 I__793 (
            .O(N__5402),
            .I(un2_D_LL_AMIGA_1));
    IoInMux I__792 (
            .O(N__5399),
            .I(N__5396));
    LocalMux I__791 (
            .O(N__5396),
            .I(N__5393));
    Span4Mux_s1_h I__790 (
            .O(N__5393),
            .I(N__5390));
    Span4Mux_h I__789 (
            .O(N__5390),
            .I(N__5387));
    Span4Mux_h I__788 (
            .O(N__5387),
            .I(N__5384));
    Odrv4 I__787 (
            .O(N__5384),
            .I(un1_D_UU_040_1));
    InMux I__786 (
            .O(N__5381),
            .I(N__5378));
    LocalMux I__785 (
            .O(N__5378),
            .I(WRITE_CYCLE_ACTIVE_rep0_i_ess));
    IoInMux I__784 (
            .O(N__5375),
            .I(N__5372));
    LocalMux I__783 (
            .O(N__5372),
            .I(N__5369));
    IoSpan4Mux I__782 (
            .O(N__5369),
            .I(N__5366));
    Span4Mux_s3_v I__781 (
            .O(N__5366),
            .I(N__5363));
    Span4Mux_v I__780 (
            .O(N__5363),
            .I(N__5360));
    Odrv4 I__779 (
            .O(N__5360),
            .I(N_212_i));
    InMux I__778 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__777 (
            .O(N__5354),
            .I(WRITE_CYCLE_ACTIVE_rep4_i_ess));
    IoInMux I__776 (
            .O(N__5351),
            .I(N__5348));
    LocalMux I__775 (
            .O(N__5348),
            .I(N__5345));
    IoSpan4Mux I__774 (
            .O(N__5345),
            .I(N__5342));
    Span4Mux_s3_v I__773 (
            .O(N__5342),
            .I(N__5339));
    Odrv4 I__772 (
            .O(N__5339),
            .I(N_216_i));
    InMux I__771 (
            .O(N__5336),
            .I(N__5333));
    LocalMux I__770 (
            .O(N__5333),
            .I(WRITE_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__769 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__768 (
            .O(N__5327),
            .I(N__5324));
    Span12Mux_s7_v I__767 (
            .O(N__5324),
            .I(N__5321));
    Odrv12 I__766 (
            .O(N__5321),
            .I(N_225_i));
    IoInMux I__765 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__764 (
            .O(N__5315),
            .I(N__5312));
    IoSpan4Mux I__763 (
            .O(N__5312),
            .I(N__5309));
    Span4Mux_s2_v I__762 (
            .O(N__5309),
            .I(N__5306));
    Span4Mux_v I__761 (
            .O(N__5306),
            .I(N__5303));
    Odrv4 I__760 (
            .O(N__5303),
            .I(LBENn_c_i));
    InMux I__759 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__758 (
            .O(N__5297),
            .I(N__5294));
    Span4Mux_v I__757 (
            .O(N__5294),
            .I(N__5291));
    Span4Mux_h I__756 (
            .O(N__5291),
            .I(N__5288));
    Span4Mux_h I__755 (
            .O(N__5288),
            .I(N__5285));
    Odrv4 I__754 (
            .O(N__5285),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__753 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__752 (
            .O(N__5279),
            .I(N__5276));
    Span4Mux_s0_h I__751 (
            .O(N__5276),
            .I(N__5273));
    Sp12to4 I__750 (
            .O(N__5273),
            .I(N__5270));
    Span12Mux_s6_v I__749 (
            .O(N__5270),
            .I(N__5267));
    Span12Mux_h I__748 (
            .O(N__5267),
            .I(N__5264));
    Odrv12 I__747 (
            .O(N__5264),
            .I(un2_D_LL_AMIGA_0));
    InMux I__746 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__745 (
            .O(N__5258),
            .I(N__5255));
    Span12Mux_h I__744 (
            .O(N__5255),
            .I(N__5252));
    Odrv12 I__743 (
            .O(N__5252),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__742 (
            .O(N__5249),
            .I(N__5246));
    LocalMux I__741 (
            .O(N__5246),
            .I(N__5243));
    Span12Mux_s8_h I__740 (
            .O(N__5243),
            .I(N__5240));
    Span12Mux_v I__739 (
            .O(N__5240),
            .I(N__5237));
    Odrv12 I__738 (
            .O(N__5237),
            .I(un2_D_LM_AMIGA_2));
    InMux I__737 (
            .O(N__5234),
            .I(N__5231));
    LocalMux I__736 (
            .O(N__5231),
            .I(WRITE_CYCLE_ACTIVE_rep13_i_ess));
    IoInMux I__735 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__734 (
            .O(N__5225),
            .I(N__5222));
    IoSpan4Mux I__733 (
            .O(N__5222),
            .I(N__5219));
    Span4Mux_s2_h I__732 (
            .O(N__5219),
            .I(N__5216));
    Sp12to4 I__731 (
            .O(N__5216),
            .I(N__5213));
    Span12Mux_s11_h I__730 (
            .O(N__5213),
            .I(N__5210));
    Span12Mux_h I__729 (
            .O(N__5210),
            .I(N__5207));
    Odrv12 I__728 (
            .O(N__5207),
            .I(un2_D_LM_AMIGA_1));
    InMux I__727 (
            .O(N__5204),
            .I(N__5201));
    LocalMux I__726 (
            .O(N__5201),
            .I(N__5198));
    Odrv12 I__725 (
            .O(N__5198),
            .I(WRITE_CYCLE_ACTIVE_rep15_i_ess));
    InMux I__724 (
            .O(N__5195),
            .I(N__5192));
    LocalMux I__723 (
            .O(N__5192),
            .I(N__5189));
    Odrv12 I__722 (
            .O(N__5189),
            .I(WRITE_CYCLE_ACTIVE_rep3_i_ess));
    InMux I__721 (
            .O(N__5186),
            .I(N__5183));
    LocalMux I__720 (
            .O(N__5183),
            .I(N__5180));
    Odrv4 I__719 (
            .O(N__5180),
            .I(WRITE_CYCLE_ACTIVE_rep7_i_ess));
    InMux I__718 (
            .O(N__5177),
            .I(N__5174));
    LocalMux I__717 (
            .O(N__5174),
            .I(N__5171));
    Span12Mux_h I__716 (
            .O(N__5171),
            .I(N__5168));
    Odrv12 I__715 (
            .O(N__5168),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__714 (
            .O(N__5165),
            .I(N__5162));
    LocalMux I__713 (
            .O(N__5162),
            .I(N__5159));
    Span4Mux_s1_h I__712 (
            .O(N__5159),
            .I(N__5156));
    Span4Mux_h I__711 (
            .O(N__5156),
            .I(N__5153));
    Sp12to4 I__710 (
            .O(N__5153),
            .I(N__5150));
    Span12Mux_v I__709 (
            .O(N__5150),
            .I(N__5147));
    Span12Mux_h I__708 (
            .O(N__5147),
            .I(N__5144));
    Odrv12 I__707 (
            .O(N__5144),
            .I(un2_D_LM_AMIGA_3));
    InMux I__706 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__705 (
            .O(N__5138),
            .I(N__5135));
    Span4Mux_v I__704 (
            .O(N__5135),
            .I(N__5132));
    Sp12to4 I__703 (
            .O(N__5132),
            .I(N__5129));
    Odrv12 I__702 (
            .O(N__5129),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__701 (
            .O(N__5126),
            .I(N__5123));
    LocalMux I__700 (
            .O(N__5123),
            .I(N__5120));
    IoSpan4Mux I__699 (
            .O(N__5120),
            .I(N__5117));
    Span4Mux_s3_h I__698 (
            .O(N__5117),
            .I(N__5114));
    Span4Mux_v I__697 (
            .O(N__5114),
            .I(N__5111));
    Sp12to4 I__696 (
            .O(N__5111),
            .I(N__5108));
    Span12Mux_h I__695 (
            .O(N__5108),
            .I(N__5105));
    Odrv12 I__694 (
            .O(N__5105),
            .I(un2_D_LM_AMIGA_5));
    IoInMux I__693 (
            .O(N__5102),
            .I(N__5099));
    LocalMux I__692 (
            .O(N__5099),
            .I(N__5096));
    Span4Mux_s1_v I__691 (
            .O(N__5096),
            .I(N__5093));
    Span4Mux_h I__690 (
            .O(N__5093),
            .I(N__5090));
    Span4Mux_v I__689 (
            .O(N__5090),
            .I(N__5087));
    Odrv4 I__688 (
            .O(N__5087),
            .I(N_214_i));
    InMux I__687 (
            .O(N__5084),
            .I(N__5081));
    LocalMux I__686 (
            .O(N__5081),
            .I(N__5078));
    Span4Mux_v I__685 (
            .O(N__5078),
            .I(N__5075));
    Span4Mux_v I__684 (
            .O(N__5075),
            .I(N__5072));
    Sp12to4 I__683 (
            .O(N__5072),
            .I(N__5069));
    Span12Mux_h I__682 (
            .O(N__5069),
            .I(N__5066));
    Odrv12 I__681 (
            .O(N__5066),
            .I(D_UU_040_in_1));
    InMux I__680 (
            .O(N__5063),
            .I(N__5059));
    IoInMux I__679 (
            .O(N__5062),
            .I(N__5056));
    LocalMux I__678 (
            .O(N__5059),
            .I(N__5053));
    LocalMux I__677 (
            .O(N__5056),
            .I(N__5050));
    Span4Mux_v I__676 (
            .O(N__5053),
            .I(N__5047));
    Span4Mux_s3_h I__675 (
            .O(N__5050),
            .I(N__5044));
    Span4Mux_h I__674 (
            .O(N__5047),
            .I(N__5041));
    Sp12to4 I__673 (
            .O(N__5044),
            .I(N__5038));
    Span4Mux_v I__672 (
            .O(N__5041),
            .I(N__5035));
    Span12Mux_v I__671 (
            .O(N__5038),
            .I(N__5032));
    Sp12to4 I__670 (
            .O(N__5035),
            .I(N__5029));
    Span12Mux_h I__669 (
            .O(N__5032),
            .I(N__5026));
    Span12Mux_h I__668 (
            .O(N__5029),
            .I(N__5023));
    Span12Mux_h I__667 (
            .O(N__5026),
            .I(N__5018));
    Span12Mux_v I__666 (
            .O(N__5023),
            .I(N__5018));
    Odrv12 I__665 (
            .O(N__5018),
            .I(D_LM_040_in_1));
    InMux I__664 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__663 (
            .O(N__5012),
            .I(N__5009));
    Span4Mux_v I__662 (
            .O(N__5009),
            .I(N__5006));
    Span4Mux_h I__661 (
            .O(N__5006),
            .I(N__5003));
    Odrv4 I__660 (
            .O(N__5003),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__659 (
            .O(N__5000),
            .I(N__4997));
    LocalMux I__658 (
            .O(N__4997),
            .I(N__4994));
    Span12Mux_s9_h I__657 (
            .O(N__4994),
            .I(N__4991));
    Span12Mux_h I__656 (
            .O(N__4991),
            .I(N__4988));
    Odrv12 I__655 (
            .O(N__4988),
            .I(un2_D_LM_AMIGA_7));
    InMux I__654 (
            .O(N__4985),
            .I(N__4982));
    LocalMux I__653 (
            .O(N__4982),
            .I(N__4979));
    Span4Mux_v I__652 (
            .O(N__4979),
            .I(N__4976));
    Odrv4 I__651 (
            .O(N__4976),
            .I(WRITE_CYCLE_ACTIVE_rep12_i_ess));
    InMux I__650 (
            .O(N__4973),
            .I(N__4970));
    LocalMux I__649 (
            .O(N__4970),
            .I(N__4967));
    Odrv4 I__648 (
            .O(N__4967),
            .I(WRITE_CYCLE_ACTIVE_rep14_i_ess));
    InMux I__647 (
            .O(N__4964),
            .I(N__4961));
    LocalMux I__646 (
            .O(N__4961),
            .I(WRITE_CYCLE_ACTIVE_rep6_i_ess));
    IoInMux I__645 (
            .O(N__4958),
            .I(N__4955));
    LocalMux I__644 (
            .O(N__4955),
            .I(N__4952));
    IoSpan4Mux I__643 (
            .O(N__4952),
            .I(N__4949));
    Span4Mux_s2_v I__642 (
            .O(N__4949),
            .I(N__4946));
    Span4Mux_v I__641 (
            .O(N__4946),
            .I(N__4943));
    Odrv4 I__640 (
            .O(N__4943),
            .I(N_218_i));
    InMux I__639 (
            .O(N__4940),
            .I(N__4937));
    LocalMux I__638 (
            .O(N__4937),
            .I(N__4934));
    Span4Mux_v I__637 (
            .O(N__4934),
            .I(N__4931));
    Sp12to4 I__636 (
            .O(N__4931),
            .I(N__4928));
    Span12Mux_h I__635 (
            .O(N__4928),
            .I(N__4925));
    Span12Mux_h I__634 (
            .O(N__4925),
            .I(N__4922));
    Odrv12 I__633 (
            .O(N__4922),
            .I(D_UU_040_in_7));
    IoInMux I__632 (
            .O(N__4919),
            .I(N__4916));
    LocalMux I__631 (
            .O(N__4916),
            .I(N__4913));
    IoSpan4Mux I__630 (
            .O(N__4913),
            .I(N__4909));
    InMux I__629 (
            .O(N__4912),
            .I(N__4906));
    Span4Mux_s2_h I__628 (
            .O(N__4909),
            .I(N__4903));
    LocalMux I__627 (
            .O(N__4906),
            .I(N__4900));
    Span4Mux_h I__626 (
            .O(N__4903),
            .I(N__4895));
    Span4Mux_v I__625 (
            .O(N__4900),
            .I(N__4895));
    Span4Mux_h I__624 (
            .O(N__4895),
            .I(N__4892));
    Sp12to4 I__623 (
            .O(N__4892),
            .I(N__4889));
    Span12Mux_h I__622 (
            .O(N__4889),
            .I(N__4886));
    Odrv12 I__621 (
            .O(N__4886),
            .I(D_LM_040_in_7));
    IoInMux I__620 (
            .O(N__4883),
            .I(N__4880));
    LocalMux I__619 (
            .O(N__4880),
            .I(N__4877));
    IoSpan4Mux I__618 (
            .O(N__4877),
            .I(N__4874));
    Span4Mux_s2_v I__617 (
            .O(N__4874),
            .I(N__4871));
    Span4Mux_v I__616 (
            .O(N__4871),
            .I(N__4868));
    Odrv4 I__615 (
            .O(N__4868),
            .I(un1_D_UU_040_7));
    IoInMux I__614 (
            .O(N__4865),
            .I(N__4862));
    LocalMux I__613 (
            .O(N__4862),
            .I(N__4859));
    Span4Mux_s3_v I__612 (
            .O(N__4859),
            .I(N__4856));
    Span4Mux_h I__611 (
            .O(N__4856),
            .I(N__4853));
    Odrv4 I__610 (
            .O(N__4853),
            .I(N_219_i));
    InMux I__609 (
            .O(N__4850),
            .I(N__4847));
    LocalMux I__608 (
            .O(N__4847),
            .I(N__4844));
    Span4Mux_v I__607 (
            .O(N__4844),
            .I(N__4841));
    Sp12to4 I__606 (
            .O(N__4841),
            .I(N__4838));
    Odrv12 I__605 (
            .O(N__4838),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__604 (
            .O(N__4835),
            .I(N__4832));
    LocalMux I__603 (
            .O(N__4832),
            .I(N__4829));
    Span4Mux_s1_h I__602 (
            .O(N__4829),
            .I(N__4826));
    Span4Mux_h I__601 (
            .O(N__4826),
            .I(N__4823));
    Sp12to4 I__600 (
            .O(N__4823),
            .I(N__4820));
    Span12Mux_s11_v I__599 (
            .O(N__4820),
            .I(N__4817));
    Span12Mux_h I__598 (
            .O(N__4817),
            .I(N__4814));
    Odrv12 I__597 (
            .O(N__4814),
            .I(un2_D_LL_AMIGA_5));
    InMux I__596 (
            .O(N__4811),
            .I(N__4808));
    LocalMux I__595 (
            .O(N__4808),
            .I(N__4805));
    Odrv12 I__594 (
            .O(N__4805),
            .I(D_LM_AMIGA_in_1));
    InMux I__593 (
            .O(N__4802),
            .I(N__4799));
    LocalMux I__592 (
            .O(N__4799),
            .I(WRITE_CYCLE_ACTIVE_rep1_i_ess));
    InMux I__591 (
            .O(N__4796),
            .I(N__4793));
    LocalMux I__590 (
            .O(N__4793),
            .I(WRITE_CYCLE_ACTIVE_rep5_i_ess));
    IoInMux I__589 (
            .O(N__4790),
            .I(N__4787));
    LocalMux I__588 (
            .O(N__4787),
            .I(N__4784));
    Span4Mux_s3_v I__587 (
            .O(N__4784),
            .I(N__4781));
    Span4Mux_h I__586 (
            .O(N__4781),
            .I(N__4778));
    Odrv4 I__585 (
            .O(N__4778),
            .I(N_215_i));
    IoInMux I__584 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__583 (
            .O(N__4772),
            .I(N__4769));
    Odrv12 I__582 (
            .O(N__4769),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__581 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__580 (
            .O(N__4763),
            .I(N__4760));
    Span4Mux_h I__579 (
            .O(N__4760),
            .I(N__4757));
    Span4Mux_v I__578 (
            .O(N__4757),
            .I(N__4754));
    Odrv4 I__577 (
            .O(N__4754),
            .I(A_040_c_0));
    IoInMux I__576 (
            .O(N__4751),
            .I(N__4748));
    LocalMux I__575 (
            .O(N__4748),
            .I(N__4745));
    IoSpan4Mux I__574 (
            .O(N__4745),
            .I(N__4742));
    Span4Mux_s2_v I__573 (
            .O(N__4742),
            .I(N__4739));
    Span4Mux_v I__572 (
            .O(N__4739),
            .I(N__4736));
    Odrv4 I__571 (
            .O(N__4736),
            .I(A_AMIGA_c_0));
    InMux I__570 (
            .O(N__4733),
            .I(N__4730));
    LocalMux I__569 (
            .O(N__4730),
            .I(N__4727));
    Span4Mux_v I__568 (
            .O(N__4727),
            .I(N__4724));
    Span4Mux_h I__567 (
            .O(N__4724),
            .I(N__4721));
    Odrv4 I__566 (
            .O(N__4721),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__565 (
            .O(N__4718),
            .I(N__4715));
    LocalMux I__564 (
            .O(N__4715),
            .I(N__4712));
    Span4Mux_s2_h I__563 (
            .O(N__4712),
            .I(N__4709));
    Span4Mux_v I__562 (
            .O(N__4709),
            .I(N__4706));
    Sp12to4 I__561 (
            .O(N__4706),
            .I(N__4703));
    Span12Mux_h I__560 (
            .O(N__4703),
            .I(N__4700));
    Span12Mux_h I__559 (
            .O(N__4700),
            .I(N__4697));
    Odrv12 I__558 (
            .O(N__4697),
            .I(un2_D_LL_AMIGA_7));
    InMux I__557 (
            .O(N__4694),
            .I(N__4690));
    IoInMux I__556 (
            .O(N__4693),
            .I(N__4687));
    LocalMux I__555 (
            .O(N__4690),
            .I(N__4684));
    LocalMux I__554 (
            .O(N__4687),
            .I(N__4681));
    Span4Mux_v I__553 (
            .O(N__4684),
            .I(N__4678));
    IoSpan4Mux I__552 (
            .O(N__4681),
            .I(N__4675));
    Sp12to4 I__551 (
            .O(N__4678),
            .I(N__4672));
    Span4Mux_s2_h I__550 (
            .O(N__4675),
            .I(N__4669));
    Span12Mux_h I__549 (
            .O(N__4672),
            .I(N__4666));
    Sp12to4 I__548 (
            .O(N__4669),
            .I(N__4663));
    Span12Mux_v I__547 (
            .O(N__4666),
            .I(N__4660));
    Span12Mux_h I__546 (
            .O(N__4663),
            .I(N__4657));
    Span12Mux_h I__545 (
            .O(N__4660),
            .I(N__4654));
    Span12Mux_h I__544 (
            .O(N__4657),
            .I(N__4651));
    Odrv12 I__543 (
            .O(N__4654),
            .I(D_LL_040_in_2));
    Odrv12 I__542 (
            .O(N__4651),
            .I(D_LL_040_in_2));
    InMux I__541 (
            .O(N__4646),
            .I(N__4643));
    LocalMux I__540 (
            .O(N__4643),
            .I(N__4640));
    Span12Mux_h I__539 (
            .O(N__4640),
            .I(N__4637));
    Span12Mux_h I__538 (
            .O(N__4637),
            .I(N__4634));
    Odrv12 I__537 (
            .O(N__4634),
            .I(D_UM_040_in_2));
    IoInMux I__536 (
            .O(N__4631),
            .I(N__4628));
    LocalMux I__535 (
            .O(N__4628),
            .I(N__4625));
    Span4Mux_s1_h I__534 (
            .O(N__4625),
            .I(N__4622));
    Span4Mux_h I__533 (
            .O(N__4622),
            .I(N__4619));
    Span4Mux_v I__532 (
            .O(N__4619),
            .I(N__4616));
    Odrv4 I__531 (
            .O(N__4616),
            .I(un1_D_UM_040_2));
    InMux I__530 (
            .O(N__4613),
            .I(N__4610));
    LocalMux I__529 (
            .O(N__4610),
            .I(N__4607));
    Odrv4 I__528 (
            .O(N__4607),
            .I(WRITE_CYCLE_ACTIVE_rep8_i_ess));
    InMux I__527 (
            .O(N__4604),
            .I(N__4601));
    LocalMux I__526 (
            .O(N__4601),
            .I(N__4598));
    Odrv4 I__525 (
            .O(N__4598),
            .I(WRITE_CYCLE_ACTIVE_rep10_i_ess));
    InMux I__524 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__523 (
            .O(N__4592),
            .I(WRITE_CYCLE_ACTIVE_rep17_i_ess));
    InMux I__522 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__521 (
            .O(N__4586),
            .I(WRITE_CYCLE_ACTIVE_rep19_i_ess));
    InMux I__520 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__519 (
            .O(N__4580),
            .I(WRITE_CYCLE_ACTIVE_rep18_i_ess));
    InMux I__518 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__517 (
            .O(N__4574),
            .I(WRITE_CYCLE_ACTIVE_rep20_i_ess));
    InMux I__516 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__515 (
            .O(N__4568),
            .I(WRITE_CYCLE_ACTIVE_rep21_i_ess));
    InMux I__514 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__513 (
            .O(N__4562),
            .I(WRITE_CYCLE_ACTIVE_rep22_i_ess));
    InMux I__512 (
            .O(N__4559),
            .I(N__4556));
    LocalMux I__511 (
            .O(N__4556),
            .I(WRITE_CYCLE_ACTIVE_rep9_i_ess));
    InMux I__510 (
            .O(N__4553),
            .I(N__4550));
    LocalMux I__509 (
            .O(N__4550),
            .I(WRITE_CYCLE_ACTIVE_rep23_i_ess));
    InMux I__508 (
            .O(N__4547),
            .I(N__4544));
    LocalMux I__507 (
            .O(N__4544),
            .I(WRITE_CYCLE_ACTIVE_rep11_i_ess));
    InMux I__506 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__505 (
            .O(N__4538),
            .I(N__4535));
    Odrv4 I__504 (
            .O(N__4535),
            .I(WRITE_CYCLE_ACTIVE_rep24_i_ess));
    InMux I__503 (
            .O(N__4532),
            .I(N__4529));
    LocalMux I__502 (
            .O(N__4529),
            .I(WRITE_CYCLE_ACTIVE_rep25_i_ess));
    InMux I__501 (
            .O(N__4526),
            .I(N__4523));
    LocalMux I__500 (
            .O(N__4523),
            .I(WRITE_CYCLE_ACTIVE_rep28_i_ess));
    InMux I__499 (
            .O(N__4520),
            .I(N__4517));
    LocalMux I__498 (
            .O(N__4517),
            .I(N__4514));
    Odrv4 I__497 (
            .O(N__4514),
            .I(WRITE_CYCLE_ACTIVE_rep27_i_ess));
    InMux I__496 (
            .O(N__4511),
            .I(N__4508));
    LocalMux I__495 (
            .O(N__4508),
            .I(N__4505));
    Odrv12 I__494 (
            .O(N__4505),
            .I(WRITE_CYCLE_ACTIVE_rep26_i_ess));
    InMux I__493 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__492 (
            .O(N__4499),
            .I(WRITE_CYCLE_ACTIVE_rep30_i_ess));
    InMux I__491 (
            .O(N__4496),
            .I(N__4493));
    LocalMux I__490 (
            .O(N__4493),
            .I(WRITE_CYCLE_ACTIVE_rep16_i_ess));
    InMux I__489 (
            .O(N__4490),
            .I(N__4487));
    LocalMux I__488 (
            .O(N__4487),
            .I(WRITE_CYCLE_ACTIVE_rep29_i_ess));
    InMux I__487 (
            .O(N__4484),
            .I(N__4481));
    LocalMux I__486 (
            .O(N__4481),
            .I(WRITE_CYCLE_ACTIVE_i_ess));
    IoInMux I__485 (
            .O(N__4478),
            .I(N__4475));
    LocalMux I__484 (
            .O(N__4475),
            .I(N__4472));
    IoSpan4Mux I__483 (
            .O(N__4472),
            .I(N__4469));
    Span4Mux_s3_h I__482 (
            .O(N__4469),
            .I(N__4466));
    Odrv4 I__481 (
            .O(N__4466),
            .I(N_235_i));
    IoInMux I__480 (
            .O(N__4463),
            .I(N__4460));
    LocalMux I__479 (
            .O(N__4460),
            .I(N__4457));
    IoSpan4Mux I__478 (
            .O(N__4457),
            .I(N__4454));
    Span4Mux_s3_h I__477 (
            .O(N__4454),
            .I(N__4451));
    Odrv4 I__476 (
            .O(N__4451),
            .I(N_213_i));
    IoInMux I__475 (
            .O(N__4448),
            .I(N__4445));
    LocalMux I__474 (
            .O(N__4445),
            .I(N__4442));
    Span4Mux_s0_h I__473 (
            .O(N__4442),
            .I(N__4439));
    Span4Mux_h I__472 (
            .O(N__4439),
            .I(N__4436));
    Odrv4 I__471 (
            .O(N__4436),
            .I(N_223_i));
    IoInMux I__470 (
            .O(N__4433),
            .I(N__4430));
    LocalMux I__469 (
            .O(N__4430),
            .I(N__4427));
    IoSpan4Mux I__468 (
            .O(N__4427),
            .I(N__4424));
    Span4Mux_s3_h I__467 (
            .O(N__4424),
            .I(N__4421));
    Odrv4 I__466 (
            .O(N__4421),
            .I(N_224_i));
    IoInMux I__465 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__464 (
            .O(N__4415),
            .I(N__4412));
    IoSpan4Mux I__463 (
            .O(N__4412),
            .I(N__4409));
    Span4Mux_s3_v I__462 (
            .O(N__4409),
            .I(N__4406));
    Span4Mux_v I__461 (
            .O(N__4406),
            .I(N__4403));
    Odrv4 I__460 (
            .O(N__4403),
            .I(N_217_i));
    IoInMux I__459 (
            .O(N__4400),
            .I(N__4397));
    LocalMux I__458 (
            .O(N__4397),
            .I(N__4394));
    Span4Mux_s0_h I__457 (
            .O(N__4394),
            .I(N__4391));
    Span4Mux_h I__456 (
            .O(N__4391),
            .I(N__4388));
    Odrv4 I__455 (
            .O(N__4388),
            .I(N_227_i));
    IoInMux I__454 (
            .O(N__4385),
            .I(N__4382));
    LocalMux I__453 (
            .O(N__4382),
            .I(N__4379));
    IoSpan4Mux I__452 (
            .O(N__4379),
            .I(N__4376));
    Span4Mux_s0_h I__451 (
            .O(N__4376),
            .I(N__4373));
    Span4Mux_h I__450 (
            .O(N__4373),
            .I(N__4370));
    Odrv4 I__449 (
            .O(N__4370),
            .I(N_226_i));
    IoInMux I__448 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__447 (
            .O(N__4364),
            .I(N__4361));
    IoSpan4Mux I__446 (
            .O(N__4361),
            .I(N__4358));
    Span4Mux_s3_h I__445 (
            .O(N__4358),
            .I(N__4355));
    Odrv4 I__444 (
            .O(N__4355),
            .I(N_236_i));
    IoInMux I__443 (
            .O(N__4352),
            .I(N__4349));
    LocalMux I__442 (
            .O(N__4349),
            .I(N__4346));
    IoSpan4Mux I__441 (
            .O(N__4346),
            .I(N__4343));
    Span4Mux_s1_h I__440 (
            .O(N__4343),
            .I(N__4340));
    Span4Mux_h I__439 (
            .O(N__4340),
            .I(N__4337));
    Odrv4 I__438 (
            .O(N__4337),
            .I(N_239_i));
    IoInMux I__437 (
            .O(N__4334),
            .I(N__4331));
    LocalMux I__436 (
            .O(N__4331),
            .I(N__4328));
    IoSpan4Mux I__435 (
            .O(N__4328),
            .I(N__4325));
    Span4Mux_s1_h I__434 (
            .O(N__4325),
            .I(N__4322));
    Span4Mux_h I__433 (
            .O(N__4322),
            .I(N__4319));
    Odrv4 I__432 (
            .O(N__4319),
            .I(N_238_i));
    IoInMux I__431 (
            .O(N__4316),
            .I(N__4313));
    LocalMux I__430 (
            .O(N__4313),
            .I(N__4310));
    Odrv12 I__429 (
            .O(N__4310),
            .I(RESETn_c_i));
    IoInMux I__428 (
            .O(N__4307),
            .I(N__4304));
    LocalMux I__427 (
            .O(N__4304),
            .I(N__4301));
    Odrv12 I__426 (
            .O(N__4301),
            .I(N_231_i));
    IoInMux I__425 (
            .O(N__4298),
            .I(N__4295));
    LocalMux I__424 (
            .O(N__4295),
            .I(N__4292));
    Odrv12 I__423 (
            .O(N__4292),
            .I(N_220_i));
    IoInMux I__422 (
            .O(N__4289),
            .I(N__4286));
    LocalMux I__421 (
            .O(N__4286),
            .I(N__4283));
    Odrv12 I__420 (
            .O(N__4283),
            .I(N_230_i));
    IoInMux I__419 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__418 (
            .O(N__4277),
            .I(N__4274));
    Span12Mux_s4_h I__417 (
            .O(N__4274),
            .I(N__4271));
    Odrv12 I__416 (
            .O(N__4271),
            .I(N_232_i));
    IoInMux I__415 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__414 (
            .O(N__4265),
            .I(N__4262));
    IoSpan4Mux I__413 (
            .O(N__4262),
            .I(N__4259));
    Span4Mux_s3_h I__412 (
            .O(N__4259),
            .I(N__4256));
    Odrv4 I__411 (
            .O(N__4256),
            .I(N_222_i));
    IoInMux I__410 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__409 (
            .O(N__4250),
            .I(N__4247));
    IoSpan4Mux I__408 (
            .O(N__4247),
            .I(N__4244));
    Span4Mux_s3_h I__407 (
            .O(N__4244),
            .I(N__4241));
    Odrv4 I__406 (
            .O(N__4241),
            .I(N_221_i));
    IoInMux I__405 (
            .O(N__4238),
            .I(N__4235));
    LocalMux I__404 (
            .O(N__4235),
            .I(N__4232));
    IoSpan4Mux I__403 (
            .O(N__4232),
            .I(N__4229));
    Span4Mux_s2_h I__402 (
            .O(N__4229),
            .I(N__4226));
    Odrv4 I__401 (
            .O(N__4226),
            .I(N_233_i));
    IoInMux I__400 (
            .O(N__4223),
            .I(N__4220));
    LocalMux I__399 (
            .O(N__4220),
            .I(N__4217));
    IoSpan4Mux I__398 (
            .O(N__4217),
            .I(N__4214));
    Span4Mux_s3_h I__397 (
            .O(N__4214),
            .I(N__4211));
    Odrv4 I__396 (
            .O(N__4211),
            .I(N_234_i));
    IoInMux I__395 (
            .O(N__4208),
            .I(N__4205));
    LocalMux I__394 (
            .O(N__4205),
            .I(N__4202));
    Span4Mux_s0_v I__393 (
            .O(N__4202),
            .I(N__4199));
    Sp12to4 I__392 (
            .O(N__4199),
            .I(N__4196));
    Span12Mux_h I__391 (
            .O(N__4196),
            .I(N__4193));
    Span12Mux_v I__390 (
            .O(N__4193),
            .I(N__4190));
    Span12Mux_v I__389 (
            .O(N__4190),
            .I(N__4187));
    Odrv12 I__388 (
            .O(N__4187),
            .I(TAn_in));
    IoInMux I__387 (
            .O(N__4184),
            .I(N__4181));
    LocalMux I__386 (
            .O(N__4181),
            .I(N__4178));
    Span12Mux_s4_h I__385 (
            .O(N__4178),
            .I(N__4175));
    Odrv12 I__384 (
            .O(N__4175),
            .I(N_237_i));
    IoInMux I__383 (
            .O(N__4172),
            .I(N__4169));
    LocalMux I__382 (
            .O(N__4169),
            .I(N__4166));
    IoSpan4Mux I__381 (
            .O(N__4166),
            .I(N__4163));
    Span4Mux_s1_h I__380 (
            .O(N__4163),
            .I(N__4160));
    Odrv4 I__379 (
            .O(N__4160),
            .I(N_240_i));
    IoInMux I__378 (
            .O(N__4157),
            .I(N__4154));
    LocalMux I__377 (
            .O(N__4154),
            .I(N__4151));
    Span4Mux_s0_h I__376 (
            .O(N__4151),
            .I(N__4148));
    Span4Mux_h I__375 (
            .O(N__4148),
            .I(N__4145));
    Odrv4 I__374 (
            .O(N__4145),
            .I(N_242_i));
    IoInMux I__373 (
            .O(N__4142),
            .I(N__4139));
    LocalMux I__372 (
            .O(N__4139),
            .I(N__4136));
    Span4Mux_s0_h I__371 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_h I__370 (
            .O(N__4133),
            .I(N__4130));
    Odrv4 I__369 (
            .O(N__4130),
            .I(N_228_i));
    IoInMux I__368 (
            .O(N__4127),
            .I(N__4124));
    LocalMux I__367 (
            .O(N__4124),
            .I(N__4121));
    IoSpan4Mux I__366 (
            .O(N__4121),
            .I(N__4118));
    Span4Mux_s3_h I__365 (
            .O(N__4118),
            .I(N__4115));
    Odrv4 I__364 (
            .O(N__4115),
            .I(N_241_i));
    IoInMux I__363 (
            .O(N__4112),
            .I(N__4109));
    LocalMux I__362 (
            .O(N__4109),
            .I(N__4106));
    Span12Mux_s4_h I__361 (
            .O(N__4106),
            .I(N__4103));
    Odrv12 I__360 (
            .O(N__4103),
            .I(N_243_i));
    IoInMux I__359 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__358 (
            .O(N__4097),
            .I(N__4094));
    Span4Mux_s0_h I__357 (
            .O(N__4094),
            .I(N__4091));
    Span4Mux_h I__356 (
            .O(N__4091),
            .I(N__4088));
    Odrv4 I__355 (
            .O(N__4088),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_0 ));
    IoInMux I__354 (
            .O(N__4085),
            .I(N__4082));
    LocalMux I__353 (
            .O(N__4082),
            .I(N__4079));
    Odrv12 I__352 (
            .O(N__4079),
            .I(N_229_i));
    IoInMux I__351 (
            .O(N__4076),
            .I(N__4073));
    LocalMux I__350 (
            .O(N__4073),
            .I(N__4070));
    IoSpan4Mux I__349 (
            .O(N__4070),
            .I(N__4067));
    Span4Mux_s3_h I__348 (
            .O(N__4067),
            .I(N__4064));
    Sp12to4 I__347 (
            .O(N__4064),
            .I(N__4061));
    Span12Mux_s8_h I__346 (
            .O(N__4061),
            .I(N__4058));
    Span12Mux_v I__345 (
            .O(N__4058),
            .I(N__4055));
    Span12Mux_v I__344 (
            .O(N__4055),
            .I(N__4052));
    Span12Mux_h I__343 (
            .O(N__4052),
            .I(N__4049));
    Odrv12 I__342 (
            .O(N__4049),
            .I(TCIn_c));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__10601));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__4316),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4100),
            .GLOBALBUFFEROUTPUT(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_3_1.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_3_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_1_LC_1_3_1 (
            .in0(N__4532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_237_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_1_3_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_1_3_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_1_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_4_LC_1_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4526),
            .lcout(N_240_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4502),
            .lcout(N_242_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_4.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_4.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_0_LC_1_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(N_228_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_7_6.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_7_6.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_5_LC_1_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4490),
            .lcout(N_241_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_9_1.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_9_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_7_LC_1_9_1 (
            .in0(N__4484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_243_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_0  (
            .in0(N__10319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6779),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_10_5.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_1_LC_1_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4595),
            .lcout(N_229_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_10_6 (
            .in0(N__6709),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_1_11_5.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_1_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_3_LC_1_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4589),
            .lcout(N_231_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_1.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_0_LC_1_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4613),
            .lcout(N_220_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_1_12_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_1_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_2_LC_1_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4583),
            .lcout(N_230_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_4_LC_1_13_1 (
            .in0(N__4577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_232_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_6.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_2_LC_1_13_6 (
            .in0(N__4604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_222_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_0.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_0.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_1_LC_1_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4559),
            .lcout(N_221_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_7.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_7.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_5_LC_1_15_7 (
            .in0(N__4571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_233_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_16_0.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_16_0.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_16_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_6_LC_1_16_0 (
            .in0(N__4565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_234_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_7_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4553),
            .lcout(N_235_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_6.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_6.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_1_LC_1_18_6 (
            .in0(N__4802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_213_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_18_7.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_18_7.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_18_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_3_LC_1_18_7 (
            .in0(N__4547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_223_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_0.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_0.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_4_LC_1_19_0 (
            .in0(N__4985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_224_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_1_19_1.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_1_19_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_5_LC_1_19_1 (
            .in0(N__4796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_217_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_2.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_2.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_7_LC_1_19_2 (
            .in0(N__5204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_227_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_4.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_19_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_6_LC_1_19_4 (
            .in0(N__4973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_226_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_2_1_6.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_2_1_6.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_2_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_0_LC_2_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4541),
            .lcout(N_236_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_2_2_4.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_2_2_4.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_2_2_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_3_LC_2_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4520),
            .lcout(N_239_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_2_2_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_2_2_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_2_2_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_2_LC_2_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4511),
            .lcout(N_238_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_2_3_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_2_3_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_2_3_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_2_3_3  (
            .in0(N__12545),
            .in1(N__11117),
            .in2(N__12184),
            .in3(N__11231),
            .lcout(WRITE_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10625),
            .ce(N__10422),
            .sr(N__10283));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_3_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_3_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_3_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_3_4  (
            .in0(N__11232),
            .in1(N__11079),
            .in2(N__12185),
            .in3(N__12546),
            .lcout(WRITE_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10625),
            .ce(N__10422),
            .sr(N__10283));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_2_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_2_3_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_2_3_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_2_3_7  (
            .in0(N__12547),
            .in1(N__12183),
            .in2(N__11113),
            .in3(N__11233),
            .lcout(WRITE_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10625),
            .ce(N__10422),
            .sr(N__10283));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_2_4_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_2_4_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_2_4_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_2_4_2  (
            .in0(N__12168),
            .in1(N__11116),
            .in2(N__12722),
            .in3(N__11430),
            .lcout(WRITE_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10622),
            .ce(N__10419),
            .sr(N__10281));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_2_5_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_2_5_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_2_5_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_2_5_6  (
            .in0(N__11115),
            .in1(N__12167),
            .in2(N__11509),
            .in3(N__12713),
            .lcout(WRITE_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10621),
            .ce(N__10417),
            .sr(N__10279));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_6  (
            .in0(N__12166),
            .in1(N__11114),
            .in2(N__12721),
            .in3(N__11434),
            .lcout(WRITE_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10619),
            .ce(N__10416),
            .sr(N__10277));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_7_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_7_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_7_6  (
            .in0(N__11093),
            .in1(N__12165),
            .in2(N__11510),
            .in3(N__12717),
            .lcout(WRITE_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10617),
            .ce(N__10414),
            .sr(N__10274));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_2_8_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_2_8_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_2_8_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_2_8_0  (
            .in0(N__11092),
            .in1(N__12144),
            .in2(N__11564),
            .in3(N__12689),
            .lcout(WRITE_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10616),
            .ce(N__10412),
            .sr(N__10272));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_9_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_9_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_9_4  (
            .in0(N__11091),
            .in1(N__11514),
            .in2(N__12164),
            .in3(N__12679),
            .lcout(WRITE_CYCLE_ACTIVE_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10614),
            .ce(N__10409),
            .sr(N__10270));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_2_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_2_10_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_2_10_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_2_10_5  (
            .in0(N__11090),
            .in1(N__12678),
            .in2(N__12163),
            .in3(N__11515),
            .lcout(WRITE_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10610),
            .ce(N__10407),
            .sr(N__10269));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_2_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_2_11_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_2_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_2_11_5  (
            .in0(N__11033),
            .in1(N__12137),
            .in2(N__12720),
            .in3(N__11516),
            .lcout(WRITE_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10609),
            .ce(N__10406),
            .sr(N__10271));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_2_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_2_12_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_2_12_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_2_12_3  (
            .in0(N__11032),
            .in1(N__12620),
            .in2(N__11606),
            .in3(N__12106),
            .lcout(WRITE_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10607),
            .ce(N__10408),
            .sr(N__10273));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_0  (
            .in0(N__12099),
            .in1(N__11030),
            .in2(N__12677),
            .in3(N__11570),
            .lcout(WRITE_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10605),
            .ce(N__10410),
            .sr(N__10275));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_2_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_2_15_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_2_15_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_2_15_0  (
            .in0(N__11057),
            .in1(N__12096),
            .in2(N__12544),
            .in3(N__11571),
            .lcout(WRITE_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10603),
            .ce(N__10415),
            .sr(N__10280));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_15_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_15_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_15_2  (
            .in0(N__12467),
            .in1(N__12097),
            .in2(N__11106),
            .in3(N__11572),
            .lcout(WRITE_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10603),
            .ce(N__10415),
            .sr(N__10280));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_2_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_2_15_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_2_15_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_2_15_6  (
            .in0(N__12468),
            .in1(N__12098),
            .in2(N__11107),
            .in3(N__11573),
            .lcout(WRITE_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10603),
            .ce(N__10415),
            .sr(N__10280));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_2_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_2_17_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_2_17_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_2_17_5  (
            .in0(N__12640),
            .in1(N__11065),
            .in2(N__12095),
            .in3(N__11608),
            .lcout(WRITE_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10600),
            .ce(N__10418),
            .sr(N__10282));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_18_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_18_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_18_1  (
            .in0(N__11108),
            .in1(N__12641),
            .in2(N__11629),
            .in3(N__12034),
            .lcout(WRITE_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10595),
            .ce(N__10420),
            .sr(N__10284));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_3  (
            .in0(N__11109),
            .in1(N__12642),
            .in2(N__11630),
            .in3(N__12035),
            .lcout(WRITE_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10595),
            .ce(N__10420),
            .sr(N__10284));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_19_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_19_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_19_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_19_6  (
            .in0(N__11112),
            .in1(N__12033),
            .in2(N__12695),
            .in3(N__11617),
            .lcout(WRITE_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10588),
            .ce(N__10421),
            .sr(N__10285));
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_6.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_6.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_3_LC_2_20_6 (
            .in0(N__5195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_215_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_2  (
            .in0(_gnd_net_),
            .in1(N__5818),
            .in2(_gnd_net_),
            .in3(N__6812),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_4  (
            .in0(N__4766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6811),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_3_7_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_3_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_3_7_0  (
            .in0(N__8958),
            .in1(N__7145),
            .in2(_gnd_net_),
            .in3(N__4733),
            .lcout(un2_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_3_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_3_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_3_10_1  (
            .in0(N__8959),
            .in1(N__4694),
            .in2(_gnd_net_),
            .in3(N__4646),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_3_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_3_12_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_3_12_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_3_12_1  (
            .in0(N__11565),
            .in1(N__11031),
            .in2(N__12136),
            .in3(N__12670),
            .lcout(WRITE_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10606),
            .ce(N__10411),
            .sr(N__10276));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_3_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_3_13_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_3_13_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_3_13_1  (
            .in0(N__11566),
            .in1(N__11029),
            .in2(N__12019),
            .in3(N__12669),
            .lcout(WRITE_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10604),
            .ce(N__10413),
            .sr(N__10278));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_3_17_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_3_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_3_17_4  (
            .in0(N__5015),
            .in1(N__6993),
            .in2(_gnd_net_),
            .in3(N__8963),
            .lcout(un2_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_3_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_3_18_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_3_18_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_3_18_2  (
            .in0(N__11064),
            .in1(N__11607),
            .in2(N__12709),
            .in3(N__12032),
            .lcout(WRITE_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10589),
            .ce(N__10423),
            .sr(N__10286));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_3_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_3_19_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_3_19_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_3_19_5  (
            .in0(N__11958),
            .in1(N__11111),
            .in2(N__12694),
            .in3(N__11616),
            .lcout(WRITE_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10584),
            .ce(N__10424),
            .sr(N__10288));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_3_19_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_3_19_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_3_19_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_3_19_7  (
            .in0(N__11957),
            .in1(N__11110),
            .in2(N__12693),
            .in3(N__11615),
            .lcout(WRITE_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10584),
            .ce(N__10424),
            .sr(N__10288));
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_0.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_0.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_6_LC_3_20_0 (
            .in0(N__4964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_218_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_3_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_3_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_3_20_1  (
            .in0(N__8964),
            .in1(N__4940),
            .in2(_gnd_net_),
            .in3(N__4912),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_20_6.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_20_6.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_20_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_7_LC_3_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5186),
            .lcout(N_219_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_2  (
            .in0(N__4850),
            .in1(N__7214),
            .in2(_gnd_net_),
            .in3(N__8980),
            .lcout(un2_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_0  (
            .in0(N__9007),
            .in1(N__5987),
            .in2(_gnd_net_),
            .in3(N__4811),
            .lcout(un2_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_19_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_19_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_19_1  (
            .in0(N__11619),
            .in1(N__11085),
            .in2(N__11990),
            .in3(N__12603),
            .lcout(WRITE_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10579),
            .ce(N__10425),
            .sr(N__10294));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_5_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_5_19_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_5_19_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_5_19_5  (
            .in0(N__11620),
            .in1(N__11086),
            .in2(N__11991),
            .in3(N__12604),
            .lcout(WRITE_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10579),
            .ce(N__10425),
            .sr(N__10294));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_5_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_5_20_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_5_20_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_5_20_1  (
            .in0(N__12699),
            .in1(N__11087),
            .in2(N__11988),
            .in3(N__11631),
            .lcout(WRITE_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10575),
            .ce(N__10427),
            .sr(N__10297));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_5_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_5_20_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_5_20_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_5_20_6  (
            .in0(N__11089),
            .in1(N__11633),
            .in2(N__12719),
            .in3(N__11905),
            .lcout(WRITE_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10575),
            .ce(N__10427),
            .sr(N__10297));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_7  (
            .in0(N__12700),
            .in1(N__11088),
            .in2(N__11989),
            .in3(N__11632),
            .lcout(WRITE_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10575),
            .ce(N__10427),
            .sr(N__10297));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_11_3  (
            .in0(N__5177),
            .in1(N__7783),
            .in2(_gnd_net_),
            .in3(N__8973),
            .lcout(un2_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_15_7  (
            .in0(N__5141),
            .in1(N__8602),
            .in2(_gnd_net_),
            .in3(N__9005),
            .lcout(un2_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_6_18_3.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_6_18_3.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_6_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_2_LC_6_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5336),
            .lcout(N_214_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_6_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_6_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_6_18_5  (
            .in0(N__9020),
            .in1(N__5084),
            .in2(_gnd_net_),
            .in3(N__5063),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_6_19_2.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_6_19_2.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_6_19_2.LUT_INIT=16'b0011001100110011;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_0_LC_6_19_2 (
            .in0(_gnd_net_),
            .in1(N__5381),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_212_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_4.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_4.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_4_LC_6_20_4 (
            .in0(N__5357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_216_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_18_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_18_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_18_5  (
            .in0(N__11505),
            .in1(N__11016),
            .in2(N__12031),
            .in3(N__12528),
            .lcout(WRITE_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10573),
            .ce(N__10426),
            .sr(N__10295));
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_7_19_2.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_7_19_2.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_7_19_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_5_LC_7_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5234),
            .lcout(N_225_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BUFENn_obuf_RNO_LC_7_20_1.C_ON=1'b0;
    defparam BUFENn_obuf_RNO_LC_7_20_1.SEQ_MODE=4'b0000;
    defparam BUFENn_obuf_RNO_LC_7_20_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 BUFENn_obuf_RNO_LC_7_20_1 (
            .in0(N__11563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_1_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_1_0  (
            .in0(N__9004),
            .in1(N__5300),
            .in2(_gnd_net_),
            .in3(N__7289),
            .lcout(un2_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_4  (
            .in0(N__8969),
            .in1(N__6926),
            .in2(_gnd_net_),
            .in3(N__5261),
            .lcout(un2_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_8_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_8_19_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_8_19_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_8_19_2  (
            .in0(N__11015),
            .in1(N__11875),
            .in2(N__11618),
            .in3(N__12452),
            .lcout(WRITE_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(N__10428),
            .sr(N__10298));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_8_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_8_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_8_20_7  (
            .in0(N__5765),
            .in1(N__5737),
            .in2(_gnd_net_),
            .in3(N__9003),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_9_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_9_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_9_6_0  (
            .in0(N__7403),
            .in1(N__5681),
            .in2(_gnd_net_),
            .in3(N__8919),
            .lcout(un2_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_5  (
            .in0(N__8890),
            .in1(N__7073),
            .in2(_gnd_net_),
            .in3(N__5642),
            .lcout(un2_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_1  (
            .in0(N__5603),
            .in1(N__7702),
            .in2(_gnd_net_),
            .in3(N__8979),
            .lcout(un2_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_10_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_10_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_10_3_5  (
            .in0(N__7636),
            .in1(N__5561),
            .in2(_gnd_net_),
            .in3(N__8965),
            .lcout(un2_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_10_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_10_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_10_13_1  (
            .in0(N__5528),
            .in1(N__8552),
            .in2(_gnd_net_),
            .in3(N__8993),
            .lcout(un2_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_20_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_20_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_1.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_1 (
            .in0(N__11216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_11_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_11_3_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_11_3_0  (
            .in0(N__8935),
            .in1(N__5441),
            .in2(_gnd_net_),
            .in3(N__6617),
            .lcout(un2_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_6  (
            .in0(N__7504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5825),
            .lcout(\U111_CYCLE_SM.FLIP_WORD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_11_7_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_11_7_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_11_7_7  (
            .in0(N__6723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5785),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_11_8_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_8_2 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_11_8_2  (
            .in0(N__5786),
            .in1(N__6791),
            .in2(N__5834),
            .in3(N__5855),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10596),
            .ce(),
            .sr(N__10289));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_9_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_9_1  (
            .in0(N__6230),
            .in1(N__6161),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_9_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_9_2 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_9_2  (
            .in0(N__6732),
            .in1(N__5848),
            .in2(N__5774),
            .in3(N__6061),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10591),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_11_10_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_11_10_0  (
            .in0(N__6247),
            .in1(N__6428),
            .in2(_gnd_net_),
            .in3(N__6056),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_11_10_1 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_11_10_1  (
            .in0(N__6758),
            .in1(N__5869),
            .in2(N__5771),
            .in3(N__6710),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_11_10_2 .LUT_INIT=16'b1111111100011111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_11_10_2  (
            .in0(N__6029),
            .in1(N__6192),
            .in2(N__5768),
            .in3(N__6449),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10586),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_11_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_11_10_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_11_10_4  (
            .in0(N__11083),
            .in1(N__12134),
            .in2(N__11408),
            .in3(N__6757),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN6_LC_11_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN6_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN6_LC_11_10_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN6_LC_11_10_5  (
            .in0(N__12135),
            .in1(N__11084),
            .in2(_gnd_net_),
            .in3(N__11308),
            .lcout(\U111_CYCLE_SM.TS_ENZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_11_12_3 .LUT_INIT=16'b0000000001011000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_11_12_3  (
            .in0(N__6316),
            .in1(N__6443),
            .in2(N__6362),
            .in3(N__6395),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10580),
            .ce(),
            .sr(N__10290));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_11_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5986),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(N__7905),
            .sr(N__7871));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_11_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_11_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_11_18_5  (
            .in0(N__5979),
            .in1(N__5942),
            .in2(_gnd_net_),
            .in3(N__8450),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_5  (
            .in0(N__8915),
            .in1(N__7331),
            .in2(_gnd_net_),
            .in3(N__5912),
            .lcout(un2_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_12_8_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_12_8_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_2_LC_12_8_0  (
            .in0(N__6265),
            .in1(N__6182),
            .in2(_gnd_net_),
            .in3(N__6055),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_8_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_8_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_8_1  (
            .in0(N__5873),
            .in1(N__6771),
            .in2(N__5858),
            .in3(N__6645),
            .lcout(\U111_CYCLE_SM.N_130_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_5  (
            .in0(N__6847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6717),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10590),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_8_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_8_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_8_7  (
            .in0(N__6846),
            .in1(N__7471),
            .in2(N__5849),
            .in3(N__6441),
            .lcout(\U111_CYCLE_SM.TS_EN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_12_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_12_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__6848),
            .in2(_gnd_net_),
            .in3(N__6390),
            .lcout(\U111_CYCLE_SM.un1_CYCLE_STATE_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_9_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_9_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_9_3  (
            .in0(N__6167),
            .in1(N__6266),
            .in2(_gnd_net_),
            .in3(N__6060),
            .lcout(\U111_CYCLE_SM.N_160 ),
            .ltout(\U111_CYCLE_SM.N_160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_9_4 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_9_4  (
            .in0(N__6718),
            .in1(N__6439),
            .in2(N__6119),
            .in3(N__6391),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10585),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_7  (
            .in0(N__6719),
            .in1(N__7448),
            .in2(_gnd_net_),
            .in3(N__6320),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10585),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_LC_12_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_12_10_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_12_10_0  (
            .in0(N__6115),
            .in1(N__6440),
            .in2(N__6092),
            .in3(N__6392),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10582),
            .ce(),
            .sr(N__10287));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_12_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_12_10_1 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_12_10_1  (
            .in0(N__6393),
            .in1(N__6116),
            .in2(N__7538),
            .in3(N__6091),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10582),
            .ce(),
            .sr(N__10287));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_12_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_12_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__7516),
            .in2(_gnd_net_),
            .in3(N__7533),
            .lcout(),
            .ltout(\U111_CYCLE_SM.PORT_MISMATCH_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_12_10_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_12_10_3  (
            .in0(N__7822),
            .in1(N__6850),
            .in2(N__6065),
            .in3(N__7472),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10582),
            .ce(),
            .sr(N__10287));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__6062),
            .in2(_gnd_net_),
            .in3(N__6646),
            .lcout(\U111_CYCLE_SM.N_142_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_11_3 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_11_3  (
            .in0(N__6337),
            .in1(N__6429),
            .in2(N__6023),
            .in3(N__6357),
            .lcout(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ),
            .ltout(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_11_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_11_4  (
            .in0(N__6276),
            .in1(N__7439),
            .in2(N__6452),
            .in3(N__6647),
            .lcout(\U111_CYCLE_SM.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNO_0_1_LC_12_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNO_0_1_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNO_0_1_LC_12_12_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNO_0_1_LC_12_12_3  (
            .in0(N__6314),
            .in1(N__6442),
            .in2(_gnd_net_),
            .in3(N__6394),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_132_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_12_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_12_12_4 .LUT_INIT=16'b0110000010100000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_12_12_4  (
            .in0(N__6338),
            .in1(N__6358),
            .in2(N__6341),
            .in3(N__6315),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10576),
            .ce(),
            .sr(N__10291));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7392),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10572),
            .ce(N__7903),
            .sr(N__7861));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_14_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_14_1  (
            .in0(N__6285),
            .in1(N__6201),
            .in2(_gnd_net_),
            .in3(N__6635),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2 ),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_12_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_12_14_2 .LUT_INIT=16'b0011001111110011;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__6734),
            .in2(N__6326),
            .in3(N__7234),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_12_14_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_12_14_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6323),
            .in3(N__6313),
            .lcout(\U111_CYCLE_SM.N_159_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_14_4 .LUT_INIT=16'b0010111100111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_14_4  (
            .in0(N__7447),
            .in1(N__6286),
            .in2(N__6206),
            .in3(N__6128),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_14_5 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_14_5  (
            .in0(N__6733),
            .in1(N__7484),
            .in2(N__6650),
            .in3(N__6636),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6995),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7141),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_12_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_12_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_12_15_3  (
            .in0(N__7066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_12_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_12_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_12_15_5  (
            .in0(N__6613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6918),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7200),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(N__7904),
            .sr(N__7872));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_12_16_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_12_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_12_16_1  (
            .in0(N__6600),
            .in1(N__6575),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_17_5.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6548),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_12_17_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_12_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_12_17_6  (
            .in0(N__8487),
            .in1(N__6491),
            .in2(_gnd_net_),
            .in3(N__8975),
            .lcout(un2_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_19_0  (
            .in0(N__7223),
            .in1(N__7210),
            .in2(_gnd_net_),
            .in3(N__8442),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_6  (
            .in0(N__7140),
            .in1(N__7106),
            .in2(_gnd_net_),
            .in3(N__8443),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_12_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_12_20_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_12_20_1  (
            .in0(N__7065),
            .in1(N__7031),
            .in2(_gnd_net_),
            .in3(N__8446),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_20_5  (
            .in0(N__7007),
            .in1(N__6994),
            .in2(_gnd_net_),
            .in3(N__8445),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_20_6  (
            .in0(N__8444),
            .in1(N__6935),
            .in2(_gnd_net_),
            .in3(N__6925),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_13_8_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_13_8_6 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_13_8_6  (
            .in0(N__8763),
            .in1(N__6851),
            .in2(N__6866),
            .in3(N__7473),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10597),
            .ce(),
            .sr(N__10296));
    defparam \U111_CYCLE_SM.A2_EN_LC_13_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_13_9_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_13_9_6  (
            .in0(N__6802),
            .in1(N__6849),
            .in2(_gnd_net_),
            .in3(N__6818),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10592),
            .ce(),
            .sr(N__10292));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_13_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_13_9_7 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_13_9_7  (
            .in0(N__7238),
            .in1(N__6790),
            .in2(N__8384),
            .in3(N__6778),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10592),
            .ce(),
            .sr(N__10292));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_13_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_13_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_13_10_1  (
            .in0(N__7247),
            .in1(N__7282),
            .in2(_gnd_net_),
            .in3(N__8368),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_3  (
            .in0(N__7443),
            .in1(N__7537),
            .in2(N__7520),
            .in3(N__7480),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10583),
            .ce(),
            .sr(N__10293));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_12_2  (
            .in0(N__8385),
            .in1(N__7295),
            .in2(_gnd_net_),
            .in3(N__7324),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_12_7  (
            .in0(N__7393),
            .in1(N__7358),
            .in2(_gnd_net_),
            .in3(N__8386),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7323),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10577),
            .ce(N__7906),
            .sr(N__7877));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7281),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10577),
            .ce(N__7906),
            .sr(N__7877));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_13_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_13_14_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_13_14_0  (
            .in0(N__10823),
            .in1(N__12088),
            .in2(N__11553),
            .in3(N__12527),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10574),
            .ce(N__10429),
            .sr(N__10299));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8492),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_15_1  (
            .in0(N__7637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8544),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_13_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_13_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7703),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7784),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8618),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(N__7907),
            .sr(N__7876));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_13_16_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_13_16_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__11554),
            .in2(_gnd_net_),
            .in3(N__7829),
            .lcout(TAn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_17_5  (
            .in0(N__8407),
            .in1(N__7793),
            .in2(_gnd_net_),
            .in3(N__7773),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_13_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_13_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_13_18_5  (
            .in0(N__8437),
            .in1(N__7712),
            .in2(_gnd_net_),
            .in3(N__7698),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_19_2  (
            .in0(N__7632),
            .in1(N__7592),
            .in2(_gnd_net_),
            .in3(N__8438),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_19_5  (
            .in0(N__8439),
            .in1(N__8630),
            .in2(_gnd_net_),
            .in3(N__8614),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_1  (
            .in0(N__8440),
            .in1(N__8561),
            .in2(_gnd_net_),
            .in3(N__8551),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_20_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_20_2  (
            .in0(N__8491),
            .in1(N__8441),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_14_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_14_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_14_20_3  (
            .in0(N__8308),
            .in1(N__8279),
            .in2(_gnd_net_),
            .in3(N__8997),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_15_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_15_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_15_12_0  (
            .in0(N__8240),
            .in1(N__8215),
            .in2(_gnd_net_),
            .in3(N__9008),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_15_19_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_15_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_15_19_7  (
            .in0(N__9006),
            .in1(N__8156),
            .in2(_gnd_net_),
            .in3(N__8111),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_15_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_15_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_15_20_2  (
            .in0(N__8075),
            .in1(N__8047),
            .in2(_gnd_net_),
            .in3(N__8998),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_16_15_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_16_15_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_16_15_7  (
            .in0(N__8974),
            .in1(N__7981),
            .in2(_gnd_net_),
            .in3(N__7946),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_16_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_16_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_16_20_1  (
            .in0(N__9512),
            .in1(N__9476),
            .in2(_gnd_net_),
            .in3(N__9000),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_16_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_16_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_16_20_7  (
            .in0(N__9434),
            .in1(N__9412),
            .in2(_gnd_net_),
            .in3(N__8999),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_17_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_17_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_17_20_6  (
            .in0(N__9337),
            .in1(N__9302),
            .in2(_gnd_net_),
            .in3(N__9001),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_17_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_17_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_17_20_7  (
            .in0(N__9002),
            .in1(N__9260),
            .in2(_gnd_net_),
            .in3(N__9235),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_18_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_18_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_18_9_6  (
            .in0(N__9185),
            .in1(N__9163),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_18_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_18_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_18_18_2  (
            .in0(N__9110),
            .in1(N__9091),
            .in2(_gnd_net_),
            .in3(N__9018),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_2  (
            .in0(N__9019),
            .in1(N__8716),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_3  (
            .in0(N__12526),
            .in1(N__11013),
            .in2(N__11932),
            .in3(N__11475),
            .lcout(READ_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10578),
            .ce(N__10432),
            .sr(N__10304));
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_2.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_2.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_4_LC_19_20_2 (
            .in0(N__9620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_184_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_4  (
            .in0(N__12505),
            .in1(N__10930),
            .in2(N__11942),
            .in3(N__11476),
            .lcout(READ_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10581),
            .ce(N__10434),
            .sr(N__10305));
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_1.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_1.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_2_LC_20_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(N_182_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_18_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_18_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_18_0  (
            .in0(N__10867),
            .in1(N__12443),
            .in2(N__12094),
            .in3(N__11503),
            .lcout(READ_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10593),
            .ce(N__10436),
            .sr(N__10308));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_19_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_19_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_19_0  (
            .in0(N__10821),
            .in1(N__12444),
            .in2(N__11943),
            .in3(N__11477),
            .lcout(READ_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10587),
            .ce(N__10437),
            .sr(N__10310));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_22_19_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_22_19_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_22_19_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_22_19_6  (
            .in0(N__10822),
            .in1(N__12445),
            .in2(N__11944),
            .in3(N__11478),
            .lcout(READ_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10587),
            .ce(N__10437),
            .sr(N__10310));
    defparam D_UU_040_iobuf_RNO_0_LC_22_20_3.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_0_LC_22_20_3.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_0_LC_22_20_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_0_LC_22_20_3 (
            .in0(N__9578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_180_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_5.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_5.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_5.LUT_INIT=16'b0011001100110011;
    LogicCell40 D_UU_040_iobuf_RNO_7_LC_22_20_5 (
            .in0(_gnd_net_),
            .in1(N__9554),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_187_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_6_LC_22_20_6.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_6_LC_22_20_6.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_6_LC_22_20_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_6_LC_22_20_6 (
            .in0(N__9533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_186_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_3_LC_23_2_2.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_3_LC_23_2_2.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_3_LC_23_2_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_3_LC_23_2_2 (
            .in0(N__9713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_1_LC_23_2_7.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_1_LC_23_2_7.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_1_LC_23_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_1_LC_23_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9707),
            .lcout(N_205_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_23_3_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_23_3_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_23_3_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_23_3_6  (
            .in0(N__11014),
            .in1(N__12132),
            .in2(N__11349),
            .in3(N__12705),
            .lcout(READ_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10626),
            .ce(N__10443),
            .sr(N__10309));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_23_4_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_23_4_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_23_4_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_23_4_3  (
            .in0(N__12595),
            .in1(N__11001),
            .in2(N__12162),
            .in3(N__11465),
            .lcout(READ_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10623),
            .ce(N__10438),
            .sr(N__10306));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_23_4_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_23_4_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_23_4_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_23_4_6  (
            .in0(N__11002),
            .in1(N__12131),
            .in2(N__11548),
            .in3(N__12596),
            .lcout(READ_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10623),
            .ce(N__10438),
            .sr(N__10306));
    defparam D_LM_040_iobuf_RNO_0_LC_23_5_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_0_LC_23_5_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_0_LC_23_5_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_0_LC_23_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9680),
            .lcout(N_196_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_23_6_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_23_6_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_23_6_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_23_6_4  (
            .in0(N__10925),
            .in1(N__12076),
            .in2(N__11549),
            .in3(N__12591),
            .lcout(READ_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10620),
            .ce(N__10435),
            .sr(N__10302));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_10_6.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_10_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10631),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_18_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_18_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_18_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_18_3  (
            .in0(N__10866),
            .in1(N__11953),
            .in2(N__12504),
            .in3(N__11504),
            .lcout(READ_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10598),
            .ce(N__10439),
            .sr(N__10311));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_23_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_23_19_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_23_19_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_23_19_4  (
            .in0(N__10931),
            .in1(N__11945),
            .in2(N__11550),
            .in3(N__12430),
            .lcout(READ_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10594),
            .ce(N__10442),
            .sr(N__10314));
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_1.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_1.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_5_LC_23_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9887),
            .lcout(N_185_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_3.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_3.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_5_LC_23_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9863),
            .lcout(N_193_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_4_LC_24_2_4.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_4_LC_24_2_4.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_4_LC_24_2_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_4_LC_24_2_4 (
            .in0(N__9827),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_208_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_24_3_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_24_3_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_24_3_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_24_3_2  (
            .in0(N__10929),
            .in1(N__12133),
            .in2(N__12704),
            .in3(N__11358),
            .lcout(READ_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10627),
            .ce(N__10445),
            .sr(N__10313));
    defparam D_LL_040_iobuf_RNO_0_LC_24_4_1.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_0_LC_24_4_1.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_0_LC_24_4_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_0_LC_24_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9974),
            .lcout(N_204_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_2.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_2.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_6_LC_24_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9803),
            .lcout(N_210_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_3.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_3.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_2_LC_24_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9968),
            .lcout(N_206_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_5_LC_24_4_5.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_5_LC_24_4_5.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_5_LC_24_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_5_LC_24_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9980),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_5_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_5_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_5_5 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_5_5  (
            .in0(N__12594),
            .in1(N__10928),
            .in2(N__11913),
            .in3(N__11363),
            .lcout(READ_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10624),
            .ce(N__10440),
            .sr(N__10307));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_5_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_5_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_5_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_5_6  (
            .in0(N__10926),
            .in1(N__11817),
            .in2(N__11472),
            .in3(N__12592),
            .lcout(READ_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10624),
            .ce(N__10440),
            .sr(N__10307));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_24_5_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_24_5_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_24_5_7 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_24_5_7  (
            .in0(N__12593),
            .in1(N__10927),
            .in2(N__11912),
            .in3(N__11362),
            .lcout(READ_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10624),
            .ce(N__10440),
            .sr(N__10307));
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_1.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_1.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_1_LC_24_6_1 (
            .in0(N__10064),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_197_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_4.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_4.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_7_LC_24_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9902),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_2_LC_24_7_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_2_LC_24_7_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_2_LC_24_7_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_2_LC_24_7_2 (
            .in0(N__10070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_198_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_3_LC_24_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9893),
            .lcout(N_199_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_24_8_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_24_8_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_24_8_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_24_8_0  (
            .in0(N__12074),
            .in1(N__10848),
            .in2(N__12503),
            .in3(N__11369),
            .lcout(READ_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10618),
            .ce(N__10433),
            .sr(N__10301));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_8_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_8_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_8_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_8_3  (
            .in0(N__10849),
            .in1(N__12426),
            .in2(N__11474),
            .in3(N__12075),
            .lcout(READ_CYCLE_ACTIVE_rep31_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10618),
            .ce(N__10433),
            .sr(N__10301));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_4  (
            .in0(N__12073),
            .in1(N__10847),
            .in2(N__12502),
            .in3(N__11368),
            .lcout(READ_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10618),
            .ce(N__10433),
            .sr(N__10301));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_24_8_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_24_8_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_24_8_5 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_24_8_5  (
            .in0(N__10846),
            .in1(N__12419),
            .in2(N__11473),
            .in3(N__12072),
            .lcout(READ_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10618),
            .ce(N__10433),
            .sr(N__10301));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_24_8_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_24_8_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_24_8_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_24_8_6  (
            .in0(N__12071),
            .in1(N__10845),
            .in2(N__12501),
            .in3(N__11364),
            .lcout(READ_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10618),
            .ce(N__10433),
            .sr(N__10301));
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_1.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_1.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_4_LC_24_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10016),
            .lcout(N_200_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_3.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_3.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_0_LC_24_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10010),
            .lcout(N_188_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_5_LC_24_9_5.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_5_LC_24_9_5.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_5_LC_24_9_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_5_LC_24_9_5 (
            .in0(N__10031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_201_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_10_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_10_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_10_4  (
            .in0(N__11373),
            .in1(N__10840),
            .in2(N__12069),
            .in3(N__12414),
            .lcout(READ_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10615),
            .ce(N__10430),
            .sr(N__10300));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_10_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_10_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_10_7  (
            .in0(N__10841),
            .in1(N__12415),
            .in2(N__12070),
            .in3(N__11374),
            .lcout(READ_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10615),
            .ce(N__10430),
            .sr(N__10300));
    defparam D_UM_040_iobuf_RNO_2_LC_24_12_4.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_2_LC_24_12_4.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_2_LC_24_12_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_2_LC_24_12_4 (
            .in0(N__10115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_190_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_6_LC_24_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10121),
            .lcout(N_194_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_1  (
            .in0(N__10764),
            .in1(N__12327),
            .in2(N__11914),
            .in3(N__11377),
            .lcout(READ_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10608),
            .ce(N__10431),
            .sr(N__10303));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_2  (
            .in0(N__11378),
            .in1(N__10765),
            .in2(N__12412),
            .in3(N__11829),
            .lcout(READ_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10608),
            .ce(N__10431),
            .sr(N__10303));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_4  (
            .in0(N__11376),
            .in1(N__10763),
            .in2(N__12411),
            .in3(N__11825),
            .lcout(READ_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10608),
            .ce(N__10431),
            .sr(N__10303));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_13_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_13_6 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_13_6  (
            .in0(N__11375),
            .in1(N__10762),
            .in2(N__12410),
            .in3(N__11824),
            .lcout(READ_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10608),
            .ce(N__10431),
            .sr(N__10303));
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_1.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_1.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_6_LC_24_14_1 (
            .in0(N__10109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_202_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_5.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_5.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_7_LC_24_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10091),
            .lcout(N_203_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_24_17_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_24_17_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_24_17_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_24_17_0  (
            .in0(N__10794),
            .in1(N__12334),
            .in2(N__11816),
            .in3(N__11483),
            .lcout(READ_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10602),
            .ce(N__10441),
            .sr(N__10312));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_17_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_17_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_17_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_17_6  (
            .in0(N__10795),
            .in1(N__11746),
            .in2(N__11551),
            .in3(N__12335),
            .lcout(READ_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10602),
            .ce(N__10441),
            .sr(N__10312));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_17_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_17_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_17_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_17_7  (
            .in0(N__11482),
            .in1(N__10793),
            .in2(N__12413),
            .in3(N__11742),
            .lcout(READ_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10602),
            .ce(N__10441),
            .sr(N__10312));
    defparam D_UM_040_iobuf_RNO_1_LC_24_18_3.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_1_LC_24_18_3.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_1_LC_24_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_1_LC_24_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12782),
            .lcout(N_189_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_3_LC_24_18_4.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_3_LC_24_18_4.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_3_LC_24_18_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_3_LC_24_18_4 (
            .in0(N__12761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_191_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_7_LC_24_18_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_7_LC_24_18_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_7_LC_24_18_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_7_LC_24_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12740),
            .lcout(N_195_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_19_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_19_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_19_2  (
            .in0(N__10864),
            .in1(N__12337),
            .in2(N__12030),
            .in3(N__11488),
            .lcout(READ_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10599),
            .ce(N__10444),
            .sr(N__10315));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_19_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_19_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_19_4  (
            .in0(N__10863),
            .in1(N__12336),
            .in2(N__12029),
            .in3(N__11487),
            .lcout(READ_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10599),
            .ce(N__10444),
            .sr(N__10315));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_19_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_19_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_19_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_19_7  (
            .in0(N__12338),
            .in1(N__11952),
            .in2(N__11552),
            .in3(N__10865),
            .lcout(READ_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10599),
            .ce(N__10444),
            .sr(N__10315));
    defparam D_UU_040_iobuf_RNO_1_LC_24_20_2.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_1_LC_24_20_2.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_1_LC_24_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_1_LC_24_20_2 (
            .in0(N__10163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_181_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_4_LC_24_20_3.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_4_LC_24_20_3.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_4_LC_24_20_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_4_LC_24_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10142),
            .lcout(N_192_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_3_LC_24_20_5.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_3_LC_24_20_5.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_3_LC_24_20_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_3_LC_24_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12800),
            .lcout(N_183_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 31 2025 15:09:50

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_UU_AMIGA,
    D_LL_AMIGA,
    D_UM_AMIGA,
    D_LM_AMIGA,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    D_LL_040,
    A_AMIGA,
    A_040,
    SIZ,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    TBIn,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LL_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TEAn;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    input TBIn;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    inout TACKn;
    input BGn;

    wire N__8833;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8808;
    wire N__8807;
    wire N__8806;
    wire N__8799;
    wire N__8798;
    wire N__8797;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8754;
    wire N__8753;
    wire N__8752;
    wire N__8745;
    wire N__8744;
    wire N__8743;
    wire N__8736;
    wire N__8735;
    wire N__8734;
    wire N__8727;
    wire N__8726;
    wire N__8725;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8709;
    wire N__8708;
    wire N__8707;
    wire N__8700;
    wire N__8699;
    wire N__8698;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8655;
    wire N__8654;
    wire N__8653;
    wire N__8646;
    wire N__8645;
    wire N__8644;
    wire N__8637;
    wire N__8636;
    wire N__8635;
    wire N__8628;
    wire N__8627;
    wire N__8626;
    wire N__8619;
    wire N__8618;
    wire N__8617;
    wire N__8610;
    wire N__8609;
    wire N__8608;
    wire N__8601;
    wire N__8600;
    wire N__8599;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8574;
    wire N__8573;
    wire N__8572;
    wire N__8565;
    wire N__8564;
    wire N__8563;
    wire N__8556;
    wire N__8555;
    wire N__8554;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8529;
    wire N__8528;
    wire N__8527;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8511;
    wire N__8510;
    wire N__8509;
    wire N__8502;
    wire N__8501;
    wire N__8500;
    wire N__8493;
    wire N__8492;
    wire N__8491;
    wire N__8484;
    wire N__8483;
    wire N__8482;
    wire N__8475;
    wire N__8474;
    wire N__8473;
    wire N__8466;
    wire N__8465;
    wire N__8464;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8448;
    wire N__8447;
    wire N__8446;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8421;
    wire N__8420;
    wire N__8419;
    wire N__8412;
    wire N__8411;
    wire N__8410;
    wire N__8403;
    wire N__8402;
    wire N__8401;
    wire N__8394;
    wire N__8393;
    wire N__8392;
    wire N__8385;
    wire N__8384;
    wire N__8383;
    wire N__8376;
    wire N__8375;
    wire N__8374;
    wire N__8367;
    wire N__8366;
    wire N__8365;
    wire N__8358;
    wire N__8357;
    wire N__8356;
    wire N__8349;
    wire N__8348;
    wire N__8347;
    wire N__8340;
    wire N__8339;
    wire N__8338;
    wire N__8331;
    wire N__8330;
    wire N__8329;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8313;
    wire N__8312;
    wire N__8311;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8295;
    wire N__8294;
    wire N__8293;
    wire N__8286;
    wire N__8285;
    wire N__8284;
    wire N__8277;
    wire N__8276;
    wire N__8275;
    wire N__8268;
    wire N__8267;
    wire N__8266;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8241;
    wire N__8240;
    wire N__8239;
    wire N__8232;
    wire N__8231;
    wire N__8230;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8205;
    wire N__8204;
    wire N__8203;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8178;
    wire N__8177;
    wire N__8176;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8160;
    wire N__8159;
    wire N__8158;
    wire N__8151;
    wire N__8150;
    wire N__8149;
    wire N__8142;
    wire N__8141;
    wire N__8140;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8106;
    wire N__8105;
    wire N__8104;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8088;
    wire N__8087;
    wire N__8086;
    wire N__8079;
    wire N__8078;
    wire N__8077;
    wire N__8070;
    wire N__8069;
    wire N__8068;
    wire N__8061;
    wire N__8060;
    wire N__8059;
    wire N__8052;
    wire N__8051;
    wire N__8050;
    wire N__8043;
    wire N__8042;
    wire N__8041;
    wire N__8034;
    wire N__8033;
    wire N__8032;
    wire N__8025;
    wire N__8024;
    wire N__8023;
    wire N__8016;
    wire N__8015;
    wire N__8014;
    wire N__8007;
    wire N__8006;
    wire N__8005;
    wire N__7998;
    wire N__7997;
    wire N__7996;
    wire N__7989;
    wire N__7988;
    wire N__7987;
    wire N__7980;
    wire N__7979;
    wire N__7978;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7921;
    wire N__7918;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7891;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7811;
    wire N__7810;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7806;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7791;
    wire N__7786;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7742;
    wire N__7741;
    wire N__7740;
    wire N__7739;
    wire N__7738;
    wire N__7737;
    wire N__7736;
    wire N__7703;
    wire N__7700;
    wire N__7699;
    wire N__7696;
    wire N__7695;
    wire N__7692;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7673;
    wire N__7670;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7649;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7637;
    wire N__7636;
    wire N__7635;
    wire N__7630;
    wire N__7627;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7586;
    wire N__7585;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7579;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7552;
    wire N__7549;
    wire N__7548;
    wire N__7545;
    wire N__7544;
    wire N__7543;
    wire N__7542;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7496;
    wire N__7493;
    wire N__7488;
    wire N__7485;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7471;
    wire N__7470;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7448;
    wire N__7445;
    wire N__7444;
    wire N__7443;
    wire N__7442;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7427;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7399;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7264;
    wire N__7263;
    wire N__7260;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7213;
    wire N__7210;
    wire N__7209;
    wire N__7208;
    wire N__7207;
    wire N__7202;
    wire N__7199;
    wire N__7194;
    wire N__7193;
    wire N__7192;
    wire N__7191;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7187;
    wire N__7180;
    wire N__7173;
    wire N__7172;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7147;
    wire N__7142;
    wire N__7137;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7125;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6956;
    wire N__6955;
    wire N__6950;
    wire N__6949;
    wire N__6948;
    wire N__6947;
    wire N__6946;
    wire N__6945;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6932;
    wire N__6927;
    wire N__6922;
    wire N__6921;
    wire N__6920;
    wire N__6919;
    wire N__6918;
    wire N__6917;
    wire N__6916;
    wire N__6915;
    wire N__6912;
    wire N__6907;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6895;
    wire N__6890;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6877;
    wire N__6870;
    wire N__6865;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6835;
    wire N__6834;
    wire N__6833;
    wire N__6832;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6802;
    wire N__6797;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6773;
    wire N__6770;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6700;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6549;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6532;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6495;
    wire N__6490;
    wire N__6487;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6437;
    wire N__6436;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6401;
    wire N__6398;
    wire N__6397;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6379;
    wire N__6376;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6332;
    wire N__6331;
    wire N__6330;
    wire N__6329;
    wire N__6328;
    wire N__6323;
    wire N__6320;
    wire N__6315;
    wire N__6308;
    wire N__6307;
    wire N__6306;
    wire N__6303;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6274;
    wire N__6271;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6215;
    wire N__6210;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6186;
    wire N__6181;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5656;
    wire N__5655;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5628;
    wire N__5625;
    wire N__5620;
    wire N__5615;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5461;
    wire N__5458;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5446;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5432;
    wire N__5429;
    wire N__5428;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5393;
    wire N__5390;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5349;
    wire N__5348;
    wire N__5347;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5314;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5287;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5266;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5215;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5050;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4824;
    wire N__4819;
    wire N__4816;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4759;
    wire N__4754;
    wire N__4751;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4743;
    wire N__4742;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4730;
    wire N__4729;
    wire N__4728;
    wire N__4727;
    wire N__4726;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4703;
    wire N__4702;
    wire N__4701;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4678;
    wire N__4675;
    wire N__4674;
    wire N__4667;
    wire N__4664;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4660;
    wire N__4659;
    wire N__4658;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4650;
    wire N__4649;
    wire N__4648;
    wire N__4643;
    wire N__4640;
    wire N__4639;
    wire N__4638;
    wire N__4637;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4585;
    wire N__4584;
    wire N__4575;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4559;
    wire N__4552;
    wire N__4549;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4468;
    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4375;
    wire N__4374;
    wire N__4373;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4356;
    wire N__4355;
    wire N__4354;
    wire N__4353;
    wire N__4342;
    wire N__4341;
    wire N__4340;
    wire N__4339;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4323;
    wire N__4322;
    wire N__4321;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4304;
    wire N__4303;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4287;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4262;
    wire N__4259;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4246;
    wire N__4245;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4229;
    wire N__4226;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4174;
    wire N__4171;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4155;
    wire N__4150;
    wire N__4145;
    wire N__4142;
    wire N__4135;
    wire N__4130;
    wire N__4127;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3988;
    wire N__3985;
    wire N__3984;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3914;
    wire N__3911;
    wire N__3910;
    wire N__3909;
    wire N__3906;
    wire N__3901;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3339;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3277;
    wire N__3276;
    wire N__3273;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire TCIn_c;
    wire VCCG0;
    wire GNDG0;
    wire TAn_in;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire D_LL_AMIGA_in_0;
    wire un1_D_LL_AMIGA_0;
    wire D_LL_AMIGA_in_1;
    wire un1_D_LL_AMIGA_1;
    wire D_LL_AMIGA_in_3;
    wire un1_D_LL_AMIGA_3;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire LBENn_c_i;
    wire D_LM_AMIGA_in_4;
    wire un1_D_LM_AMIGA_4;
    wire D_LM_AMIGA_in_5;
    wire un1_D_LM_AMIGA_5;
    wire D_LM_AMIGA_in_7;
    wire un1_D_LM_AMIGA_7;
    wire D_LM_AMIGA_in_6;
    wire un1_D_LM_AMIGA_6;
    wire CONSTANT_ONE_NET;
    wire D_LM_040_in_7;
    wire D_UU_040_in_7;
    wire un1_D_UU_040_7;
    wire D_LM_AMIGA_in_3;
    wire un1_D_LM_AMIGA_3;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_UU_040_in_1;
    wire D_LM_040_in_1;
    wire un1_D_UU_040_1;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_UU_040_in_0;
    wire D_LM_040_in_0;
    wire un1_D_UU_040_0;
    wire un1_D_UM_AMIGA_0;
    wire D_LM_AMIGA_in_1;
    wire un1_D_LM_AMIGA_1;
    wire D_UM_AMIGA_in_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire un1_D_UM_AMIGA_1;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UU_AMIGA_1;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire un1_D_UM_040_5;
    wire LBENn_c_i_0;
    wire D_LL_AMIGA_in_6;
    wire un1_D_LL_AMIGA_6;
    wire D_LL_AMIGA_in_5;
    wire un1_D_LL_AMIGA_5;
    wire A_040_c_1;
    wire D_LL_AMIGA_in_7;
    wire un1_D_LL_AMIGA_7;
    wire D_LM_AMIGA_in_0;
    wire un1_D_LM_AMIGA_0;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire D_UU_AMIGA_1_i;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire \U111_CYCLE_SM.FLIP_WORD_2 ;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire \U111_CYCLE_SM.PORT_MISMATCH_2 ;
    wire \U111_CYCLE_SM.N_123_0_cascade_ ;
    wire \U111_CYCLE_SM.N_121_0 ;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_0 ;
    wire D_UU_040_1_i;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire un1_D_UU_AMIGA_6;
    wire D_UU_AMIGA_in_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire un1_D_UU_AMIGA_0;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire un1_D_UU_AMIGA_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire D_UM_AMIGA_in_5;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire D_UU_AMIGA_in_7;
    wire un1_D_UU_AMIGA_7;
    wire D_LL_AMIGA_in_2;
    wire un1_D_LL_AMIGA_2;
    wire D_LL_AMIGA_in_4;
    wire un1_D_LL_AMIGA_4;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire \U111_CYCLE_SM.N_148 ;
    wire \U111_CYCLE_SM.N_148_cascade_ ;
    wire \U111_CYCLE_SM.TS_EN_6 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ;
    wire LBENn_c;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire TAn_1_i;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire \U111_CYCLE_SM.N_135_cascade_ ;
    wire \U111_CYCLE_SM.N_128_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire TEAn_c;
    wire RESETn_c;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire D_LM_AMIGA_in_2;
    wire D_UU_AMIGA_in_2;
    wire un1_D_LM_AMIGA_2;
    wire \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ;
    wire D_UM_AMIGA_in_4;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire un1_D_UM_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire D_UU_AMIGA_in_3;
    wire un1_D_UU_AMIGA_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire D_UM_AMIGA_in_3;
    wire un1_D_UM_AMIGA_3;
    wire D_UM_040_in_3;
    wire D_LL_040_in_3;
    wire un1_D_UM_040_3;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire D_UM_040_in_4;
    wire D_LL_040_in_4;
    wire un1_D_UM_040_4;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire PORTSIZE_c;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ;
    wire TS_CPUn_c;
    wire RnW_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ;
    wire CLK40;
    wire RESETn_c_i;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire TBIn_c;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0 ;
    wire TACKn_in;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire \U111_CYCLE_SM.N_136 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire D_UM_AMIGA_in_2;
    wire un1_D_UM_AMIGA_2;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire un1_D_UM_AMIGA_6;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LM_040_in_5;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire D_UU_040_in_5;
    wire un1_D_UU_040_5;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__3121),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__8833));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__8833),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__8817),
            .DIN(N__8816),
            .DOUT(N__8815),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__8817),
            .PADOUT(N__8816),
            .PADIN(N__8815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__8808),
            .DIN(N__8807),
            .DOUT(N__8806),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__8808),
            .PADOUT(N__8807),
            .PADIN(N__8806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4585),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__6005),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__8799),
            .DIN(N__8798),
            .DOUT(N__8797),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__8799),
            .PADOUT(N__8798),
            .PADIN(N__8797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5372),
            .DIN0(TAn_in),
            .DOUT0(N__7553),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__8790),
            .DIN(N__8789),
            .DOUT(N__8788),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__8790),
            .PADOUT(N__8789),
            .PADIN(N__8788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4373),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__7334),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__8781),
            .DIN(N__8780),
            .DOUT(N__8779),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__8781),
            .PADOUT(N__8780),
            .PADIN(N__8779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4337),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__7943),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__8772),
            .DIN(N__8771),
            .DOUT(N__8770),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__8772),
            .PADOUT(N__8771),
            .PADIN(N__8770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4660),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__4964),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__8763),
            .DIN(N__8762),
            .DOUT(N__8761),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__8763),
            .PADOUT(N__8762),
            .PADIN(N__8761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__8754),
            .DIN(N__8753),
            .DOUT(N__8752),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__8754),
            .PADOUT(N__8753),
            .PADIN(N__8752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4726),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__3590),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__8745),
            .DIN(N__8744),
            .DOUT(N__8743),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__8745),
            .PADOUT(N__8744),
            .PADIN(N__8743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4372),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__5797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__8736),
            .DIN(N__8735),
            .DOUT(N__8734),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8736),
            .PADOUT(N__8735),
            .PADIN(N__8734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4246),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__5924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__8727),
            .DIN(N__8726),
            .DOUT(N__8725),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__8727),
            .PADOUT(N__8726),
            .PADIN(N__8725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4701),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__6077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__8718),
            .DIN(N__8717),
            .DOUT(N__8716),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__8718),
            .PADOUT(N__8717),
            .PADIN(N__8716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5276),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__8709),
            .DIN(N__8708),
            .DOUT(N__8707),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__8709),
            .PADOUT(N__8708),
            .PADIN(N__8707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__8700),
            .DIN(N__8699),
            .DOUT(N__8698),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__8700),
            .PADOUT(N__8699),
            .PADIN(N__8698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4304),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__6662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__8691),
            .DIN(N__8690),
            .DOUT(N__8689),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__8691),
            .PADOUT(N__8690),
            .PADIN(N__8689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4727),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__4418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__8682),
            .DIN(N__8681),
            .DOUT(N__8680),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8682),
            .PADOUT(N__8681),
            .PADIN(N__8680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4336),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__2612),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__8673),
            .DIN(N__8672),
            .DOUT(N__8671),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8673),
            .PADOUT(N__8672),
            .PADIN(N__8671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4257),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__3551),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__8664),
            .DIN(N__8663),
            .DOUT(N__8662),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__8664),
            .PADOUT(N__8663),
            .PADIN(N__8662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2795),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__8655),
            .DIN(N__8654),
            .DOUT(N__8653),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__8655),
            .PADOUT(N__8654),
            .PADIN(N__8653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4663),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__3167),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__8646),
            .DIN(N__8645),
            .DOUT(N__8644),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__8646),
            .PADOUT(N__8645),
            .PADIN(N__8644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4702),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__6149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__8637),
            .DIN(N__8636),
            .DOUT(N__8635),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__8637),
            .PADOUT(N__8636),
            .PADIN(N__8635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3984),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__8628),
            .DIN(N__8627),
            .DOUT(N__8626),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__8628),
            .PADOUT(N__8627),
            .PADIN(N__8626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4355),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__3431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__8619),
            .DIN(N__8618),
            .DOUT(N__8617),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__8619),
            .PADOUT(N__8618),
            .PADIN(N__8617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4678),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__3308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__8610),
            .DIN(N__8609),
            .DOUT(N__8608),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__8610),
            .PADOUT(N__8609),
            .PADIN(N__8608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__8601),
            .DIN(N__8600),
            .DOUT(N__8599),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__8601),
            .PADOUT(N__8600),
            .PADIN(N__8599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4743),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__5072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__8592),
            .DIN(N__8591),
            .DOUT(N__8590),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__8592),
            .PADOUT(N__8591),
            .PADIN(N__8590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4338),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__5711),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__8583),
            .DIN(N__8582),
            .DOUT(N__8581),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__8583),
            .PADOUT(N__8582),
            .PADIN(N__8581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4253),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__3032),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__8574),
            .DIN(N__8573),
            .DOUT(N__8572),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__8574),
            .PADOUT(N__8573),
            .PADIN(N__8572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7877),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__8565),
            .DIN(N__8564),
            .DOUT(N__8563),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__8565),
            .PADOUT(N__8564),
            .PADIN(N__8563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4657),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__6518),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__8556),
            .DIN(N__8555),
            .DOUT(N__8554),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__8556),
            .PADOUT(N__8555),
            .PADIN(N__8554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__8547),
            .DIN(N__8546),
            .DOUT(N__8545),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__8547),
            .PADOUT(N__8546),
            .PADIN(N__8545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__8538),
            .DIN(N__8537),
            .DOUT(N__8536),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__8538),
            .PADOUT(N__8537),
            .PADIN(N__8536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4742),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__2723),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__8529),
            .DIN(N__8528),
            .DOUT(N__8527),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__8529),
            .PADOUT(N__8528),
            .PADIN(N__8527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4356),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__3737),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__8520),
            .DIN(N__8519),
            .DOUT(N__8518),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__8520),
            .PADOUT(N__8519),
            .PADIN(N__8518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4703),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__3239),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__8511),
            .DIN(N__8510),
            .DOUT(N__8509),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__8511),
            .PADOUT(N__8510),
            .PADIN(N__8509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4256),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__2885),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__8502),
            .DIN(N__8501),
            .DOUT(N__8500),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__8502),
            .PADOUT(N__8501),
            .PADIN(N__8500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4637),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__5477),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__8493),
            .DIN(N__8492),
            .DOUT(N__8491),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__8493),
            .PADOUT(N__8492),
            .PADIN(N__8491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4728),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__3653),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__8484),
            .DIN(N__8483),
            .DOUT(N__8482),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__8484),
            .PADOUT(N__8483),
            .PADIN(N__8482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4340),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__2657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__8475),
            .DIN(N__8474),
            .DOUT(N__8473),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__8475),
            .PADOUT(N__8474),
            .PADIN(N__8473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4254),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__7025),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__8466),
            .DIN(N__8465),
            .DOUT(N__8464),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__8466),
            .PADOUT(N__8465),
            .PADIN(N__8464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4286),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__7286),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__8457),
            .DIN(N__8456),
            .DOUT(N__8455),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__8457),
            .PADOUT(N__8456),
            .PADIN(N__8455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4662),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__6683),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__8448),
            .DIN(N__8447),
            .DOUT(N__8446),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__8448),
            .PADOUT(N__8447),
            .PADIN(N__8446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3719),
            .DIN0(TACKn_in),
            .DOUT0(N__2546),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__8439),
            .DIN(N__8438),
            .DOUT(N__8437),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__8439),
            .PADOUT(N__8438),
            .PADIN(N__8437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3992),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__8430),
            .DIN(N__8429),
            .DOUT(N__8428),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__8430),
            .PADOUT(N__8429),
            .PADIN(N__8428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4648),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__7370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__8421),
            .DIN(N__8420),
            .DOUT(N__8419),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__8421),
            .PADOUT(N__8420),
            .PADIN(N__8419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4730),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__5111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__8412),
            .DIN(N__8411),
            .DOUT(N__8410),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__8412),
            .PADOUT(N__8411),
            .PADIN(N__8410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2522),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__8403),
            .DIN(N__8402),
            .DOUT(N__8401),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__8403),
            .PADOUT(N__8402),
            .PADIN(N__8401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5576),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__8394),
            .DIN(N__8393),
            .DOUT(N__8392),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__8394),
            .PADOUT(N__8393),
            .PADIN(N__8392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4375),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__4055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__8385),
            .DIN(N__8384),
            .DOUT(N__8383),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8385),
            .PADOUT(N__8384),
            .PADIN(N__8383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4303),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__5753),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__8376),
            .DIN(N__8375),
            .DOUT(N__8374),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__8376),
            .PADOUT(N__8375),
            .PADIN(N__8374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4354),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__3821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TEAn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__8367),
            .DIN(N__8366),
            .DOUT(N__8365),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__8367),
            .PADOUT(N__8366),
            .PADIN(N__8365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__8358),
            .DIN(N__8357),
            .DOUT(N__8356),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__8358),
            .PADOUT(N__8357),
            .PADIN(N__8356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__8349),
            .DIN(N__8348),
            .DOUT(N__8347),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8349),
            .PADOUT(N__8348),
            .PADIN(N__8347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4323),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__7067),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__8340),
            .DIN(N__8339),
            .DOUT(N__8338),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__8340),
            .PADOUT(N__8339),
            .PADIN(N__8338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__8331),
            .DIN(N__8330),
            .DOUT(N__8329),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__8331),
            .PADOUT(N__8330),
            .PADIN(N__8329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4650),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3203),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__8322),
            .DIN(N__8321),
            .DOUT(N__8320),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__8322),
            .PADOUT(N__8321),
            .PADIN(N__8320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4638),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__7103),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__8313),
            .DIN(N__8312),
            .DOUT(N__8311),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__8313),
            .PADOUT(N__8312),
            .PADIN(N__8311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__8304),
            .DIN(N__8303),
            .DOUT(N__8302),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__8304),
            .PADOUT(N__8303),
            .PADIN(N__8302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4729),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__3692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__8295),
            .DIN(N__8294),
            .DOUT(N__8293),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__8295),
            .PADOUT(N__8294),
            .PADIN(N__8293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4341),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__3803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__8286),
            .DIN(N__8285),
            .DOUT(N__8284),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8286),
            .PADOUT(N__8285),
            .PADIN(N__8284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4321),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__2924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__8277),
            .DIN(N__8276),
            .DOUT(N__8275),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__8277),
            .PADOUT(N__8276),
            .PADIN(N__8275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4574),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__4868),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__8268),
            .DIN(N__8267),
            .DOUT(N__8266),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__8268),
            .PADOUT(N__8267),
            .PADIN(N__8266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4320),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__3857),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__8259),
            .DIN(N__8258),
            .DOUT(N__8257),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__8259),
            .PADOUT(N__8258),
            .PADIN(N__8257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5572),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__8250),
            .DIN(N__8249),
            .DOUT(N__8248),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__8250),
            .PADOUT(N__8249),
            .PADIN(N__8248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4750),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__2690),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__8241),
            .DIN(N__8240),
            .DOUT(N__8239),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__8241),
            .PADOUT(N__8240),
            .PADIN(N__8239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4636),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__3383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_obuf_iopad (
            .OE(N__8232),
            .DIN(N__8231),
            .DOUT(N__8230),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__8232),
            .PADOUT(N__8231),
            .PADIN(N__8230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4394),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__8223),
            .DIN(N__8222),
            .DOUT(N__8221),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__8223),
            .PADOUT(N__8222),
            .PADIN(N__8221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4302),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__5672),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__8214),
            .DIN(N__8213),
            .DOUT(N__8212),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__8214),
            .PADOUT(N__8213),
            .PADIN(N__8212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4322),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__3089),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__8205),
            .DIN(N__8204),
            .DOUT(N__8203),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__8205),
            .PADOUT(N__8204),
            .PADIN(N__8203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__8196),
            .DIN(N__8195),
            .DOUT(N__8194),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__8196),
            .PADOUT(N__8195),
            .PADIN(N__8194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__8187),
            .DIN(N__8186),
            .DOUT(N__8185),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__8187),
            .PADOUT(N__8186),
            .PADIN(N__8185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4674),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__2567),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__8178),
            .DIN(N__8177),
            .DOUT(N__8176),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__8178),
            .PADOUT(N__8177),
            .PADIN(N__8176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4584),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__5843),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__8169),
            .DIN(N__8168),
            .DOUT(N__8167),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__8169),
            .PADOUT(N__8168),
            .PADIN(N__8167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__8160),
            .DIN(N__8159),
            .DOUT(N__8158),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__8160),
            .PADOUT(N__8159),
            .PADIN(N__8158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4245),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__2843),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__8151),
            .DIN(N__8150),
            .DOUT(N__8149),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__8151),
            .PADOUT(N__8150),
            .PADIN(N__8149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3983),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__8142),
            .DIN(N__8141),
            .DOUT(N__8140),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__8142),
            .PADOUT(N__8141),
            .PADIN(N__8140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4649),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__3413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__8133),
            .DIN(N__8132),
            .DOUT(N__8131),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__8133),
            .PADOUT(N__8132),
            .PADIN(N__8131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4376),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__2963),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__8124),
            .DIN(N__8123),
            .DOUT(N__8122),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__8124),
            .PADOUT(N__8123),
            .PADIN(N__8122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4353),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__3512),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__8115),
            .DIN(N__8114),
            .DOUT(N__8113),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__8115),
            .PADOUT(N__8114),
            .PADIN(N__8113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4659),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__5150),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__8106),
            .DIN(N__8105),
            .DOUT(N__8104),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__8106),
            .PADOUT(N__8105),
            .PADIN(N__8104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__8097),
            .DIN(N__8096),
            .DOUT(N__8095),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__8097),
            .PADOUT(N__8096),
            .PADIN(N__8095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4751),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__2762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__8088),
            .DIN(N__8087),
            .DOUT(N__8086),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__8088),
            .PADOUT(N__8087),
            .PADIN(N__8086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4258),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__4013),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__8079),
            .DIN(N__8078),
            .DOUT(N__8077),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__8079),
            .PADOUT(N__8078),
            .PADIN(N__8077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4658),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__4898),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__8070),
            .DIN(N__8069),
            .DOUT(N__8068),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__8070),
            .PADOUT(N__8069),
            .PADIN(N__8068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__8061),
            .DIN(N__8060),
            .DOUT(N__8059),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__8061),
            .PADOUT(N__8060),
            .PADIN(N__8059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__8052),
            .DIN(N__8051),
            .DOUT(N__8050),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8052),
            .PADOUT(N__8051),
            .PADIN(N__8050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4339),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__3473),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__8043),
            .DIN(N__8042),
            .DOUT(N__8041),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__8043),
            .PADOUT(N__8042),
            .PADIN(N__8041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__8034),
            .DIN(N__8033),
            .DOUT(N__8032),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__8034),
            .PADOUT(N__8033),
            .PADIN(N__8032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__8025),
            .DIN(N__8024),
            .DOUT(N__8023),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__8025),
            .PADOUT(N__8024),
            .PADIN(N__8023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4592),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__3002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__8016),
            .DIN(N__8015),
            .DOUT(N__8014),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__8016),
            .PADOUT(N__8015),
            .PADIN(N__8014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4279),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__7001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__8007),
            .DIN(N__8006),
            .DOUT(N__8005),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__8007),
            .PADOUT(N__8006),
            .PADIN(N__8005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4639),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__3134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__7998),
            .DIN(N__7997),
            .DOUT(N__7996),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__7998),
            .PADOUT(N__7997),
            .PADIN(N__7996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4661),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__4796),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__7989),
            .DIN(N__7988),
            .DOUT(N__7987),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__7989),
            .PADOUT(N__7988),
            .PADIN(N__7987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4374),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__5960),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__7980),
            .DIN(N__7979),
            .DOUT(N__7978),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__7980),
            .PADOUT(N__7979),
            .PADIN(N__7978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4255),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__6593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2033 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__2032 (
            .O(N__7958),
            .I(N__7955));
    Sp12to4 I__2031 (
            .O(N__7955),
            .I(N__7952));
    Span12Mux_v I__2030 (
            .O(N__7952),
            .I(N__7949));
    Span12Mux_h I__2029 (
            .O(N__7949),
            .I(N__7946));
    Odrv12 I__2028 (
            .O(N__7946),
            .I(D_UU_040_in_5));
    IoInMux I__2027 (
            .O(N__7943),
            .I(N__7940));
    LocalMux I__2026 (
            .O(N__7940),
            .I(N__7937));
    Span4Mux_s3_h I__2025 (
            .O(N__7937),
            .I(N__7934));
    Span4Mux_v I__2024 (
            .O(N__7934),
            .I(N__7931));
    Sp12to4 I__2023 (
            .O(N__7931),
            .I(N__7928));
    Span12Mux_s9_h I__2022 (
            .O(N__7928),
            .I(N__7925));
    Odrv12 I__2021 (
            .O(N__7925),
            .I(un1_D_UU_040_5));
    InMux I__2020 (
            .O(N__7922),
            .I(N__7918));
    InMux I__2019 (
            .O(N__7921),
            .I(N__7912));
    LocalMux I__2018 (
            .O(N__7918),
            .I(N__7909));
    InMux I__2017 (
            .O(N__7917),
            .I(N__7904));
    InMux I__2016 (
            .O(N__7916),
            .I(N__7904));
    InMux I__2015 (
            .O(N__7915),
            .I(N__7901));
    LocalMux I__2014 (
            .O(N__7912),
            .I(N__7898));
    Span4Mux_v I__2013 (
            .O(N__7909),
            .I(N__7891));
    LocalMux I__2012 (
            .O(N__7904),
            .I(N__7891));
    LocalMux I__2011 (
            .O(N__7901),
            .I(N__7891));
    Span4Mux_h I__2010 (
            .O(N__7898),
            .I(N__7886));
    Span4Mux_h I__2009 (
            .O(N__7891),
            .I(N__7886));
    Sp12to4 I__2008 (
            .O(N__7886),
            .I(N__7883));
    Span12Mux_v I__2007 (
            .O(N__7883),
            .I(N__7880));
    Odrv12 I__2006 (
            .O(N__7880),
            .I(TS_CPUn_c));
    IoInMux I__2005 (
            .O(N__7877),
            .I(N__7874));
    LocalMux I__2004 (
            .O(N__7874),
            .I(N__7869));
    CascadeMux I__2003 (
            .O(N__7873),
            .I(N__7866));
    CascadeMux I__2002 (
            .O(N__7872),
            .I(N__7863));
    Span4Mux_s3_v I__2001 (
            .O(N__7869),
            .I(N__7860));
    InMux I__2000 (
            .O(N__7866),
            .I(N__7857));
    InMux I__1999 (
            .O(N__7863),
            .I(N__7854));
    Span4Mux_v I__1998 (
            .O(N__7860),
            .I(N__7851));
    LocalMux I__1997 (
            .O(N__7857),
            .I(N__7848));
    LocalMux I__1996 (
            .O(N__7854),
            .I(N__7845));
    Span4Mux_v I__1995 (
            .O(N__7851),
            .I(N__7842));
    Span4Mux_h I__1994 (
            .O(N__7848),
            .I(N__7839));
    Span4Mux_v I__1993 (
            .O(N__7845),
            .I(N__7836));
    Sp12to4 I__1992 (
            .O(N__7842),
            .I(N__7833));
    Span4Mux_v I__1991 (
            .O(N__7839),
            .I(N__7830));
    Sp12to4 I__1990 (
            .O(N__7836),
            .I(N__7827));
    Span12Mux_h I__1989 (
            .O(N__7833),
            .I(N__7822));
    Sp12to4 I__1988 (
            .O(N__7830),
            .I(N__7822));
    Span12Mux_h I__1987 (
            .O(N__7827),
            .I(N__7819));
    Span12Mux_h I__1986 (
            .O(N__7822),
            .I(N__7816));
    Odrv12 I__1985 (
            .O(N__7819),
            .I(RnW_c));
    Odrv12 I__1984 (
            .O(N__7816),
            .I(RnW_c));
    InMux I__1983 (
            .O(N__7811),
            .I(N__7802));
    InMux I__1982 (
            .O(N__7810),
            .I(N__7799));
    InMux I__1981 (
            .O(N__7809),
            .I(N__7796));
    InMux I__1980 (
            .O(N__7808),
            .I(N__7791));
    InMux I__1979 (
            .O(N__7807),
            .I(N__7791));
    InMux I__1978 (
            .O(N__7806),
            .I(N__7786));
    InMux I__1977 (
            .O(N__7805),
            .I(N__7786));
    LocalMux I__1976 (
            .O(N__7802),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1975 (
            .O(N__7799),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1974 (
            .O(N__7796),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1973 (
            .O(N__7791),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1972 (
            .O(N__7786),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1971 (
            .O(N__7775),
            .I(N__7772));
    LocalMux I__1970 (
            .O(N__7772),
            .I(N__7769));
    Span4Mux_v I__1969 (
            .O(N__7769),
            .I(N__7765));
    InMux I__1968 (
            .O(N__7768),
            .I(N__7762));
    Odrv4 I__1967 (
            .O(N__7765),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    LocalMux I__1966 (
            .O(N__7762),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    InMux I__1965 (
            .O(N__7757),
            .I(N__7754));
    LocalMux I__1964 (
            .O(N__7754),
            .I(N__7745));
    ClkMux I__1963 (
            .O(N__7753),
            .I(N__7703));
    ClkMux I__1962 (
            .O(N__7752),
            .I(N__7703));
    ClkMux I__1961 (
            .O(N__7751),
            .I(N__7703));
    ClkMux I__1960 (
            .O(N__7750),
            .I(N__7703));
    ClkMux I__1959 (
            .O(N__7749),
            .I(N__7703));
    ClkMux I__1958 (
            .O(N__7748),
            .I(N__7703));
    Glb2LocalMux I__1957 (
            .O(N__7745),
            .I(N__7703));
    ClkMux I__1956 (
            .O(N__7744),
            .I(N__7703));
    ClkMux I__1955 (
            .O(N__7743),
            .I(N__7703));
    ClkMux I__1954 (
            .O(N__7742),
            .I(N__7703));
    ClkMux I__1953 (
            .O(N__7741),
            .I(N__7703));
    ClkMux I__1952 (
            .O(N__7740),
            .I(N__7703));
    ClkMux I__1951 (
            .O(N__7739),
            .I(N__7703));
    ClkMux I__1950 (
            .O(N__7738),
            .I(N__7703));
    ClkMux I__1949 (
            .O(N__7737),
            .I(N__7703));
    ClkMux I__1948 (
            .O(N__7736),
            .I(N__7703));
    GlobalMux I__1947 (
            .O(N__7703),
            .I(CLK40));
    SRMux I__1946 (
            .O(N__7700),
            .I(N__7696));
    SRMux I__1945 (
            .O(N__7699),
            .I(N__7692));
    LocalMux I__1944 (
            .O(N__7696),
            .I(N__7688));
    SRMux I__1943 (
            .O(N__7695),
            .I(N__7685));
    LocalMux I__1942 (
            .O(N__7692),
            .I(N__7681));
    SRMux I__1941 (
            .O(N__7691),
            .I(N__7678));
    Span4Mux_h I__1940 (
            .O(N__7688),
            .I(N__7673));
    LocalMux I__1939 (
            .O(N__7685),
            .I(N__7673));
    SRMux I__1938 (
            .O(N__7684),
            .I(N__7670));
    Span4Mux_h I__1937 (
            .O(N__7681),
            .I(N__7665));
    LocalMux I__1936 (
            .O(N__7678),
            .I(N__7665));
    Span4Mux_h I__1935 (
            .O(N__7673),
            .I(N__7662));
    LocalMux I__1934 (
            .O(N__7670),
            .I(N__7659));
    Span4Mux_v I__1933 (
            .O(N__7665),
            .I(N__7656));
    Odrv4 I__1932 (
            .O(N__7662),
            .I(RESETn_c_i));
    Odrv12 I__1931 (
            .O(N__7659),
            .I(RESETn_c_i));
    Odrv4 I__1930 (
            .O(N__7656),
            .I(RESETn_c_i));
    InMux I__1929 (
            .O(N__7649),
            .I(N__7645));
    InMux I__1928 (
            .O(N__7648),
            .I(N__7642));
    LocalMux I__1927 (
            .O(N__7645),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    LocalMux I__1926 (
            .O(N__7642),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    InMux I__1925 (
            .O(N__7637),
            .I(N__7630));
    InMux I__1924 (
            .O(N__7636),
            .I(N__7630));
    InMux I__1923 (
            .O(N__7635),
            .I(N__7627));
    LocalMux I__1922 (
            .O(N__7630),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1921 (
            .O(N__7627),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    CascadeMux I__1920 (
            .O(N__7622),
            .I(N__7619));
    InMux I__1919 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__1918 (
            .O(N__7616),
            .I(N__7613));
    Span4Mux_v I__1917 (
            .O(N__7613),
            .I(N__7610));
    Span4Mux_h I__1916 (
            .O(N__7610),
            .I(N__7606));
    IoInMux I__1915 (
            .O(N__7609),
            .I(N__7603));
    Sp12to4 I__1914 (
            .O(N__7606),
            .I(N__7600));
    LocalMux I__1913 (
            .O(N__7603),
            .I(N__7597));
    Span12Mux_v I__1912 (
            .O(N__7600),
            .I(N__7594));
    IoSpan4Mux I__1911 (
            .O(N__7597),
            .I(N__7591));
    Odrv12 I__1910 (
            .O(N__7594),
            .I(TBIn_c));
    Odrv4 I__1909 (
            .O(N__7591),
            .I(TBIn_c));
    InMux I__1908 (
            .O(N__7586),
            .I(N__7579));
    InMux I__1907 (
            .O(N__7585),
            .I(N__7574));
    InMux I__1906 (
            .O(N__7584),
            .I(N__7574));
    InMux I__1905 (
            .O(N__7583),
            .I(N__7571));
    InMux I__1904 (
            .O(N__7582),
            .I(N__7568));
    LocalMux I__1903 (
            .O(N__7579),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1902 (
            .O(N__7574),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1901 (
            .O(N__7571),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1900 (
            .O(N__7568),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    InMux I__1899 (
            .O(N__7559),
            .I(N__7556));
    LocalMux I__1898 (
            .O(N__7556),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ));
    IoInMux I__1897 (
            .O(N__7553),
            .I(N__7549));
    CascadeMux I__1896 (
            .O(N__7552),
            .I(N__7545));
    LocalMux I__1895 (
            .O(N__7549),
            .I(N__7538));
    InMux I__1894 (
            .O(N__7548),
            .I(N__7535));
    InMux I__1893 (
            .O(N__7545),
            .I(N__7532));
    InMux I__1892 (
            .O(N__7544),
            .I(N__7529));
    InMux I__1891 (
            .O(N__7543),
            .I(N__7526));
    InMux I__1890 (
            .O(N__7542),
            .I(N__7521));
    InMux I__1889 (
            .O(N__7541),
            .I(N__7521));
    Span4Mux_s1_v I__1888 (
            .O(N__7538),
            .I(N__7518));
    LocalMux I__1887 (
            .O(N__7535),
            .I(N__7515));
    LocalMux I__1886 (
            .O(N__7532),
            .I(N__7506));
    LocalMux I__1885 (
            .O(N__7529),
            .I(N__7506));
    LocalMux I__1884 (
            .O(N__7526),
            .I(N__7506));
    LocalMux I__1883 (
            .O(N__7521),
            .I(N__7506));
    Sp12to4 I__1882 (
            .O(N__7518),
            .I(N__7503));
    Span4Mux_v I__1881 (
            .O(N__7515),
            .I(N__7500));
    Span4Mux_v I__1880 (
            .O(N__7506),
            .I(N__7497));
    Span12Mux_h I__1879 (
            .O(N__7503),
            .I(N__7493));
    Sp12to4 I__1878 (
            .O(N__7500),
            .I(N__7488));
    Sp12to4 I__1877 (
            .O(N__7497),
            .I(N__7488));
    InMux I__1876 (
            .O(N__7496),
            .I(N__7485));
    Span12Mux_v I__1875 (
            .O(N__7493),
            .I(N__7478));
    Span12Mux_h I__1874 (
            .O(N__7488),
            .I(N__7478));
    LocalMux I__1873 (
            .O(N__7485),
            .I(N__7478));
    Span12Mux_v I__1872 (
            .O(N__7478),
            .I(N__7475));
    Odrv12 I__1871 (
            .O(N__7475),
            .I(TACKn_in));
    InMux I__1870 (
            .O(N__7472),
            .I(N__7466));
    InMux I__1869 (
            .O(N__7471),
            .I(N__7463));
    InMux I__1868 (
            .O(N__7470),
            .I(N__7460));
    InMux I__1867 (
            .O(N__7469),
            .I(N__7457));
    LocalMux I__1866 (
            .O(N__7466),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1865 (
            .O(N__7463),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1864 (
            .O(N__7460),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1863 (
            .O(N__7457),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    CascadeMux I__1862 (
            .O(N__7448),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ));
    InMux I__1861 (
            .O(N__7445),
            .I(N__7438));
    InMux I__1860 (
            .O(N__7444),
            .I(N__7435));
    InMux I__1859 (
            .O(N__7443),
            .I(N__7432));
    InMux I__1858 (
            .O(N__7442),
            .I(N__7427));
    InMux I__1857 (
            .O(N__7441),
            .I(N__7427));
    LocalMux I__1856 (
            .O(N__7438),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1855 (
            .O(N__7435),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1854 (
            .O(N__7432),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1853 (
            .O(N__7427),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    InMux I__1852 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__1851 (
            .O(N__7415),
            .I(\U111_CYCLE_SM.N_136 ));
    InMux I__1850 (
            .O(N__7412),
            .I(N__7409));
    LocalMux I__1849 (
            .O(N__7409),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    InMux I__1848 (
            .O(N__7406),
            .I(N__7403));
    LocalMux I__1847 (
            .O(N__7403),
            .I(N__7400));
    Span4Mux_v I__1846 (
            .O(N__7400),
            .I(N__7395));
    InMux I__1845 (
            .O(N__7399),
            .I(N__7392));
    InMux I__1844 (
            .O(N__7398),
            .I(N__7389));
    Span4Mux_v I__1843 (
            .O(N__7395),
            .I(N__7382));
    LocalMux I__1842 (
            .O(N__7392),
            .I(N__7382));
    LocalMux I__1841 (
            .O(N__7389),
            .I(N__7382));
    Span4Mux_v I__1840 (
            .O(N__7382),
            .I(N__7379));
    Sp12to4 I__1839 (
            .O(N__7379),
            .I(N__7376));
    Span12Mux_h I__1838 (
            .O(N__7376),
            .I(N__7373));
    Odrv12 I__1837 (
            .O(N__7373),
            .I(D_UM_AMIGA_in_2));
    IoInMux I__1836 (
            .O(N__7370),
            .I(N__7367));
    LocalMux I__1835 (
            .O(N__7367),
            .I(N__7364));
    IoSpan4Mux I__1834 (
            .O(N__7364),
            .I(N__7361));
    Span4Mux_s2_h I__1833 (
            .O(N__7361),
            .I(N__7358));
    Sp12to4 I__1832 (
            .O(N__7358),
            .I(N__7355));
    Odrv12 I__1831 (
            .O(N__7355),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1830 (
            .O(N__7352),
            .I(N__7349));
    LocalMux I__1829 (
            .O(N__7349),
            .I(N__7346));
    Sp12to4 I__1828 (
            .O(N__7346),
            .I(N__7343));
    Span12Mux_v I__1827 (
            .O(N__7343),
            .I(N__7340));
    Span12Mux_h I__1826 (
            .O(N__7340),
            .I(N__7337));
    Odrv12 I__1825 (
            .O(N__7337),
            .I(D_UM_040_in_1));
    IoInMux I__1824 (
            .O(N__7334),
            .I(N__7330));
    InMux I__1823 (
            .O(N__7333),
            .I(N__7327));
    LocalMux I__1822 (
            .O(N__7330),
            .I(N__7324));
    LocalMux I__1821 (
            .O(N__7327),
            .I(N__7321));
    Span4Mux_s3_h I__1820 (
            .O(N__7324),
            .I(N__7318));
    Span4Mux_h I__1819 (
            .O(N__7321),
            .I(N__7315));
    Sp12to4 I__1818 (
            .O(N__7318),
            .I(N__7312));
    Sp12to4 I__1817 (
            .O(N__7315),
            .I(N__7309));
    Span12Mux_v I__1816 (
            .O(N__7312),
            .I(N__7306));
    Span12Mux_v I__1815 (
            .O(N__7309),
            .I(N__7303));
    Span12Mux_h I__1814 (
            .O(N__7306),
            .I(N__7300));
    Span12Mux_v I__1813 (
            .O(N__7303),
            .I(N__7297));
    Span12Mux_h I__1812 (
            .O(N__7300),
            .I(N__7294));
    Span12Mux_h I__1811 (
            .O(N__7297),
            .I(N__7291));
    Odrv12 I__1810 (
            .O(N__7294),
            .I(D_LL_040_in_1));
    Odrv12 I__1809 (
            .O(N__7291),
            .I(D_LL_040_in_1));
    IoInMux I__1808 (
            .O(N__7286),
            .I(N__7283));
    LocalMux I__1807 (
            .O(N__7283),
            .I(N__7280));
    IoSpan4Mux I__1806 (
            .O(N__7280),
            .I(N__7277));
    Sp12to4 I__1805 (
            .O(N__7277),
            .I(N__7274));
    Span12Mux_h I__1804 (
            .O(N__7274),
            .I(N__7271));
    Odrv12 I__1803 (
            .O(N__7271),
            .I(un1_D_UM_040_1));
    InMux I__1802 (
            .O(N__7268),
            .I(N__7265));
    LocalMux I__1801 (
            .O(N__7265),
            .I(N__7260));
    InMux I__1800 (
            .O(N__7264),
            .I(N__7257));
    InMux I__1799 (
            .O(N__7263),
            .I(N__7254));
    Span4Mux_v I__1798 (
            .O(N__7260),
            .I(N__7251));
    LocalMux I__1797 (
            .O(N__7257),
            .I(N__7246));
    LocalMux I__1796 (
            .O(N__7254),
            .I(N__7246));
    Span4Mux_v I__1795 (
            .O(N__7251),
            .I(N__7243));
    Span4Mux_v I__1794 (
            .O(N__7246),
            .I(N__7240));
    Sp12to4 I__1793 (
            .O(N__7243),
            .I(N__7235));
    Sp12to4 I__1792 (
            .O(N__7240),
            .I(N__7235));
    Span12Mux_h I__1791 (
            .O(N__7235),
            .I(N__7232));
    Span12Mux_v I__1790 (
            .O(N__7232),
            .I(N__7229));
    Odrv12 I__1789 (
            .O(N__7229),
            .I(D_UM_AMIGA_in_6));
    InMux I__1788 (
            .O(N__7226),
            .I(N__7223));
    LocalMux I__1787 (
            .O(N__7223),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__1786 (
            .O(N__7220),
            .I(N__7213));
    InMux I__1785 (
            .O(N__7219),
            .I(N__7213));
    InMux I__1784 (
            .O(N__7218),
            .I(N__7210));
    LocalMux I__1783 (
            .O(N__7213),
            .I(N__7202));
    LocalMux I__1782 (
            .O(N__7210),
            .I(N__7202));
    InMux I__1781 (
            .O(N__7209),
            .I(N__7199));
    InMux I__1780 (
            .O(N__7208),
            .I(N__7194));
    InMux I__1779 (
            .O(N__7207),
            .I(N__7194));
    Span4Mux_v I__1778 (
            .O(N__7202),
            .I(N__7180));
    LocalMux I__1777 (
            .O(N__7199),
            .I(N__7180));
    LocalMux I__1776 (
            .O(N__7194),
            .I(N__7180));
    InMux I__1775 (
            .O(N__7193),
            .I(N__7173));
    InMux I__1774 (
            .O(N__7192),
            .I(N__7173));
    InMux I__1773 (
            .O(N__7191),
            .I(N__7173));
    InMux I__1772 (
            .O(N__7190),
            .I(N__7168));
    InMux I__1771 (
            .O(N__7189),
            .I(N__7165));
    InMux I__1770 (
            .O(N__7188),
            .I(N__7162));
    InMux I__1769 (
            .O(N__7187),
            .I(N__7159));
    Span4Mux_v I__1768 (
            .O(N__7180),
            .I(N__7155));
    LocalMux I__1767 (
            .O(N__7173),
            .I(N__7152));
    InMux I__1766 (
            .O(N__7172),
            .I(N__7147));
    InMux I__1765 (
            .O(N__7171),
            .I(N__7147));
    LocalMux I__1764 (
            .O(N__7168),
            .I(N__7142));
    LocalMux I__1763 (
            .O(N__7165),
            .I(N__7142));
    LocalMux I__1762 (
            .O(N__7162),
            .I(N__7137));
    LocalMux I__1761 (
            .O(N__7159),
            .I(N__7137));
    CascadeMux I__1760 (
            .O(N__7158),
            .I(N__7133));
    Span4Mux_v I__1759 (
            .O(N__7155),
            .I(N__7130));
    Span12Mux_s8_v I__1758 (
            .O(N__7152),
            .I(N__7125));
    LocalMux I__1757 (
            .O(N__7147),
            .I(N__7125));
    Span4Mux_v I__1756 (
            .O(N__7142),
            .I(N__7120));
    Span4Mux_v I__1755 (
            .O(N__7137),
            .I(N__7120));
    InMux I__1754 (
            .O(N__7136),
            .I(N__7117));
    InMux I__1753 (
            .O(N__7133),
            .I(N__7114));
    Odrv4 I__1752 (
            .O(N__7130),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv12 I__1751 (
            .O(N__7125),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__1750 (
            .O(N__7120),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1749 (
            .O(N__7117),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1748 (
            .O(N__7114),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    IoInMux I__1747 (
            .O(N__7103),
            .I(N__7100));
    LocalMux I__1746 (
            .O(N__7100),
            .I(N__7097));
    IoSpan4Mux I__1745 (
            .O(N__7097),
            .I(N__7094));
    Span4Mux_s3_h I__1744 (
            .O(N__7094),
            .I(N__7091));
    Span4Mux_h I__1743 (
            .O(N__7091),
            .I(N__7088));
    Span4Mux_h I__1742 (
            .O(N__7088),
            .I(N__7085));
    Odrv4 I__1741 (
            .O(N__7085),
            .I(un1_D_UM_AMIGA_6));
    InMux I__1740 (
            .O(N__7082),
            .I(N__7079));
    LocalMux I__1739 (
            .O(N__7079),
            .I(N__7076));
    Span12Mux_v I__1738 (
            .O(N__7076),
            .I(N__7073));
    Span12Mux_h I__1737 (
            .O(N__7073),
            .I(N__7070));
    Odrv12 I__1736 (
            .O(N__7070),
            .I(D_UU_040_in_6));
    IoInMux I__1735 (
            .O(N__7067),
            .I(N__7064));
    LocalMux I__1734 (
            .O(N__7064),
            .I(N__7061));
    Span4Mux_s2_h I__1733 (
            .O(N__7061),
            .I(N__7057));
    InMux I__1732 (
            .O(N__7060),
            .I(N__7054));
    Span4Mux_v I__1731 (
            .O(N__7057),
            .I(N__7051));
    LocalMux I__1730 (
            .O(N__7054),
            .I(N__7048));
    Sp12to4 I__1729 (
            .O(N__7051),
            .I(N__7045));
    Sp12to4 I__1728 (
            .O(N__7048),
            .I(N__7042));
    Span12Mux_h I__1727 (
            .O(N__7045),
            .I(N__7039));
    Span12Mux_s11_v I__1726 (
            .O(N__7042),
            .I(N__7036));
    Span12Mux_h I__1725 (
            .O(N__7039),
            .I(N__7033));
    Span12Mux_h I__1724 (
            .O(N__7036),
            .I(N__7030));
    Odrv12 I__1723 (
            .O(N__7033),
            .I(D_LM_040_in_6));
    Odrv12 I__1722 (
            .O(N__7030),
            .I(D_LM_040_in_6));
    IoInMux I__1721 (
            .O(N__7025),
            .I(N__7022));
    LocalMux I__1720 (
            .O(N__7022),
            .I(N__7019));
    IoSpan4Mux I__1719 (
            .O(N__7019),
            .I(N__7016));
    IoSpan4Mux I__1718 (
            .O(N__7016),
            .I(N__7013));
    Span4Mux_s2_v I__1717 (
            .O(N__7013),
            .I(N__7010));
    Span4Mux_h I__1716 (
            .O(N__7010),
            .I(N__7007));
    Span4Mux_v I__1715 (
            .O(N__7007),
            .I(N__7004));
    Odrv4 I__1714 (
            .O(N__7004),
            .I(un1_D_UU_040_6));
    IoInMux I__1713 (
            .O(N__7001),
            .I(N__6998));
    LocalMux I__1712 (
            .O(N__6998),
            .I(N__6995));
    IoSpan4Mux I__1711 (
            .O(N__6995),
            .I(N__6992));
    Span4Mux_s2_h I__1710 (
            .O(N__6992),
            .I(N__6988));
    InMux I__1709 (
            .O(N__6991),
            .I(N__6985));
    Span4Mux_v I__1708 (
            .O(N__6988),
            .I(N__6982));
    LocalMux I__1707 (
            .O(N__6985),
            .I(N__6979));
    Sp12to4 I__1706 (
            .O(N__6982),
            .I(N__6976));
    Sp12to4 I__1705 (
            .O(N__6979),
            .I(N__6973));
    Span12Mux_s9_h I__1704 (
            .O(N__6976),
            .I(N__6970));
    Span12Mux_v I__1703 (
            .O(N__6973),
            .I(N__6967));
    Span12Mux_h I__1702 (
            .O(N__6970),
            .I(N__6964));
    Span12Mux_h I__1701 (
            .O(N__6967),
            .I(N__6961));
    Odrv12 I__1700 (
            .O(N__6964),
            .I(D_LM_040_in_5));
    Odrv12 I__1699 (
            .O(N__6961),
            .I(D_LM_040_in_5));
    InMux I__1698 (
            .O(N__6956),
            .I(N__6950));
    InMux I__1697 (
            .O(N__6955),
            .I(N__6950));
    LocalMux I__1696 (
            .O(N__6950),
            .I(N__6941));
    InMux I__1695 (
            .O(N__6949),
            .I(N__6938));
    InMux I__1694 (
            .O(N__6948),
            .I(N__6927));
    InMux I__1693 (
            .O(N__6947),
            .I(N__6927));
    InMux I__1692 (
            .O(N__6946),
            .I(N__6922));
    InMux I__1691 (
            .O(N__6945),
            .I(N__6922));
    InMux I__1690 (
            .O(N__6944),
            .I(N__6912));
    Span4Mux_v I__1689 (
            .O(N__6941),
            .I(N__6907));
    LocalMux I__1688 (
            .O(N__6938),
            .I(N__6907));
    InMux I__1687 (
            .O(N__6937),
            .I(N__6900));
    InMux I__1686 (
            .O(N__6936),
            .I(N__6900));
    InMux I__1685 (
            .O(N__6935),
            .I(N__6900));
    InMux I__1684 (
            .O(N__6934),
            .I(N__6895));
    InMux I__1683 (
            .O(N__6933),
            .I(N__6890));
    InMux I__1682 (
            .O(N__6932),
            .I(N__6890));
    LocalMux I__1681 (
            .O(N__6927),
            .I(N__6885));
    LocalMux I__1680 (
            .O(N__6922),
            .I(N__6885));
    InMux I__1679 (
            .O(N__6921),
            .I(N__6882));
    InMux I__1678 (
            .O(N__6920),
            .I(N__6877));
    InMux I__1677 (
            .O(N__6919),
            .I(N__6870));
    InMux I__1676 (
            .O(N__6918),
            .I(N__6870));
    InMux I__1675 (
            .O(N__6917),
            .I(N__6870));
    InMux I__1674 (
            .O(N__6916),
            .I(N__6865));
    InMux I__1673 (
            .O(N__6915),
            .I(N__6865));
    LocalMux I__1672 (
            .O(N__6912),
            .I(N__6858));
    Span4Mux_h I__1671 (
            .O(N__6907),
            .I(N__6858));
    LocalMux I__1670 (
            .O(N__6900),
            .I(N__6858));
    InMux I__1669 (
            .O(N__6899),
            .I(N__6855));
    InMux I__1668 (
            .O(N__6898),
            .I(N__6852));
    LocalMux I__1667 (
            .O(N__6895),
            .I(N__6847));
    LocalMux I__1666 (
            .O(N__6890),
            .I(N__6847));
    Span4Mux_v I__1665 (
            .O(N__6885),
            .I(N__6843));
    LocalMux I__1664 (
            .O(N__6882),
            .I(N__6840));
    InMux I__1663 (
            .O(N__6881),
            .I(N__6835));
    InMux I__1662 (
            .O(N__6880),
            .I(N__6835));
    LocalMux I__1661 (
            .O(N__6877),
            .I(N__6828));
    LocalMux I__1660 (
            .O(N__6870),
            .I(N__6825));
    LocalMux I__1659 (
            .O(N__6865),
            .I(N__6822));
    Span4Mux_v I__1658 (
            .O(N__6858),
            .I(N__6815));
    LocalMux I__1657 (
            .O(N__6855),
            .I(N__6815));
    LocalMux I__1656 (
            .O(N__6852),
            .I(N__6815));
    Span4Mux_v I__1655 (
            .O(N__6847),
            .I(N__6812));
    InMux I__1654 (
            .O(N__6846),
            .I(N__6809));
    Span4Mux_v I__1653 (
            .O(N__6843),
            .I(N__6802));
    Span4Mux_h I__1652 (
            .O(N__6840),
            .I(N__6802));
    LocalMux I__1651 (
            .O(N__6835),
            .I(N__6802));
    InMux I__1650 (
            .O(N__6834),
            .I(N__6797));
    InMux I__1649 (
            .O(N__6833),
            .I(N__6797));
    InMux I__1648 (
            .O(N__6832),
            .I(N__6792));
    InMux I__1647 (
            .O(N__6831),
            .I(N__6792));
    Span12Mux_v I__1646 (
            .O(N__6828),
            .I(N__6784));
    Span12Mux_v I__1645 (
            .O(N__6825),
            .I(N__6784));
    Span12Mux_v I__1644 (
            .O(N__6822),
            .I(N__6781));
    Span4Mux_v I__1643 (
            .O(N__6815),
            .I(N__6778));
    Span4Mux_v I__1642 (
            .O(N__6812),
            .I(N__6773));
    LocalMux I__1641 (
            .O(N__6809),
            .I(N__6773));
    Span4Mux_v I__1640 (
            .O(N__6802),
            .I(N__6770));
    LocalMux I__1639 (
            .O(N__6797),
            .I(N__6765));
    LocalMux I__1638 (
            .O(N__6792),
            .I(N__6765));
    InMux I__1637 (
            .O(N__6791),
            .I(N__6762));
    InMux I__1636 (
            .O(N__6790),
            .I(N__6759));
    InMux I__1635 (
            .O(N__6789),
            .I(N__6756));
    Odrv12 I__1634 (
            .O(N__6784),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1633 (
            .O(N__6781),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1632 (
            .O(N__6778),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1631 (
            .O(N__6773),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1630 (
            .O(N__6770),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1629 (
            .O(N__6765),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1628 (
            .O(N__6762),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1627 (
            .O(N__6759),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1626 (
            .O(N__6756),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    InMux I__1625 (
            .O(N__6737),
            .I(N__6734));
    LocalMux I__1624 (
            .O(N__6734),
            .I(N__6731));
    Odrv12 I__1623 (
            .O(N__6731),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1622 (
            .O(N__6728),
            .I(N__6724));
    InMux I__1621 (
            .O(N__6727),
            .I(N__6721));
    LocalMux I__1620 (
            .O(N__6724),
            .I(N__6718));
    LocalMux I__1619 (
            .O(N__6721),
            .I(N__6714));
    Span4Mux_v I__1618 (
            .O(N__6718),
            .I(N__6711));
    InMux I__1617 (
            .O(N__6717),
            .I(N__6708));
    Span4Mux_v I__1616 (
            .O(N__6714),
            .I(N__6705));
    Span4Mux_v I__1615 (
            .O(N__6711),
            .I(N__6700));
    LocalMux I__1614 (
            .O(N__6708),
            .I(N__6700));
    Span4Mux_v I__1613 (
            .O(N__6705),
            .I(N__6695));
    Span4Mux_h I__1612 (
            .O(N__6700),
            .I(N__6695));
    Span4Mux_v I__1611 (
            .O(N__6695),
            .I(N__6692));
    Sp12to4 I__1610 (
            .O(N__6692),
            .I(N__6689));
    Span12Mux_h I__1609 (
            .O(N__6689),
            .I(N__6686));
    Odrv12 I__1608 (
            .O(N__6686),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1607 (
            .O(N__6683),
            .I(N__6680));
    LocalMux I__1606 (
            .O(N__6680),
            .I(N__6677));
    IoSpan4Mux I__1605 (
            .O(N__6677),
            .I(N__6674));
    IoSpan4Mux I__1604 (
            .O(N__6674),
            .I(N__6671));
    Sp12to4 I__1603 (
            .O(N__6671),
            .I(N__6668));
    Span12Mux_s6_v I__1602 (
            .O(N__6668),
            .I(N__6665));
    Odrv12 I__1601 (
            .O(N__6665),
            .I(un1_D_UU_AMIGA_5));
    IoInMux I__1600 (
            .O(N__6662),
            .I(N__6659));
    LocalMux I__1599 (
            .O(N__6659),
            .I(N__6656));
    IoSpan4Mux I__1598 (
            .O(N__6656),
            .I(N__6652));
    InMux I__1597 (
            .O(N__6655),
            .I(N__6649));
    IoSpan4Mux I__1596 (
            .O(N__6652),
            .I(N__6646));
    LocalMux I__1595 (
            .O(N__6649),
            .I(N__6643));
    Span4Mux_s2_h I__1594 (
            .O(N__6646),
            .I(N__6640));
    Span4Mux_v I__1593 (
            .O(N__6643),
            .I(N__6637));
    Sp12to4 I__1592 (
            .O(N__6640),
            .I(N__6634));
    Sp12to4 I__1591 (
            .O(N__6637),
            .I(N__6631));
    Span12Mux_h I__1590 (
            .O(N__6634),
            .I(N__6628));
    Span12Mux_h I__1589 (
            .O(N__6631),
            .I(N__6625));
    Span12Mux_h I__1588 (
            .O(N__6628),
            .I(N__6622));
    Span12Mux_v I__1587 (
            .O(N__6625),
            .I(N__6619));
    Odrv12 I__1586 (
            .O(N__6622),
            .I(D_LM_040_in_3));
    Odrv12 I__1585 (
            .O(N__6619),
            .I(D_LM_040_in_3));
    InMux I__1584 (
            .O(N__6614),
            .I(N__6611));
    LocalMux I__1583 (
            .O(N__6611),
            .I(N__6608));
    Span4Mux_v I__1582 (
            .O(N__6608),
            .I(N__6605));
    Span4Mux_h I__1581 (
            .O(N__6605),
            .I(N__6602));
    Sp12to4 I__1580 (
            .O(N__6602),
            .I(N__6599));
    Span12Mux_h I__1579 (
            .O(N__6599),
            .I(N__6596));
    Odrv12 I__1578 (
            .O(N__6596),
            .I(D_UU_040_in_3));
    IoInMux I__1577 (
            .O(N__6593),
            .I(N__6590));
    LocalMux I__1576 (
            .O(N__6590),
            .I(N__6587));
    Span4Mux_s2_v I__1575 (
            .O(N__6587),
            .I(N__6584));
    Span4Mux_v I__1574 (
            .O(N__6584),
            .I(N__6581));
    Sp12to4 I__1573 (
            .O(N__6581),
            .I(N__6578));
    Span12Mux_h I__1572 (
            .O(N__6578),
            .I(N__6575));
    Odrv12 I__1571 (
            .O(N__6575),
            .I(un1_D_UU_040_3));
    InMux I__1570 (
            .O(N__6572),
            .I(N__6569));
    LocalMux I__1569 (
            .O(N__6569),
            .I(N__6566));
    Odrv12 I__1568 (
            .O(N__6566),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    InMux I__1567 (
            .O(N__6563),
            .I(N__6559));
    InMux I__1566 (
            .O(N__6562),
            .I(N__6556));
    LocalMux I__1565 (
            .O(N__6559),
            .I(N__6553));
    LocalMux I__1564 (
            .O(N__6556),
            .I(N__6550));
    Span4Mux_v I__1563 (
            .O(N__6553),
            .I(N__6546));
    Span4Mux_v I__1562 (
            .O(N__6550),
            .I(N__6543));
    InMux I__1561 (
            .O(N__6549),
            .I(N__6540));
    Span4Mux_v I__1560 (
            .O(N__6546),
            .I(N__6537));
    Span4Mux_v I__1559 (
            .O(N__6543),
            .I(N__6532));
    LocalMux I__1558 (
            .O(N__6540),
            .I(N__6532));
    Span4Mux_v I__1557 (
            .O(N__6537),
            .I(N__6527));
    Span4Mux_v I__1556 (
            .O(N__6532),
            .I(N__6527));
    Sp12to4 I__1555 (
            .O(N__6527),
            .I(N__6524));
    Span12Mux_h I__1554 (
            .O(N__6524),
            .I(N__6521));
    Odrv12 I__1553 (
            .O(N__6521),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1552 (
            .O(N__6518),
            .I(N__6515));
    LocalMux I__1551 (
            .O(N__6515),
            .I(N__6512));
    IoSpan4Mux I__1550 (
            .O(N__6512),
            .I(N__6509));
    Sp12to4 I__1549 (
            .O(N__6509),
            .I(N__6506));
    Span12Mux_s6_v I__1548 (
            .O(N__6506),
            .I(N__6503));
    Odrv12 I__1547 (
            .O(N__6503),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1546 (
            .O(N__6500),
            .I(N__6495));
    InMux I__1545 (
            .O(N__6499),
            .I(N__6490));
    InMux I__1544 (
            .O(N__6498),
            .I(N__6490));
    LocalMux I__1543 (
            .O(N__6495),
            .I(N__6487));
    LocalMux I__1542 (
            .O(N__6490),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    Odrv4 I__1541 (
            .O(N__6487),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    CascadeMux I__1540 (
            .O(N__6482),
            .I(N__6478));
    InMux I__1539 (
            .O(N__6481),
            .I(N__6474));
    InMux I__1538 (
            .O(N__6478),
            .I(N__6471));
    InMux I__1537 (
            .O(N__6477),
            .I(N__6467));
    LocalMux I__1536 (
            .O(N__6474),
            .I(N__6464));
    LocalMux I__1535 (
            .O(N__6471),
            .I(N__6460));
    InMux I__1534 (
            .O(N__6470),
            .I(N__6457));
    LocalMux I__1533 (
            .O(N__6467),
            .I(N__6454));
    Span4Mux_h I__1532 (
            .O(N__6464),
            .I(N__6451));
    InMux I__1531 (
            .O(N__6463),
            .I(N__6448));
    Odrv4 I__1530 (
            .O(N__6460),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1529 (
            .O(N__6457),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    Odrv4 I__1528 (
            .O(N__6454),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    Odrv4 I__1527 (
            .O(N__6451),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1526 (
            .O(N__6448),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    InMux I__1525 (
            .O(N__6437),
            .I(N__6432));
    InMux I__1524 (
            .O(N__6436),
            .I(N__6429));
    InMux I__1523 (
            .O(N__6435),
            .I(N__6426));
    LocalMux I__1522 (
            .O(N__6432),
            .I(N__6421));
    LocalMux I__1521 (
            .O(N__6429),
            .I(N__6421));
    LocalMux I__1520 (
            .O(N__6426),
            .I(N__6418));
    Span12Mux_h I__1519 (
            .O(N__6421),
            .I(N__6415));
    Span12Mux_h I__1518 (
            .O(N__6418),
            .I(N__6412));
    Span12Mux_v I__1517 (
            .O(N__6415),
            .I(N__6409));
    Span12Mux_v I__1516 (
            .O(N__6412),
            .I(N__6406));
    Odrv12 I__1515 (
            .O(N__6409),
            .I(PORTSIZE_c));
    Odrv12 I__1514 (
            .O(N__6406),
            .I(PORTSIZE_c));
    CascadeMux I__1513 (
            .O(N__6401),
            .I(N__6398));
    InMux I__1512 (
            .O(N__6398),
            .I(N__6392));
    InMux I__1511 (
            .O(N__6397),
            .I(N__6392));
    LocalMux I__1510 (
            .O(N__6392),
            .I(N__6389));
    Span12Mux_h I__1509 (
            .O(N__6389),
            .I(N__6386));
    Span12Mux_v I__1508 (
            .O(N__6386),
            .I(N__6383));
    Odrv12 I__1507 (
            .O(N__6383),
            .I(SIZ_c_1));
    CascadeMux I__1506 (
            .O(N__6380),
            .I(N__6376));
    InMux I__1505 (
            .O(N__6379),
            .I(N__6371));
    InMux I__1504 (
            .O(N__6376),
            .I(N__6371));
    LocalMux I__1503 (
            .O(N__6371),
            .I(N__6368));
    Span12Mux_h I__1502 (
            .O(N__6368),
            .I(N__6365));
    Span12Mux_v I__1501 (
            .O(N__6365),
            .I(N__6362));
    Odrv12 I__1500 (
            .O(N__6362),
            .I(SIZ_c_0));
    CascadeMux I__1499 (
            .O(N__6359),
            .I(N__6354));
    InMux I__1498 (
            .O(N__6358),
            .I(N__6343));
    InMux I__1497 (
            .O(N__6357),
            .I(N__6343));
    InMux I__1496 (
            .O(N__6354),
            .I(N__6343));
    InMux I__1495 (
            .O(N__6353),
            .I(N__6343));
    InMux I__1494 (
            .O(N__6352),
            .I(N__6340));
    LocalMux I__1493 (
            .O(N__6343),
            .I(N__6337));
    LocalMux I__1492 (
            .O(N__6340),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    Odrv4 I__1491 (
            .O(N__6337),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    InMux I__1490 (
            .O(N__6332),
            .I(N__6323));
    InMux I__1489 (
            .O(N__6331),
            .I(N__6323));
    InMux I__1488 (
            .O(N__6330),
            .I(N__6320));
    InMux I__1487 (
            .O(N__6329),
            .I(N__6315));
    InMux I__1486 (
            .O(N__6328),
            .I(N__6315));
    LocalMux I__1485 (
            .O(N__6323),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    LocalMux I__1484 (
            .O(N__6320),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    LocalMux I__1483 (
            .O(N__6315),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    CEMux I__1482 (
            .O(N__6308),
            .I(N__6303));
    CEMux I__1481 (
            .O(N__6307),
            .I(N__6299));
    CEMux I__1480 (
            .O(N__6306),
            .I(N__6296));
    LocalMux I__1479 (
            .O(N__6303),
            .I(N__6292));
    CEMux I__1478 (
            .O(N__6302),
            .I(N__6289));
    LocalMux I__1477 (
            .O(N__6299),
            .I(N__6285));
    LocalMux I__1476 (
            .O(N__6296),
            .I(N__6282));
    CEMux I__1475 (
            .O(N__6295),
            .I(N__6279));
    Span4Mux_h I__1474 (
            .O(N__6292),
            .I(N__6274));
    LocalMux I__1473 (
            .O(N__6289),
            .I(N__6274));
    CEMux I__1472 (
            .O(N__6288),
            .I(N__6271));
    Span4Mux_v I__1471 (
            .O(N__6285),
            .I(N__6266));
    Span4Mux_v I__1470 (
            .O(N__6282),
            .I(N__6266));
    LocalMux I__1469 (
            .O(N__6279),
            .I(N__6263));
    Span4Mux_h I__1468 (
            .O(N__6274),
            .I(N__6260));
    LocalMux I__1467 (
            .O(N__6271),
            .I(N__6257));
    Odrv4 I__1466 (
            .O(N__6266),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1465 (
            .O(N__6263),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1464 (
            .O(N__6260),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1463 (
            .O(N__6257),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    SRMux I__1462 (
            .O(N__6248),
            .I(N__6240));
    SRMux I__1461 (
            .O(N__6247),
            .I(N__6237));
    SRMux I__1460 (
            .O(N__6246),
            .I(N__6234));
    SRMux I__1459 (
            .O(N__6245),
            .I(N__6231));
    SRMux I__1458 (
            .O(N__6244),
            .I(N__6228));
    SRMux I__1457 (
            .O(N__6243),
            .I(N__6225));
    LocalMux I__1456 (
            .O(N__6240),
            .I(N__6222));
    LocalMux I__1455 (
            .O(N__6237),
            .I(N__6215));
    LocalMux I__1454 (
            .O(N__6234),
            .I(N__6215));
    LocalMux I__1453 (
            .O(N__6231),
            .I(N__6215));
    LocalMux I__1452 (
            .O(N__6228),
            .I(N__6210));
    LocalMux I__1451 (
            .O(N__6225),
            .I(N__6210));
    Odrv4 I__1450 (
            .O(N__6222),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    Odrv4 I__1449 (
            .O(N__6215),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    Odrv4 I__1448 (
            .O(N__6210),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ));
    InMux I__1447 (
            .O(N__6203),
            .I(N__6200));
    LocalMux I__1446 (
            .O(N__6200),
            .I(N__6197));
    Span4Mux_v I__1445 (
            .O(N__6197),
            .I(N__6194));
    Span4Mux_v I__1444 (
            .O(N__6194),
            .I(N__6190));
    InMux I__1443 (
            .O(N__6193),
            .I(N__6187));
    Span4Mux_v I__1442 (
            .O(N__6190),
            .I(N__6181));
    LocalMux I__1441 (
            .O(N__6187),
            .I(N__6181));
    InMux I__1440 (
            .O(N__6186),
            .I(N__6178));
    Span4Mux_h I__1439 (
            .O(N__6181),
            .I(N__6173));
    LocalMux I__1438 (
            .O(N__6178),
            .I(N__6173));
    Span4Mux_v I__1437 (
            .O(N__6173),
            .I(N__6170));
    Span4Mux_v I__1436 (
            .O(N__6170),
            .I(N__6167));
    Sp12to4 I__1435 (
            .O(N__6167),
            .I(N__6164));
    Span12Mux_h I__1434 (
            .O(N__6164),
            .I(N__6161));
    Odrv12 I__1433 (
            .O(N__6161),
            .I(D_UM_AMIGA_in_4));
    InMux I__1432 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__1431 (
            .O(N__6155),
            .I(N__6152));
    Odrv4 I__1430 (
            .O(N__6152),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    IoInMux I__1429 (
            .O(N__6149),
            .I(N__6146));
    LocalMux I__1428 (
            .O(N__6146),
            .I(N__6143));
    IoSpan4Mux I__1427 (
            .O(N__6143),
            .I(N__6140));
    Sp12to4 I__1426 (
            .O(N__6140),
            .I(N__6137));
    Span12Mux_s6_v I__1425 (
            .O(N__6137),
            .I(N__6134));
    Span12Mux_h I__1424 (
            .O(N__6134),
            .I(N__6131));
    Odrv12 I__1423 (
            .O(N__6131),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1422 (
            .O(N__6128),
            .I(N__6125));
    LocalMux I__1421 (
            .O(N__6125),
            .I(N__6122));
    Odrv4 I__1420 (
            .O(N__6122),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    InMux I__1419 (
            .O(N__6119),
            .I(N__6115));
    InMux I__1418 (
            .O(N__6118),
            .I(N__6112));
    LocalMux I__1417 (
            .O(N__6115),
            .I(N__6109));
    LocalMux I__1416 (
            .O(N__6112),
            .I(N__6105));
    Span4Mux_v I__1415 (
            .O(N__6109),
            .I(N__6102));
    InMux I__1414 (
            .O(N__6108),
            .I(N__6099));
    Span4Mux_v I__1413 (
            .O(N__6105),
            .I(N__6096));
    Span4Mux_v I__1412 (
            .O(N__6102),
            .I(N__6093));
    LocalMux I__1411 (
            .O(N__6099),
            .I(N__6090));
    Sp12to4 I__1410 (
            .O(N__6096),
            .I(N__6083));
    Sp12to4 I__1409 (
            .O(N__6093),
            .I(N__6083));
    Span12Mux_h I__1408 (
            .O(N__6090),
            .I(N__6083));
    Span12Mux_h I__1407 (
            .O(N__6083),
            .I(N__6080));
    Odrv12 I__1406 (
            .O(N__6080),
            .I(D_UU_AMIGA_in_3));
    IoInMux I__1405 (
            .O(N__6077),
            .I(N__6074));
    LocalMux I__1404 (
            .O(N__6074),
            .I(N__6071));
    Span12Mux_s9_v I__1403 (
            .O(N__6071),
            .I(N__6068));
    Span12Mux_h I__1402 (
            .O(N__6068),
            .I(N__6065));
    Odrv12 I__1401 (
            .O(N__6065),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1400 (
            .O(N__6062),
            .I(N__6059));
    LocalMux I__1399 (
            .O(N__6059),
            .I(N__6056));
    Odrv12 I__1398 (
            .O(N__6056),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    InMux I__1397 (
            .O(N__6053),
            .I(N__6049));
    InMux I__1396 (
            .O(N__6052),
            .I(N__6046));
    LocalMux I__1395 (
            .O(N__6049),
            .I(N__6042));
    LocalMux I__1394 (
            .O(N__6046),
            .I(N__6039));
    InMux I__1393 (
            .O(N__6045),
            .I(N__6036));
    Span4Mux_h I__1392 (
            .O(N__6042),
            .I(N__6033));
    Span4Mux_v I__1391 (
            .O(N__6039),
            .I(N__6028));
    LocalMux I__1390 (
            .O(N__6036),
            .I(N__6028));
    Span4Mux_v I__1389 (
            .O(N__6033),
            .I(N__6025));
    Span4Mux_v I__1388 (
            .O(N__6028),
            .I(N__6022));
    Sp12to4 I__1387 (
            .O(N__6025),
            .I(N__6019));
    Sp12to4 I__1386 (
            .O(N__6022),
            .I(N__6016));
    Span12Mux_v I__1385 (
            .O(N__6019),
            .I(N__6013));
    Span12Mux_h I__1384 (
            .O(N__6016),
            .I(N__6010));
    Odrv12 I__1383 (
            .O(N__6013),
            .I(D_UM_AMIGA_in_3));
    Odrv12 I__1382 (
            .O(N__6010),
            .I(D_UM_AMIGA_in_3));
    IoInMux I__1381 (
            .O(N__6005),
            .I(N__6002));
    LocalMux I__1380 (
            .O(N__6002),
            .I(N__5999));
    Span4Mux_s3_h I__1379 (
            .O(N__5999),
            .I(N__5996));
    Span4Mux_h I__1378 (
            .O(N__5996),
            .I(N__5993));
    Span4Mux_h I__1377 (
            .O(N__5993),
            .I(N__5990));
    Span4Mux_h I__1376 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_v I__1375 (
            .O(N__5987),
            .I(N__5984));
    Odrv4 I__1374 (
            .O(N__5984),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1373 (
            .O(N__5981),
            .I(N__5978));
    LocalMux I__1372 (
            .O(N__5978),
            .I(N__5975));
    Span4Mux_v I__1371 (
            .O(N__5975),
            .I(N__5972));
    Span4Mux_v I__1370 (
            .O(N__5972),
            .I(N__5969));
    Sp12to4 I__1369 (
            .O(N__5969),
            .I(N__5966));
    Span12Mux_h I__1368 (
            .O(N__5966),
            .I(N__5963));
    Odrv12 I__1367 (
            .O(N__5963),
            .I(D_UM_040_in_3));
    IoInMux I__1366 (
            .O(N__5960),
            .I(N__5957));
    LocalMux I__1365 (
            .O(N__5957),
            .I(N__5953));
    InMux I__1364 (
            .O(N__5956),
            .I(N__5950));
    Span4Mux_s3_h I__1363 (
            .O(N__5953),
            .I(N__5947));
    LocalMux I__1362 (
            .O(N__5950),
            .I(N__5944));
    Sp12to4 I__1361 (
            .O(N__5947),
            .I(N__5941));
    Span12Mux_v I__1360 (
            .O(N__5944),
            .I(N__5938));
    Span12Mux_v I__1359 (
            .O(N__5941),
            .I(N__5935));
    Span12Mux_v I__1358 (
            .O(N__5938),
            .I(N__5930));
    Span12Mux_h I__1357 (
            .O(N__5935),
            .I(N__5930));
    Span12Mux_h I__1356 (
            .O(N__5930),
            .I(N__5927));
    Odrv12 I__1355 (
            .O(N__5927),
            .I(D_LL_040_in_3));
    IoInMux I__1354 (
            .O(N__5924),
            .I(N__5921));
    LocalMux I__1353 (
            .O(N__5921),
            .I(N__5918));
    Span4Mux_s3_h I__1352 (
            .O(N__5918),
            .I(N__5915));
    Span4Mux_h I__1351 (
            .O(N__5915),
            .I(N__5912));
    Span4Mux_h I__1350 (
            .O(N__5912),
            .I(N__5909));
    Span4Mux_h I__1349 (
            .O(N__5909),
            .I(N__5906));
    Odrv4 I__1348 (
            .O(N__5906),
            .I(un1_D_UM_040_3));
    InMux I__1347 (
            .O(N__5903),
            .I(N__5899));
    InMux I__1346 (
            .O(N__5902),
            .I(N__5896));
    LocalMux I__1345 (
            .O(N__5899),
            .I(N__5893));
    LocalMux I__1344 (
            .O(N__5896),
            .I(N__5889));
    Span4Mux_h I__1343 (
            .O(N__5893),
            .I(N__5886));
    InMux I__1342 (
            .O(N__5892),
            .I(N__5883));
    Span4Mux_v I__1341 (
            .O(N__5889),
            .I(N__5880));
    Span4Mux_v I__1340 (
            .O(N__5886),
            .I(N__5875));
    LocalMux I__1339 (
            .O(N__5883),
            .I(N__5875));
    Sp12to4 I__1338 (
            .O(N__5880),
            .I(N__5872));
    Span4Mux_v I__1337 (
            .O(N__5875),
            .I(N__5869));
    Span12Mux_h I__1336 (
            .O(N__5872),
            .I(N__5866));
    Sp12to4 I__1335 (
            .O(N__5869),
            .I(N__5863));
    Span12Mux_v I__1334 (
            .O(N__5866),
            .I(N__5858));
    Span12Mux_h I__1333 (
            .O(N__5863),
            .I(N__5858));
    Odrv12 I__1332 (
            .O(N__5858),
            .I(D_UM_AMIGA_in_7));
    InMux I__1331 (
            .O(N__5855),
            .I(N__5852));
    LocalMux I__1330 (
            .O(N__5852),
            .I(N__5849));
    Span4Mux_v I__1329 (
            .O(N__5849),
            .I(N__5846));
    Odrv4 I__1328 (
            .O(N__5846),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1327 (
            .O(N__5843),
            .I(N__5840));
    LocalMux I__1326 (
            .O(N__5840),
            .I(N__5837));
    IoSpan4Mux I__1325 (
            .O(N__5837),
            .I(N__5834));
    Span4Mux_s3_h I__1324 (
            .O(N__5834),
            .I(N__5831));
    Span4Mux_h I__1323 (
            .O(N__5831),
            .I(N__5828));
    Span4Mux_h I__1322 (
            .O(N__5828),
            .I(N__5825));
    Span4Mux_h I__1321 (
            .O(N__5825),
            .I(N__5822));
    Odrv4 I__1320 (
            .O(N__5822),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1319 (
            .O(N__5819),
            .I(N__5816));
    LocalMux I__1318 (
            .O(N__5816),
            .I(N__5813));
    Span4Mux_h I__1317 (
            .O(N__5813),
            .I(N__5810));
    Sp12to4 I__1316 (
            .O(N__5810),
            .I(N__5807));
    Span12Mux_v I__1315 (
            .O(N__5807),
            .I(N__5804));
    Span12Mux_h I__1314 (
            .O(N__5804),
            .I(N__5801));
    Odrv12 I__1313 (
            .O(N__5801),
            .I(D_UM_040_in_4));
    InMux I__1312 (
            .O(N__5798),
            .I(N__5794));
    IoInMux I__1311 (
            .O(N__5797),
            .I(N__5791));
    LocalMux I__1310 (
            .O(N__5794),
            .I(N__5788));
    LocalMux I__1309 (
            .O(N__5791),
            .I(N__5785));
    Span4Mux_v I__1308 (
            .O(N__5788),
            .I(N__5782));
    Span4Mux_s2_h I__1307 (
            .O(N__5785),
            .I(N__5779));
    Sp12to4 I__1306 (
            .O(N__5782),
            .I(N__5776));
    Span4Mux_v I__1305 (
            .O(N__5779),
            .I(N__5773));
    Span12Mux_h I__1304 (
            .O(N__5776),
            .I(N__5770));
    Sp12to4 I__1303 (
            .O(N__5773),
            .I(N__5767));
    Span12Mux_v I__1302 (
            .O(N__5770),
            .I(N__5764));
    Span12Mux_h I__1301 (
            .O(N__5767),
            .I(N__5761));
    Span12Mux_v I__1300 (
            .O(N__5764),
            .I(N__5756));
    Span12Mux_h I__1299 (
            .O(N__5761),
            .I(N__5756));
    Odrv12 I__1298 (
            .O(N__5756),
            .I(D_LL_040_in_4));
    IoInMux I__1297 (
            .O(N__5753),
            .I(N__5750));
    LocalMux I__1296 (
            .O(N__5750),
            .I(N__5747));
    Span4Mux_s3_h I__1295 (
            .O(N__5747),
            .I(N__5744));
    Span4Mux_h I__1294 (
            .O(N__5744),
            .I(N__5741));
    Span4Mux_h I__1293 (
            .O(N__5741),
            .I(N__5738));
    Span4Mux_h I__1292 (
            .O(N__5738),
            .I(N__5735));
    Odrv4 I__1291 (
            .O(N__5735),
            .I(un1_D_UM_040_4));
    InMux I__1290 (
            .O(N__5732),
            .I(N__5729));
    LocalMux I__1289 (
            .O(N__5729),
            .I(N__5726));
    Span4Mux_v I__1288 (
            .O(N__5726),
            .I(N__5723));
    Span4Mux_v I__1287 (
            .O(N__5723),
            .I(N__5720));
    Sp12to4 I__1286 (
            .O(N__5720),
            .I(N__5717));
    Span12Mux_h I__1285 (
            .O(N__5717),
            .I(N__5714));
    Odrv12 I__1284 (
            .O(N__5714),
            .I(D_UM_040_in_7));
    IoInMux I__1283 (
            .O(N__5711),
            .I(N__5708));
    LocalMux I__1282 (
            .O(N__5708),
            .I(N__5705));
    IoSpan4Mux I__1281 (
            .O(N__5705),
            .I(N__5702));
    Span4Mux_s3_h I__1280 (
            .O(N__5702),
            .I(N__5698));
    InMux I__1279 (
            .O(N__5701),
            .I(N__5695));
    Sp12to4 I__1278 (
            .O(N__5698),
            .I(N__5692));
    LocalMux I__1277 (
            .O(N__5695),
            .I(N__5689));
    Span12Mux_v I__1276 (
            .O(N__5692),
            .I(N__5686));
    Span12Mux_v I__1275 (
            .O(N__5689),
            .I(N__5683));
    Span12Mux_h I__1274 (
            .O(N__5686),
            .I(N__5678));
    Span12Mux_v I__1273 (
            .O(N__5683),
            .I(N__5678));
    Span12Mux_h I__1272 (
            .O(N__5678),
            .I(N__5675));
    Odrv12 I__1271 (
            .O(N__5675),
            .I(D_LL_040_in_7));
    IoInMux I__1270 (
            .O(N__5672),
            .I(N__5669));
    LocalMux I__1269 (
            .O(N__5669),
            .I(N__5666));
    Span12Mux_s3_h I__1268 (
            .O(N__5666),
            .I(N__5663));
    Span12Mux_h I__1267 (
            .O(N__5663),
            .I(N__5660));
    Odrv12 I__1266 (
            .O(N__5660),
            .I(un1_D_UM_040_7));
    InMux I__1265 (
            .O(N__5657),
            .I(N__5651));
    InMux I__1264 (
            .O(N__5656),
            .I(N__5648));
    InMux I__1263 (
            .O(N__5655),
            .I(N__5645));
    InMux I__1262 (
            .O(N__5654),
            .I(N__5642));
    LocalMux I__1261 (
            .O(N__5651),
            .I(N__5628));
    LocalMux I__1260 (
            .O(N__5648),
            .I(N__5628));
    LocalMux I__1259 (
            .O(N__5645),
            .I(N__5628));
    LocalMux I__1258 (
            .O(N__5642),
            .I(N__5628));
    InMux I__1257 (
            .O(N__5641),
            .I(N__5625));
    InMux I__1256 (
            .O(N__5640),
            .I(N__5620));
    InMux I__1255 (
            .O(N__5639),
            .I(N__5620));
    InMux I__1254 (
            .O(N__5638),
            .I(N__5615));
    InMux I__1253 (
            .O(N__5637),
            .I(N__5615));
    Span4Mux_v I__1252 (
            .O(N__5628),
            .I(N__5606));
    LocalMux I__1251 (
            .O(N__5625),
            .I(N__5606));
    LocalMux I__1250 (
            .O(N__5620),
            .I(N__5606));
    LocalMux I__1249 (
            .O(N__5615),
            .I(N__5606));
    Span4Mux_v I__1248 (
            .O(N__5606),
            .I(N__5603));
    Span4Mux_h I__1247 (
            .O(N__5603),
            .I(N__5600));
    Sp12to4 I__1246 (
            .O(N__5600),
            .I(N__5597));
    Span12Mux_v I__1245 (
            .O(N__5597),
            .I(N__5594));
    Odrv12 I__1244 (
            .O(N__5594),
            .I(RESETn_c));
    CascadeMux I__1243 (
            .O(N__5591),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ));
    InMux I__1242 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__1241 (
            .O(N__5585),
            .I(N__5582));
    Glb2LocalMux I__1240 (
            .O(N__5582),
            .I(N__5579));
    GlobalMux I__1239 (
            .O(N__5579),
            .I(CLK80));
    IoInMux I__1238 (
            .O(N__5576),
            .I(N__5573));
    LocalMux I__1237 (
            .O(N__5573),
            .I(N__5569));
    IoInMux I__1236 (
            .O(N__5572),
            .I(N__5566));
    Span4Mux_s1_v I__1235 (
            .O(N__5569),
            .I(N__5563));
    LocalMux I__1234 (
            .O(N__5566),
            .I(N__5560));
    Span4Mux_v I__1233 (
            .O(N__5563),
            .I(N__5557));
    IoSpan4Mux I__1232 (
            .O(N__5560),
            .I(N__5554));
    Span4Mux_v I__1231 (
            .O(N__5557),
            .I(N__5551));
    Span4Mux_s3_h I__1230 (
            .O(N__5554),
            .I(N__5548));
    Span4Mux_v I__1229 (
            .O(N__5551),
            .I(N__5545));
    Sp12to4 I__1228 (
            .O(N__5548),
            .I(N__5542));
    Odrv4 I__1227 (
            .O(N__5545),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1226 (
            .O(N__5542),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1225 (
            .O(N__5537),
            .I(N__5534));
    LocalMux I__1224 (
            .O(N__5534),
            .I(N__5531));
    Span12Mux_h I__1223 (
            .O(N__5531),
            .I(N__5528));
    Odrv12 I__1222 (
            .O(N__5528),
            .I(D_LM_AMIGA_in_2));
    InMux I__1221 (
            .O(N__5525),
            .I(N__5521));
    InMux I__1220 (
            .O(N__5524),
            .I(N__5518));
    LocalMux I__1219 (
            .O(N__5521),
            .I(N__5515));
    LocalMux I__1218 (
            .O(N__5518),
            .I(N__5512));
    Span4Mux_v I__1217 (
            .O(N__5515),
            .I(N__5508));
    Span4Mux_v I__1216 (
            .O(N__5512),
            .I(N__5505));
    InMux I__1215 (
            .O(N__5511),
            .I(N__5502));
    Span4Mux_v I__1214 (
            .O(N__5508),
            .I(N__5499));
    Span4Mux_v I__1213 (
            .O(N__5505),
            .I(N__5494));
    LocalMux I__1212 (
            .O(N__5502),
            .I(N__5494));
    Span4Mux_v I__1211 (
            .O(N__5499),
            .I(N__5491));
    Span4Mux_v I__1210 (
            .O(N__5494),
            .I(N__5488));
    Sp12to4 I__1209 (
            .O(N__5491),
            .I(N__5483));
    Sp12to4 I__1208 (
            .O(N__5488),
            .I(N__5483));
    Span12Mux_h I__1207 (
            .O(N__5483),
            .I(N__5480));
    Odrv12 I__1206 (
            .O(N__5480),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1205 (
            .O(N__5477),
            .I(N__5474));
    LocalMux I__1204 (
            .O(N__5474),
            .I(N__5471));
    Span12Mux_s7_h I__1203 (
            .O(N__5471),
            .I(N__5468));
    Span12Mux_v I__1202 (
            .O(N__5468),
            .I(N__5465));
    Odrv12 I__1201 (
            .O(N__5465),
            .I(un1_D_LM_AMIGA_2));
    CascadeMux I__1200 (
            .O(N__5462),
            .I(N__5458));
    InMux I__1199 (
            .O(N__5461),
            .I(N__5453));
    InMux I__1198 (
            .O(N__5458),
            .I(N__5453));
    LocalMux I__1197 (
            .O(N__5453),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    CascadeMux I__1196 (
            .O(N__5450),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ));
    InMux I__1195 (
            .O(N__5447),
            .I(N__5443));
    InMux I__1194 (
            .O(N__5446),
            .I(N__5439));
    LocalMux I__1193 (
            .O(N__5443),
            .I(N__5436));
    InMux I__1192 (
            .O(N__5442),
            .I(N__5433));
    LocalMux I__1191 (
            .O(N__5439),
            .I(N__5429));
    Span4Mux_h I__1190 (
            .O(N__5436),
            .I(N__5423));
    LocalMux I__1189 (
            .O(N__5433),
            .I(N__5423));
    InMux I__1188 (
            .O(N__5432),
            .I(N__5420));
    Span4Mux_v I__1187 (
            .O(N__5429),
            .I(N__5417));
    InMux I__1186 (
            .O(N__5428),
            .I(N__5414));
    Sp12to4 I__1185 (
            .O(N__5423),
            .I(N__5409));
    LocalMux I__1184 (
            .O(N__5420),
            .I(N__5409));
    Span4Mux_v I__1183 (
            .O(N__5417),
            .I(N__5404));
    LocalMux I__1182 (
            .O(N__5414),
            .I(N__5404));
    Span12Mux_v I__1181 (
            .O(N__5409),
            .I(N__5401));
    Span4Mux_v I__1180 (
            .O(N__5404),
            .I(N__5398));
    Odrv12 I__1179 (
            .O(N__5401),
            .I(LBENn_c));
    Odrv4 I__1178 (
            .O(N__5398),
            .I(LBENn_c));
    InMux I__1177 (
            .O(N__5393),
            .I(N__5390));
    LocalMux I__1176 (
            .O(N__5390),
            .I(N__5386));
    CascadeMux I__1175 (
            .O(N__5389),
            .I(N__5383));
    Span4Mux_h I__1174 (
            .O(N__5386),
            .I(N__5380));
    InMux I__1173 (
            .O(N__5383),
            .I(N__5377));
    Odrv4 I__1172 (
            .O(N__5380),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1171 (
            .O(N__5377),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    IoInMux I__1170 (
            .O(N__5372),
            .I(N__5369));
    LocalMux I__1169 (
            .O(N__5369),
            .I(N__5366));
    Span4Mux_s3_v I__1168 (
            .O(N__5366),
            .I(N__5363));
    Span4Mux_v I__1167 (
            .O(N__5363),
            .I(N__5360));
    Span4Mux_v I__1166 (
            .O(N__5360),
            .I(N__5357));
    Span4Mux_v I__1165 (
            .O(N__5357),
            .I(N__5354));
    Odrv4 I__1164 (
            .O(N__5354),
            .I(TAn_1_i));
    InMux I__1163 (
            .O(N__5351),
            .I(N__5342));
    InMux I__1162 (
            .O(N__5350),
            .I(N__5342));
    InMux I__1161 (
            .O(N__5349),
            .I(N__5339));
    InMux I__1160 (
            .O(N__5348),
            .I(N__5334));
    InMux I__1159 (
            .O(N__5347),
            .I(N__5334));
    LocalMux I__1158 (
            .O(N__5342),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1157 (
            .O(N__5339),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1156 (
            .O(N__5334),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    CascadeMux I__1155 (
            .O(N__5327),
            .I(\U111_CYCLE_SM.N_135_cascade_ ));
    InMux I__1154 (
            .O(N__5324),
            .I(N__5321));
    LocalMux I__1153 (
            .O(N__5321),
            .I(\U111_CYCLE_SM.N_128_0 ));
    CascadeMux I__1152 (
            .O(N__5318),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ));
    InMux I__1151 (
            .O(N__5315),
            .I(N__5310));
    InMux I__1150 (
            .O(N__5314),
            .I(N__5307));
    InMux I__1149 (
            .O(N__5313),
            .I(N__5301));
    LocalMux I__1148 (
            .O(N__5310),
            .I(N__5298));
    LocalMux I__1147 (
            .O(N__5307),
            .I(N__5295));
    InMux I__1146 (
            .O(N__5306),
            .I(N__5292));
    InMux I__1145 (
            .O(N__5305),
            .I(N__5287));
    InMux I__1144 (
            .O(N__5304),
            .I(N__5287));
    LocalMux I__1143 (
            .O(N__5301),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    Odrv4 I__1142 (
            .O(N__5298),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    Odrv4 I__1141 (
            .O(N__5295),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1140 (
            .O(N__5292),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1139 (
            .O(N__5287),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    IoInMux I__1138 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__1137 (
            .O(N__5273),
            .I(N__5270));
    Span4Mux_s1_v I__1136 (
            .O(N__5270),
            .I(N__5261));
    InMux I__1135 (
            .O(N__5269),
            .I(N__5256));
    InMux I__1134 (
            .O(N__5268),
            .I(N__5256));
    InMux I__1133 (
            .O(N__5267),
            .I(N__5253));
    InMux I__1132 (
            .O(N__5266),
            .I(N__5250));
    InMux I__1131 (
            .O(N__5265),
            .I(N__5245));
    InMux I__1130 (
            .O(N__5264),
            .I(N__5245));
    Span4Mux_v I__1129 (
            .O(N__5261),
            .I(N__5242));
    LocalMux I__1128 (
            .O(N__5256),
            .I(N__5239));
    LocalMux I__1127 (
            .O(N__5253),
            .I(N__5232));
    LocalMux I__1126 (
            .O(N__5250),
            .I(N__5232));
    LocalMux I__1125 (
            .O(N__5245),
            .I(N__5232));
    Sp12to4 I__1124 (
            .O(N__5242),
            .I(N__5229));
    Span4Mux_v I__1123 (
            .O(N__5239),
            .I(N__5226));
    Span4Mux_v I__1122 (
            .O(N__5232),
            .I(N__5223));
    Span12Mux_h I__1121 (
            .O(N__5229),
            .I(N__5220));
    Sp12to4 I__1120 (
            .O(N__5226),
            .I(N__5215));
    Sp12to4 I__1119 (
            .O(N__5223),
            .I(N__5215));
    Span12Mux_v I__1118 (
            .O(N__5220),
            .I(N__5210));
    Span12Mux_h I__1117 (
            .O(N__5215),
            .I(N__5210));
    Span12Mux_v I__1116 (
            .O(N__5210),
            .I(N__5207));
    Odrv12 I__1115 (
            .O(N__5207),
            .I(TEAn_c));
    InMux I__1114 (
            .O(N__5204),
            .I(N__5201));
    LocalMux I__1113 (
            .O(N__5201),
            .I(N__5198));
    Span4Mux_v I__1112 (
            .O(N__5198),
            .I(N__5195));
    Odrv4 I__1111 (
            .O(N__5195),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    InMux I__1110 (
            .O(N__5192),
            .I(N__5188));
    InMux I__1109 (
            .O(N__5191),
            .I(N__5185));
    LocalMux I__1108 (
            .O(N__5188),
            .I(N__5182));
    LocalMux I__1107 (
            .O(N__5185),
            .I(N__5178));
    Span4Mux_v I__1106 (
            .O(N__5182),
            .I(N__5175));
    InMux I__1105 (
            .O(N__5181),
            .I(N__5172));
    Span4Mux_v I__1104 (
            .O(N__5178),
            .I(N__5169));
    Sp12to4 I__1103 (
            .O(N__5175),
            .I(N__5164));
    LocalMux I__1102 (
            .O(N__5172),
            .I(N__5164));
    Sp12to4 I__1101 (
            .O(N__5169),
            .I(N__5161));
    Span12Mux_h I__1100 (
            .O(N__5164),
            .I(N__5158));
    Span12Mux_h I__1099 (
            .O(N__5161),
            .I(N__5155));
    Odrv12 I__1098 (
            .O(N__5158),
            .I(D_UU_AMIGA_in_7));
    Odrv12 I__1097 (
            .O(N__5155),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1096 (
            .O(N__5150),
            .I(N__5147));
    LocalMux I__1095 (
            .O(N__5147),
            .I(N__5144));
    IoSpan4Mux I__1094 (
            .O(N__5144),
            .I(N__5141));
    Span4Mux_s2_v I__1093 (
            .O(N__5141),
            .I(N__5138));
    Span4Mux_v I__1092 (
            .O(N__5138),
            .I(N__5135));
    Sp12to4 I__1091 (
            .O(N__5135),
            .I(N__5132));
    Odrv12 I__1090 (
            .O(N__5132),
            .I(un1_D_UU_AMIGA_7));
    InMux I__1089 (
            .O(N__5129),
            .I(N__5126));
    LocalMux I__1088 (
            .O(N__5126),
            .I(N__5123));
    Span4Mux_v I__1087 (
            .O(N__5123),
            .I(N__5120));
    Sp12to4 I__1086 (
            .O(N__5120),
            .I(N__5117));
    Span12Mux_h I__1085 (
            .O(N__5117),
            .I(N__5114));
    Odrv12 I__1084 (
            .O(N__5114),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__1083 (
            .O(N__5111),
            .I(N__5108));
    LocalMux I__1082 (
            .O(N__5108),
            .I(N__5105));
    Span4Mux_s3_h I__1081 (
            .O(N__5105),
            .I(N__5102));
    Span4Mux_v I__1080 (
            .O(N__5102),
            .I(N__5099));
    Span4Mux_h I__1079 (
            .O(N__5099),
            .I(N__5096));
    Span4Mux_h I__1078 (
            .O(N__5096),
            .I(N__5093));
    Span4Mux_h I__1077 (
            .O(N__5093),
            .I(N__5090));
    Odrv4 I__1076 (
            .O(N__5090),
            .I(un1_D_LL_AMIGA_2));
    InMux I__1075 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__1074 (
            .O(N__5084),
            .I(N__5081));
    Span12Mux_v I__1073 (
            .O(N__5081),
            .I(N__5078));
    Span12Mux_h I__1072 (
            .O(N__5078),
            .I(N__5075));
    Odrv12 I__1071 (
            .O(N__5075),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__1070 (
            .O(N__5072),
            .I(N__5069));
    LocalMux I__1069 (
            .O(N__5069),
            .I(N__5066));
    Span4Mux_s3_h I__1068 (
            .O(N__5066),
            .I(N__5063));
    Span4Mux_h I__1067 (
            .O(N__5063),
            .I(N__5060));
    Sp12to4 I__1066 (
            .O(N__5060),
            .I(N__5057));
    Span12Mux_s8_v I__1065 (
            .O(N__5057),
            .I(N__5054));
    Odrv12 I__1064 (
            .O(N__5054),
            .I(un1_D_LL_AMIGA_4));
    InMux I__1063 (
            .O(N__5051),
            .I(N__5045));
    InMux I__1062 (
            .O(N__5050),
            .I(N__5045));
    LocalMux I__1061 (
            .O(N__5045),
            .I(N__5042));
    Span4Mux_v I__1060 (
            .O(N__5042),
            .I(N__5039));
    Sp12to4 I__1059 (
            .O(N__5039),
            .I(N__5036));
    Span12Mux_h I__1058 (
            .O(N__5036),
            .I(N__5032));
    InMux I__1057 (
            .O(N__5035),
            .I(N__5029));
    Odrv12 I__1056 (
            .O(N__5032),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__1055 (
            .O(N__5029),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    InMux I__1054 (
            .O(N__5024),
            .I(N__5021));
    LocalMux I__1053 (
            .O(N__5021),
            .I(\U111_CYCLE_SM.N_148 ));
    CascadeMux I__1052 (
            .O(N__5018),
            .I(\U111_CYCLE_SM.N_148_cascade_ ));
    InMux I__1051 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__1050 (
            .O(N__5012),
            .I(\U111_CYCLE_SM.TS_EN_6 ));
    InMux I__1049 (
            .O(N__5009),
            .I(N__5006));
    LocalMux I__1048 (
            .O(N__5006),
            .I(N__5003));
    Odrv4 I__1047 (
            .O(N__5003),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    InMux I__1046 (
            .O(N__5000),
            .I(N__4995));
    InMux I__1045 (
            .O(N__4999),
            .I(N__4992));
    InMux I__1044 (
            .O(N__4998),
            .I(N__4989));
    LocalMux I__1043 (
            .O(N__4995),
            .I(N__4984));
    LocalMux I__1042 (
            .O(N__4992),
            .I(N__4984));
    LocalMux I__1041 (
            .O(N__4989),
            .I(N__4981));
    Span4Mux_v I__1040 (
            .O(N__4984),
            .I(N__4978));
    Span4Mux_v I__1039 (
            .O(N__4981),
            .I(N__4975));
    Sp12to4 I__1038 (
            .O(N__4978),
            .I(N__4970));
    Sp12to4 I__1037 (
            .O(N__4975),
            .I(N__4970));
    Span12Mux_h I__1036 (
            .O(N__4970),
            .I(N__4967));
    Odrv12 I__1035 (
            .O(N__4967),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1034 (
            .O(N__4964),
            .I(N__4961));
    LocalMux I__1033 (
            .O(N__4961),
            .I(N__4958));
    Span4Mux_s3_v I__1032 (
            .O(N__4958),
            .I(N__4955));
    Span4Mux_v I__1031 (
            .O(N__4955),
            .I(N__4952));
    Sp12to4 I__1030 (
            .O(N__4952),
            .I(N__4949));
    Span12Mux_h I__1029 (
            .O(N__4949),
            .I(N__4946));
    Odrv12 I__1028 (
            .O(N__4946),
            .I(un1_D_UU_AMIGA_6));
    InMux I__1027 (
            .O(N__4943),
            .I(N__4940));
    LocalMux I__1026 (
            .O(N__4940),
            .I(N__4937));
    Span4Mux_v I__1025 (
            .O(N__4937),
            .I(N__4932));
    InMux I__1024 (
            .O(N__4936),
            .I(N__4929));
    InMux I__1023 (
            .O(N__4935),
            .I(N__4926));
    Span4Mux_v I__1022 (
            .O(N__4932),
            .I(N__4919));
    LocalMux I__1021 (
            .O(N__4929),
            .I(N__4919));
    LocalMux I__1020 (
            .O(N__4926),
            .I(N__4919));
    Span4Mux_v I__1019 (
            .O(N__4919),
            .I(N__4916));
    Sp12to4 I__1018 (
            .O(N__4916),
            .I(N__4913));
    Span12Mux_h I__1017 (
            .O(N__4913),
            .I(N__4910));
    Odrv12 I__1016 (
            .O(N__4910),
            .I(D_UU_AMIGA_in_0));
    InMux I__1015 (
            .O(N__4907),
            .I(N__4904));
    LocalMux I__1014 (
            .O(N__4904),
            .I(N__4901));
    Odrv4 I__1013 (
            .O(N__4901),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    IoInMux I__1012 (
            .O(N__4898),
            .I(N__4895));
    LocalMux I__1011 (
            .O(N__4895),
            .I(N__4892));
    Span4Mux_s2_v I__1010 (
            .O(N__4892),
            .I(N__4889));
    Span4Mux_v I__1009 (
            .O(N__4889),
            .I(N__4886));
    Span4Mux_v I__1008 (
            .O(N__4886),
            .I(N__4883));
    Sp12to4 I__1007 (
            .O(N__4883),
            .I(N__4880));
    Odrv12 I__1006 (
            .O(N__4880),
            .I(un1_D_UU_AMIGA_0));
    InMux I__1005 (
            .O(N__4877),
            .I(N__4874));
    LocalMux I__1004 (
            .O(N__4874),
            .I(N__4871));
    Odrv12 I__1003 (
            .O(N__4871),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    IoInMux I__1002 (
            .O(N__4868),
            .I(N__4865));
    LocalMux I__1001 (
            .O(N__4865),
            .I(N__4862));
    Span12Mux_s9_v I__1000 (
            .O(N__4862),
            .I(N__4859));
    Span12Mux_h I__999 (
            .O(N__4859),
            .I(N__4856));
    Odrv12 I__998 (
            .O(N__4856),
            .I(un1_D_UU_AMIGA_2));
    InMux I__997 (
            .O(N__4853),
            .I(N__4850));
    LocalMux I__996 (
            .O(N__4850),
            .I(N__4847));
    Odrv12 I__995 (
            .O(N__4847),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    InMux I__994 (
            .O(N__4844),
            .I(N__4841));
    LocalMux I__993 (
            .O(N__4841),
            .I(N__4838));
    Span4Mux_v I__992 (
            .O(N__4838),
            .I(N__4834));
    InMux I__991 (
            .O(N__4837),
            .I(N__4831));
    Span4Mux_v I__990 (
            .O(N__4834),
            .I(N__4828));
    LocalMux I__989 (
            .O(N__4831),
            .I(N__4825));
    Span4Mux_v I__988 (
            .O(N__4828),
            .I(N__4819));
    Span4Mux_v I__987 (
            .O(N__4825),
            .I(N__4819));
    InMux I__986 (
            .O(N__4824),
            .I(N__4816));
    Span4Mux_v I__985 (
            .O(N__4819),
            .I(N__4811));
    LocalMux I__984 (
            .O(N__4816),
            .I(N__4811));
    Span4Mux_v I__983 (
            .O(N__4811),
            .I(N__4808));
    IoSpan4Mux I__982 (
            .O(N__4808),
            .I(N__4805));
    IoSpan4Mux I__981 (
            .O(N__4805),
            .I(N__4802));
    IoSpan4Mux I__980 (
            .O(N__4802),
            .I(N__4799));
    Odrv4 I__979 (
            .O(N__4799),
            .I(D_UM_AMIGA_in_5));
    IoInMux I__978 (
            .O(N__4796),
            .I(N__4793));
    LocalMux I__977 (
            .O(N__4793),
            .I(N__4790));
    Span4Mux_s2_v I__976 (
            .O(N__4790),
            .I(N__4787));
    Span4Mux_v I__975 (
            .O(N__4787),
            .I(N__4784));
    Sp12to4 I__974 (
            .O(N__4784),
            .I(N__4781));
    Span12Mux_h I__973 (
            .O(N__4781),
            .I(N__4778));
    Odrv12 I__972 (
            .O(N__4778),
            .I(un1_D_UM_AMIGA_5));
    InMux I__971 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__970 (
            .O(N__4772),
            .I(\U111_CYCLE_SM.PORT_MISMATCH_2 ));
    CascadeMux I__969 (
            .O(N__4769),
            .I(\U111_CYCLE_SM.N_123_0_cascade_ ));
    InMux I__968 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__967 (
            .O(N__4763),
            .I(\U111_CYCLE_SM.N_121_0 ));
    InMux I__966 (
            .O(N__4760),
            .I(N__4754));
    InMux I__965 (
            .O(N__4759),
            .I(N__4754));
    LocalMux I__964 (
            .O(N__4754),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_0 ));
    IoInMux I__963 (
            .O(N__4751),
            .I(N__4747));
    IoInMux I__962 (
            .O(N__4750),
            .I(N__4744));
    LocalMux I__961 (
            .O(N__4747),
            .I(N__4737));
    LocalMux I__960 (
            .O(N__4744),
            .I(N__4737));
    IoInMux I__959 (
            .O(N__4743),
            .I(N__4734));
    IoInMux I__958 (
            .O(N__4742),
            .I(N__4731));
    IoSpan4Mux I__957 (
            .O(N__4737),
            .I(N__4719));
    LocalMux I__956 (
            .O(N__4734),
            .I(N__4719));
    LocalMux I__955 (
            .O(N__4731),
            .I(N__4719));
    IoInMux I__954 (
            .O(N__4730),
            .I(N__4716));
    IoInMux I__953 (
            .O(N__4729),
            .I(N__4713));
    IoInMux I__952 (
            .O(N__4728),
            .I(N__4710));
    IoInMux I__951 (
            .O(N__4727),
            .I(N__4707));
    IoInMux I__950 (
            .O(N__4726),
            .I(N__4704));
    IoSpan4Mux I__949 (
            .O(N__4719),
            .I(N__4688));
    LocalMux I__948 (
            .O(N__4716),
            .I(N__4688));
    LocalMux I__947 (
            .O(N__4713),
            .I(N__4688));
    LocalMux I__946 (
            .O(N__4710),
            .I(N__4688));
    LocalMux I__945 (
            .O(N__4707),
            .I(N__4688));
    LocalMux I__944 (
            .O(N__4704),
            .I(N__4688));
    IoInMux I__943 (
            .O(N__4703),
            .I(N__4685));
    IoInMux I__942 (
            .O(N__4702),
            .I(N__4682));
    IoInMux I__941 (
            .O(N__4701),
            .I(N__4679));
    IoSpan4Mux I__940 (
            .O(N__4688),
            .I(N__4675));
    LocalMux I__939 (
            .O(N__4685),
            .I(N__4667));
    LocalMux I__938 (
            .O(N__4682),
            .I(N__4667));
    LocalMux I__937 (
            .O(N__4679),
            .I(N__4667));
    IoInMux I__936 (
            .O(N__4678),
            .I(N__4664));
    IoSpan4Mux I__935 (
            .O(N__4675),
            .I(N__4654));
    IoInMux I__934 (
            .O(N__4674),
            .I(N__4651));
    IoSpan4Mux I__933 (
            .O(N__4667),
            .I(N__4643));
    LocalMux I__932 (
            .O(N__4664),
            .I(N__4643));
    IoInMux I__931 (
            .O(N__4663),
            .I(N__4640));
    IoInMux I__930 (
            .O(N__4662),
            .I(N__4633));
    IoInMux I__929 (
            .O(N__4661),
            .I(N__4630));
    IoInMux I__928 (
            .O(N__4660),
            .I(N__4627));
    IoInMux I__927 (
            .O(N__4659),
            .I(N__4624));
    IoInMux I__926 (
            .O(N__4658),
            .I(N__4621));
    IoInMux I__925 (
            .O(N__4657),
            .I(N__4618));
    IoSpan4Mux I__924 (
            .O(N__4654),
            .I(N__4613));
    LocalMux I__923 (
            .O(N__4651),
            .I(N__4613));
    IoInMux I__922 (
            .O(N__4650),
            .I(N__4610));
    IoInMux I__921 (
            .O(N__4649),
            .I(N__4607));
    IoInMux I__920 (
            .O(N__4648),
            .I(N__4604));
    IoSpan4Mux I__919 (
            .O(N__4643),
            .I(N__4599));
    LocalMux I__918 (
            .O(N__4640),
            .I(N__4599));
    IoInMux I__917 (
            .O(N__4639),
            .I(N__4596));
    IoInMux I__916 (
            .O(N__4638),
            .I(N__4593));
    IoInMux I__915 (
            .O(N__4637),
            .I(N__4589));
    IoInMux I__914 (
            .O(N__4636),
            .I(N__4586));
    LocalMux I__913 (
            .O(N__4633),
            .I(N__4575));
    LocalMux I__912 (
            .O(N__4630),
            .I(N__4575));
    LocalMux I__911 (
            .O(N__4627),
            .I(N__4575));
    LocalMux I__910 (
            .O(N__4624),
            .I(N__4575));
    LocalMux I__909 (
            .O(N__4621),
            .I(N__4571));
    LocalMux I__908 (
            .O(N__4618),
            .I(N__4568));
    IoSpan4Mux I__907 (
            .O(N__4613),
            .I(N__4559));
    LocalMux I__906 (
            .O(N__4610),
            .I(N__4559));
    LocalMux I__905 (
            .O(N__4607),
            .I(N__4559));
    LocalMux I__904 (
            .O(N__4604),
            .I(N__4559));
    IoSpan4Mux I__903 (
            .O(N__4599),
            .I(N__4552));
    LocalMux I__902 (
            .O(N__4596),
            .I(N__4552));
    LocalMux I__901 (
            .O(N__4593),
            .I(N__4552));
    IoInMux I__900 (
            .O(N__4592),
            .I(N__4549));
    LocalMux I__899 (
            .O(N__4589),
            .I(N__4544));
    LocalMux I__898 (
            .O(N__4586),
            .I(N__4544));
    IoInMux I__897 (
            .O(N__4585),
            .I(N__4541));
    IoInMux I__896 (
            .O(N__4584),
            .I(N__4538));
    IoSpan4Mux I__895 (
            .O(N__4575),
            .I(N__4535));
    IoInMux I__894 (
            .O(N__4574),
            .I(N__4532));
    Span4Mux_s2_v I__893 (
            .O(N__4571),
            .I(N__4529));
    Span4Mux_s2_v I__892 (
            .O(N__4568),
            .I(N__4526));
    IoSpan4Mux I__891 (
            .O(N__4559),
            .I(N__4521));
    IoSpan4Mux I__890 (
            .O(N__4552),
            .I(N__4521));
    LocalMux I__889 (
            .O(N__4549),
            .I(N__4518));
    Span12Mux_s5_h I__888 (
            .O(N__4544),
            .I(N__4515));
    LocalMux I__887 (
            .O(N__4541),
            .I(N__4510));
    LocalMux I__886 (
            .O(N__4538),
            .I(N__4510));
    Span4Mux_s2_v I__885 (
            .O(N__4535),
            .I(N__4507));
    LocalMux I__884 (
            .O(N__4532),
            .I(N__4504));
    Sp12to4 I__883 (
            .O(N__4529),
            .I(N__4499));
    Sp12to4 I__882 (
            .O(N__4526),
            .I(N__4499));
    Span4Mux_s2_h I__881 (
            .O(N__4521),
            .I(N__4496));
    Span12Mux_s5_h I__880 (
            .O(N__4518),
            .I(N__4493));
    Span12Mux_h I__879 (
            .O(N__4515),
            .I(N__4490));
    Span12Mux_s5_h I__878 (
            .O(N__4510),
            .I(N__4481));
    Sp12to4 I__877 (
            .O(N__4507),
            .I(N__4481));
    Span12Mux_s2_v I__876 (
            .O(N__4504),
            .I(N__4481));
    Span12Mux_h I__875 (
            .O(N__4499),
            .I(N__4481));
    Span4Mux_h I__874 (
            .O(N__4496),
            .I(N__4478));
    Span12Mux_h I__873 (
            .O(N__4493),
            .I(N__4475));
    Span12Mux_v I__872 (
            .O(N__4490),
            .I(N__4468));
    Span12Mux_v I__871 (
            .O(N__4481),
            .I(N__4468));
    Sp12to4 I__870 (
            .O(N__4478),
            .I(N__4468));
    Odrv12 I__869 (
            .O(N__4475),
            .I(D_UU_040_1_i));
    Odrv12 I__868 (
            .O(N__4468),
            .I(D_UU_040_1_i));
    InMux I__867 (
            .O(N__4463),
            .I(N__4458));
    InMux I__866 (
            .O(N__4462),
            .I(N__4452));
    InMux I__865 (
            .O(N__4461),
            .I(N__4452));
    LocalMux I__864 (
            .O(N__4458),
            .I(N__4449));
    InMux I__863 (
            .O(N__4457),
            .I(N__4446));
    LocalMux I__862 (
            .O(N__4452),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__861 (
            .O(N__4449),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__860 (
            .O(N__4446),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    CascadeMux I__859 (
            .O(N__4439),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ));
    InMux I__858 (
            .O(N__4436),
            .I(N__4433));
    LocalMux I__857 (
            .O(N__4433),
            .I(N__4430));
    Span4Mux_v I__856 (
            .O(N__4430),
            .I(N__4427));
    Sp12to4 I__855 (
            .O(N__4427),
            .I(N__4424));
    Span12Mux_h I__854 (
            .O(N__4424),
            .I(N__4421));
    Odrv12 I__853 (
            .O(N__4421),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__852 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__851 (
            .O(N__4415),
            .I(N__4412));
    Span4Mux_s2_h I__850 (
            .O(N__4412),
            .I(N__4409));
    Span4Mux_v I__849 (
            .O(N__4409),
            .I(N__4406));
    Span4Mux_v I__848 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_h I__847 (
            .O(N__4403),
            .I(N__4400));
    Sp12to4 I__846 (
            .O(N__4400),
            .I(N__4397));
    Odrv12 I__845 (
            .O(N__4397),
            .I(un1_D_LM_AMIGA_0));
    IoInMux I__844 (
            .O(N__4394),
            .I(N__4391));
    LocalMux I__843 (
            .O(N__4391),
            .I(N__4388));
    IoSpan4Mux I__842 (
            .O(N__4388),
            .I(N__4385));
    Sp12to4 I__841 (
            .O(N__4385),
            .I(N__4382));
    Span12Mux_s7_v I__840 (
            .O(N__4382),
            .I(N__4379));
    Odrv12 I__839 (
            .O(N__4379),
            .I(TSn_c));
    IoInMux I__838 (
            .O(N__4376),
            .I(N__4369));
    IoInMux I__837 (
            .O(N__4375),
            .I(N__4366));
    IoInMux I__836 (
            .O(N__4374),
            .I(N__4363));
    IoInMux I__835 (
            .O(N__4373),
            .I(N__4360));
    IoInMux I__834 (
            .O(N__4372),
            .I(N__4357));
    LocalMux I__833 (
            .O(N__4369),
            .I(N__4342));
    LocalMux I__832 (
            .O(N__4366),
            .I(N__4342));
    LocalMux I__831 (
            .O(N__4363),
            .I(N__4342));
    LocalMux I__830 (
            .O(N__4360),
            .I(N__4342));
    LocalMux I__829 (
            .O(N__4357),
            .I(N__4342));
    IoInMux I__828 (
            .O(N__4356),
            .I(N__4333));
    IoInMux I__827 (
            .O(N__4355),
            .I(N__4330));
    IoInMux I__826 (
            .O(N__4354),
            .I(N__4327));
    IoInMux I__825 (
            .O(N__4353),
            .I(N__4324));
    IoSpan4Mux I__824 (
            .O(N__4342),
            .I(N__4317));
    IoInMux I__823 (
            .O(N__4341),
            .I(N__4314));
    IoInMux I__822 (
            .O(N__4340),
            .I(N__4311));
    IoInMux I__821 (
            .O(N__4339),
            .I(N__4308));
    IoInMux I__820 (
            .O(N__4338),
            .I(N__4305));
    IoInMux I__819 (
            .O(N__4337),
            .I(N__4299));
    IoInMux I__818 (
            .O(N__4336),
            .I(N__4296));
    LocalMux I__817 (
            .O(N__4333),
            .I(N__4287));
    LocalMux I__816 (
            .O(N__4330),
            .I(N__4287));
    LocalMux I__815 (
            .O(N__4327),
            .I(N__4287));
    LocalMux I__814 (
            .O(N__4324),
            .I(N__4287));
    IoInMux I__813 (
            .O(N__4323),
            .I(N__4283));
    IoInMux I__812 (
            .O(N__4322),
            .I(N__4280));
    IoInMux I__811 (
            .O(N__4321),
            .I(N__4276));
    IoInMux I__810 (
            .O(N__4320),
            .I(N__4273));
    IoSpan4Mux I__809 (
            .O(N__4317),
            .I(N__4262));
    LocalMux I__808 (
            .O(N__4314),
            .I(N__4262));
    LocalMux I__807 (
            .O(N__4311),
            .I(N__4262));
    LocalMux I__806 (
            .O(N__4308),
            .I(N__4262));
    LocalMux I__805 (
            .O(N__4305),
            .I(N__4262));
    IoInMux I__804 (
            .O(N__4304),
            .I(N__4259));
    IoInMux I__803 (
            .O(N__4303),
            .I(N__4250));
    IoInMux I__802 (
            .O(N__4302),
            .I(N__4247));
    LocalMux I__801 (
            .O(N__4299),
            .I(N__4240));
    LocalMux I__800 (
            .O(N__4296),
            .I(N__4240));
    IoSpan4Mux I__799 (
            .O(N__4287),
            .I(N__4237));
    IoInMux I__798 (
            .O(N__4286),
            .I(N__4234));
    LocalMux I__797 (
            .O(N__4283),
            .I(N__4229));
    LocalMux I__796 (
            .O(N__4280),
            .I(N__4229));
    IoInMux I__795 (
            .O(N__4279),
            .I(N__4226));
    LocalMux I__794 (
            .O(N__4276),
            .I(N__4217));
    LocalMux I__793 (
            .O(N__4273),
            .I(N__4217));
    IoSpan4Mux I__792 (
            .O(N__4262),
            .I(N__4217));
    LocalMux I__791 (
            .O(N__4259),
            .I(N__4217));
    IoInMux I__790 (
            .O(N__4258),
            .I(N__4214));
    IoInMux I__789 (
            .O(N__4257),
            .I(N__4211));
    IoInMux I__788 (
            .O(N__4256),
            .I(N__4208));
    IoInMux I__787 (
            .O(N__4255),
            .I(N__4205));
    IoInMux I__786 (
            .O(N__4254),
            .I(N__4202));
    IoInMux I__785 (
            .O(N__4253),
            .I(N__4199));
    LocalMux I__784 (
            .O(N__4250),
            .I(N__4196));
    LocalMux I__783 (
            .O(N__4247),
            .I(N__4193));
    IoInMux I__782 (
            .O(N__4246),
            .I(N__4190));
    IoInMux I__781 (
            .O(N__4245),
            .I(N__4187));
    Span4Mux_s3_h I__780 (
            .O(N__4240),
            .I(N__4182));
    Span4Mux_s2_v I__779 (
            .O(N__4237),
            .I(N__4182));
    LocalMux I__778 (
            .O(N__4234),
            .I(N__4179));
    IoSpan4Mux I__777 (
            .O(N__4229),
            .I(N__4174));
    LocalMux I__776 (
            .O(N__4226),
            .I(N__4174));
    IoSpan4Mux I__775 (
            .O(N__4217),
            .I(N__4171));
    LocalMux I__774 (
            .O(N__4214),
            .I(N__4166));
    LocalMux I__773 (
            .O(N__4211),
            .I(N__4166));
    LocalMux I__772 (
            .O(N__4208),
            .I(N__4163));
    LocalMux I__771 (
            .O(N__4205),
            .I(N__4160));
    LocalMux I__770 (
            .O(N__4202),
            .I(N__4155));
    LocalMux I__769 (
            .O(N__4199),
            .I(N__4155));
    Span4Mux_s3_h I__768 (
            .O(N__4196),
            .I(N__4150));
    Span4Mux_s3_h I__767 (
            .O(N__4193),
            .I(N__4150));
    LocalMux I__766 (
            .O(N__4190),
            .I(N__4145));
    LocalMux I__765 (
            .O(N__4187),
            .I(N__4145));
    Span4Mux_v I__764 (
            .O(N__4182),
            .I(N__4142));
    Span4Mux_s3_h I__763 (
            .O(N__4179),
            .I(N__4135));
    Span4Mux_s3_h I__762 (
            .O(N__4174),
            .I(N__4135));
    Span4Mux_s3_h I__761 (
            .O(N__4171),
            .I(N__4135));
    Span4Mux_s3_h I__760 (
            .O(N__4166),
            .I(N__4130));
    Span4Mux_s3_h I__759 (
            .O(N__4163),
            .I(N__4130));
    Span12Mux_s10_v I__758 (
            .O(N__4160),
            .I(N__4127));
    Span12Mux_s5_v I__757 (
            .O(N__4155),
            .I(N__4114));
    Sp12to4 I__756 (
            .O(N__4150),
            .I(N__4114));
    Span12Mux_s3_h I__755 (
            .O(N__4145),
            .I(N__4114));
    Sp12to4 I__754 (
            .O(N__4142),
            .I(N__4114));
    Sp12to4 I__753 (
            .O(N__4135),
            .I(N__4114));
    Sp12to4 I__752 (
            .O(N__4130),
            .I(N__4114));
    Span12Mux_h I__751 (
            .O(N__4127),
            .I(N__4111));
    Span12Mux_v I__750 (
            .O(N__4114),
            .I(N__4108));
    Odrv12 I__749 (
            .O(N__4111),
            .I(D_UU_AMIGA_1_i));
    Odrv12 I__748 (
            .O(N__4108),
            .I(D_UU_AMIGA_1_i));
    CascadeMux I__747 (
            .O(N__4103),
            .I(N__4100));
    InMux I__746 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__745 (
            .O(N__4097),
            .I(N__4093));
    InMux I__744 (
            .O(N__4096),
            .I(N__4090));
    Odrv4 I__743 (
            .O(N__4093),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__742 (
            .O(N__4090),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    CascadeMux I__741 (
            .O(N__4085),
            .I(N__4082));
    InMux I__740 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__739 (
            .O(N__4079),
            .I(N__4076));
    Odrv12 I__738 (
            .O(N__4076),
            .I(\U111_CYCLE_SM.FLIP_WORD_2 ));
    InMux I__737 (
            .O(N__4073),
            .I(N__4070));
    LocalMux I__736 (
            .O(N__4070),
            .I(N__4067));
    Span4Mux_v I__735 (
            .O(N__4067),
            .I(N__4064));
    Sp12to4 I__734 (
            .O(N__4064),
            .I(N__4061));
    Span12Mux_h I__733 (
            .O(N__4061),
            .I(N__4058));
    Odrv12 I__732 (
            .O(N__4058),
            .I(D_UM_040_in_2));
    IoInMux I__731 (
            .O(N__4055),
            .I(N__4052));
    LocalMux I__730 (
            .O(N__4052),
            .I(N__4048));
    InMux I__729 (
            .O(N__4051),
            .I(N__4045));
    IoSpan4Mux I__728 (
            .O(N__4048),
            .I(N__4042));
    LocalMux I__727 (
            .O(N__4045),
            .I(N__4039));
    Span4Mux_s2_h I__726 (
            .O(N__4042),
            .I(N__4036));
    Span4Mux_v I__725 (
            .O(N__4039),
            .I(N__4033));
    Sp12to4 I__724 (
            .O(N__4036),
            .I(N__4030));
    Sp12to4 I__723 (
            .O(N__4033),
            .I(N__4027));
    Span12Mux_h I__722 (
            .O(N__4030),
            .I(N__4024));
    Span12Mux_h I__721 (
            .O(N__4027),
            .I(N__4021));
    Span12Mux_h I__720 (
            .O(N__4024),
            .I(N__4016));
    Span12Mux_v I__719 (
            .O(N__4021),
            .I(N__4016));
    Odrv12 I__718 (
            .O(N__4016),
            .I(D_LL_040_in_2));
    IoInMux I__717 (
            .O(N__4013),
            .I(N__4010));
    LocalMux I__716 (
            .O(N__4010),
            .I(N__4007));
    IoSpan4Mux I__715 (
            .O(N__4007),
            .I(N__4004));
    Span4Mux_s1_h I__714 (
            .O(N__4004),
            .I(N__4001));
    Sp12to4 I__713 (
            .O(N__4001),
            .I(N__3998));
    Span12Mux_s9_h I__712 (
            .O(N__3998),
            .I(N__3995));
    Odrv12 I__711 (
            .O(N__3995),
            .I(un1_D_UM_040_2));
    IoInMux I__710 (
            .O(N__3992),
            .I(N__3989));
    LocalMux I__709 (
            .O(N__3989),
            .I(N__3985));
    IoInMux I__708 (
            .O(N__3988),
            .I(N__3980));
    Span4Mux_s3_v I__707 (
            .O(N__3985),
            .I(N__3977));
    IoInMux I__706 (
            .O(N__3984),
            .I(N__3974));
    IoInMux I__705 (
            .O(N__3983),
            .I(N__3971));
    LocalMux I__704 (
            .O(N__3980),
            .I(N__3968));
    Span4Mux_h I__703 (
            .O(N__3977),
            .I(N__3965));
    LocalMux I__702 (
            .O(N__3974),
            .I(N__3962));
    LocalMux I__701 (
            .O(N__3971),
            .I(N__3959));
    IoSpan4Mux I__700 (
            .O(N__3968),
            .I(N__3956));
    Span4Mux_h I__699 (
            .O(N__3965),
            .I(N__3951));
    Span4Mux_s3_v I__698 (
            .O(N__3962),
            .I(N__3951));
    Span4Mux_s2_h I__697 (
            .O(N__3959),
            .I(N__3948));
    Span4Mux_s2_h I__696 (
            .O(N__3956),
            .I(N__3945));
    Span4Mux_v I__695 (
            .O(N__3951),
            .I(N__3942));
    Span4Mux_h I__694 (
            .O(N__3948),
            .I(N__3939));
    Sp12to4 I__693 (
            .O(N__3945),
            .I(N__3936));
    Span4Mux_v I__692 (
            .O(N__3942),
            .I(N__3933));
    Span4Mux_h I__691 (
            .O(N__3939),
            .I(N__3930));
    Span12Mux_s11_h I__690 (
            .O(N__3936),
            .I(N__3927));
    Span4Mux_v I__689 (
            .O(N__3933),
            .I(N__3924));
    Span4Mux_h I__688 (
            .O(N__3930),
            .I(N__3921));
    Odrv12 I__687 (
            .O(N__3927),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv4 I__686 (
            .O(N__3924),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv4 I__685 (
            .O(N__3921),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__684 (
            .O(N__3914),
            .I(N__3911));
    LocalMux I__683 (
            .O(N__3911),
            .I(N__3906));
    InMux I__682 (
            .O(N__3910),
            .I(N__3901));
    InMux I__681 (
            .O(N__3909),
            .I(N__3901));
    Span4Mux_v I__680 (
            .O(N__3906),
            .I(N__3896));
    LocalMux I__679 (
            .O(N__3901),
            .I(N__3896));
    Span4Mux_v I__678 (
            .O(N__3896),
            .I(N__3893));
    Span4Mux_v I__677 (
            .O(N__3893),
            .I(N__3890));
    Sp12to4 I__676 (
            .O(N__3890),
            .I(N__3887));
    Span12Mux_h I__675 (
            .O(N__3887),
            .I(N__3884));
    Odrv12 I__674 (
            .O(N__3884),
            .I(D_UU_AMIGA_in_1));
    InMux I__673 (
            .O(N__3881),
            .I(N__3878));
    LocalMux I__672 (
            .O(N__3878),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    InMux I__671 (
            .O(N__3875),
            .I(N__3872));
    LocalMux I__670 (
            .O(N__3872),
            .I(N__3869));
    Span4Mux_v I__669 (
            .O(N__3869),
            .I(N__3866));
    Sp12to4 I__668 (
            .O(N__3866),
            .I(N__3863));
    Span12Mux_h I__667 (
            .O(N__3863),
            .I(N__3860));
    Odrv12 I__666 (
            .O(N__3860),
            .I(D_UU_040_in_2));
    IoInMux I__665 (
            .O(N__3857),
            .I(N__3853));
    InMux I__664 (
            .O(N__3856),
            .I(N__3850));
    LocalMux I__663 (
            .O(N__3853),
            .I(N__3847));
    LocalMux I__662 (
            .O(N__3850),
            .I(N__3844));
    Span12Mux_s9_h I__661 (
            .O(N__3847),
            .I(N__3841));
    Span12Mux_v I__660 (
            .O(N__3844),
            .I(N__3838));
    Span12Mux_v I__659 (
            .O(N__3841),
            .I(N__3835));
    Span12Mux_v I__658 (
            .O(N__3838),
            .I(N__3832));
    Span12Mux_h I__657 (
            .O(N__3835),
            .I(N__3829));
    Span12Mux_h I__656 (
            .O(N__3832),
            .I(N__3826));
    Odrv12 I__655 (
            .O(N__3829),
            .I(D_LM_040_in_2));
    Odrv12 I__654 (
            .O(N__3826),
            .I(D_LM_040_in_2));
    IoInMux I__653 (
            .O(N__3821),
            .I(N__3818));
    LocalMux I__652 (
            .O(N__3818),
            .I(N__3815));
    IoSpan4Mux I__651 (
            .O(N__3815),
            .I(N__3812));
    Sp12to4 I__650 (
            .O(N__3812),
            .I(N__3809));
    Span12Mux_s6_v I__649 (
            .O(N__3809),
            .I(N__3806));
    Odrv12 I__648 (
            .O(N__3806),
            .I(un1_D_UU_040_2));
    IoInMux I__647 (
            .O(N__3803),
            .I(N__3799));
    InMux I__646 (
            .O(N__3802),
            .I(N__3796));
    LocalMux I__645 (
            .O(N__3799),
            .I(N__3793));
    LocalMux I__644 (
            .O(N__3796),
            .I(N__3790));
    IoSpan4Mux I__643 (
            .O(N__3793),
            .I(N__3787));
    Span4Mux_h I__642 (
            .O(N__3790),
            .I(N__3784));
    Span4Mux_s3_h I__641 (
            .O(N__3787),
            .I(N__3781));
    Sp12to4 I__640 (
            .O(N__3784),
            .I(N__3778));
    Sp12to4 I__639 (
            .O(N__3781),
            .I(N__3775));
    Span12Mux_v I__638 (
            .O(N__3778),
            .I(N__3772));
    Span12Mux_v I__637 (
            .O(N__3775),
            .I(N__3769));
    Span12Mux_v I__636 (
            .O(N__3772),
            .I(N__3764));
    Span12Mux_h I__635 (
            .O(N__3769),
            .I(N__3764));
    Span12Mux_h I__634 (
            .O(N__3764),
            .I(N__3761));
    Odrv12 I__633 (
            .O(N__3761),
            .I(D_LL_040_in_5));
    InMux I__632 (
            .O(N__3758),
            .I(N__3755));
    LocalMux I__631 (
            .O(N__3755),
            .I(N__3752));
    Span4Mux_v I__630 (
            .O(N__3752),
            .I(N__3749));
    Span4Mux_h I__629 (
            .O(N__3749),
            .I(N__3746));
    Sp12to4 I__628 (
            .O(N__3746),
            .I(N__3743));
    Span12Mux_h I__627 (
            .O(N__3743),
            .I(N__3740));
    Odrv12 I__626 (
            .O(N__3740),
            .I(D_UM_040_in_5));
    IoInMux I__625 (
            .O(N__3737),
            .I(N__3734));
    LocalMux I__624 (
            .O(N__3734),
            .I(N__3731));
    Span4Mux_s0_v I__623 (
            .O(N__3731),
            .I(N__3728));
    Sp12to4 I__622 (
            .O(N__3728),
            .I(N__3725));
    Span12Mux_h I__621 (
            .O(N__3725),
            .I(N__3722));
    Odrv12 I__620 (
            .O(N__3722),
            .I(un1_D_UM_040_5));
    IoInMux I__619 (
            .O(N__3719),
            .I(N__3716));
    LocalMux I__618 (
            .O(N__3716),
            .I(N__3713));
    Odrv12 I__617 (
            .O(N__3713),
            .I(LBENn_c_i_0));
    InMux I__616 (
            .O(N__3710),
            .I(N__3707));
    LocalMux I__615 (
            .O(N__3707),
            .I(N__3704));
    Span4Mux_v I__614 (
            .O(N__3704),
            .I(N__3701));
    Sp12to4 I__613 (
            .O(N__3701),
            .I(N__3698));
    Span12Mux_h I__612 (
            .O(N__3698),
            .I(N__3695));
    Odrv12 I__611 (
            .O(N__3695),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__610 (
            .O(N__3692),
            .I(N__3689));
    LocalMux I__609 (
            .O(N__3689),
            .I(N__3686));
    IoSpan4Mux I__608 (
            .O(N__3686),
            .I(N__3683));
    Span4Mux_s3_h I__607 (
            .O(N__3683),
            .I(N__3680));
    Sp12to4 I__606 (
            .O(N__3680),
            .I(N__3677));
    Span12Mux_h I__605 (
            .O(N__3677),
            .I(N__3674));
    Odrv12 I__604 (
            .O(N__3674),
            .I(un1_D_LL_AMIGA_6));
    InMux I__603 (
            .O(N__3671),
            .I(N__3668));
    LocalMux I__602 (
            .O(N__3668),
            .I(N__3665));
    Span4Mux_v I__601 (
            .O(N__3665),
            .I(N__3662));
    Sp12to4 I__600 (
            .O(N__3662),
            .I(N__3659));
    Span12Mux_h I__599 (
            .O(N__3659),
            .I(N__3656));
    Odrv12 I__598 (
            .O(N__3656),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__597 (
            .O(N__3653),
            .I(N__3650));
    LocalMux I__596 (
            .O(N__3650),
            .I(N__3647));
    IoSpan4Mux I__595 (
            .O(N__3647),
            .I(N__3644));
    Span4Mux_s3_h I__594 (
            .O(N__3644),
            .I(N__3641));
    Sp12to4 I__593 (
            .O(N__3641),
            .I(N__3638));
    Span12Mux_h I__592 (
            .O(N__3638),
            .I(N__3635));
    Odrv12 I__591 (
            .O(N__3635),
            .I(un1_D_LL_AMIGA_5));
    InMux I__590 (
            .O(N__3632),
            .I(N__3629));
    LocalMux I__589 (
            .O(N__3629),
            .I(N__3626));
    Sp12to4 I__588 (
            .O(N__3626),
            .I(N__3622));
    InMux I__587 (
            .O(N__3625),
            .I(N__3619));
    Span12Mux_v I__586 (
            .O(N__3622),
            .I(N__3614));
    LocalMux I__585 (
            .O(N__3619),
            .I(N__3614));
    Span12Mux_h I__584 (
            .O(N__3614),
            .I(N__3611));
    Odrv12 I__583 (
            .O(N__3611),
            .I(A_040_c_1));
    InMux I__582 (
            .O(N__3608),
            .I(N__3605));
    LocalMux I__581 (
            .O(N__3605),
            .I(N__3602));
    Span4Mux_v I__580 (
            .O(N__3602),
            .I(N__3599));
    Sp12to4 I__579 (
            .O(N__3599),
            .I(N__3596));
    Span12Mux_h I__578 (
            .O(N__3596),
            .I(N__3593));
    Odrv12 I__577 (
            .O(N__3593),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__576 (
            .O(N__3590),
            .I(N__3587));
    LocalMux I__575 (
            .O(N__3587),
            .I(N__3584));
    IoSpan4Mux I__574 (
            .O(N__3584),
            .I(N__3581));
    Span4Mux_s3_h I__573 (
            .O(N__3581),
            .I(N__3578));
    Sp12to4 I__572 (
            .O(N__3578),
            .I(N__3575));
    Span12Mux_h I__571 (
            .O(N__3575),
            .I(N__3572));
    Odrv12 I__570 (
            .O(N__3572),
            .I(un1_D_LL_AMIGA_7));
    InMux I__569 (
            .O(N__3569),
            .I(N__3566));
    LocalMux I__568 (
            .O(N__3566),
            .I(N__3563));
    Span4Mux_v I__567 (
            .O(N__3563),
            .I(N__3560));
    Sp12to4 I__566 (
            .O(N__3560),
            .I(N__3557));
    Span12Mux_h I__565 (
            .O(N__3557),
            .I(N__3554));
    Odrv12 I__564 (
            .O(N__3554),
            .I(D_UU_040_in_4));
    IoInMux I__563 (
            .O(N__3551),
            .I(N__3548));
    LocalMux I__562 (
            .O(N__3548),
            .I(N__3545));
    Span4Mux_s1_h I__561 (
            .O(N__3545),
            .I(N__3542));
    Sp12to4 I__560 (
            .O(N__3542),
            .I(N__3538));
    InMux I__559 (
            .O(N__3541),
            .I(N__3535));
    Span12Mux_v I__558 (
            .O(N__3538),
            .I(N__3532));
    LocalMux I__557 (
            .O(N__3535),
            .I(N__3529));
    Span12Mux_h I__556 (
            .O(N__3532),
            .I(N__3526));
    Span12Mux_h I__555 (
            .O(N__3529),
            .I(N__3523));
    Span12Mux_h I__554 (
            .O(N__3526),
            .I(N__3520));
    Span12Mux_v I__553 (
            .O(N__3523),
            .I(N__3517));
    Odrv12 I__552 (
            .O(N__3520),
            .I(D_LM_040_in_4));
    Odrv12 I__551 (
            .O(N__3517),
            .I(D_LM_040_in_4));
    IoInMux I__550 (
            .O(N__3512),
            .I(N__3509));
    LocalMux I__549 (
            .O(N__3509),
            .I(N__3506));
    Span4Mux_s2_v I__548 (
            .O(N__3506),
            .I(N__3503));
    Span4Mux_h I__547 (
            .O(N__3503),
            .I(N__3500));
    Span4Mux_v I__546 (
            .O(N__3500),
            .I(N__3497));
    Odrv4 I__545 (
            .O(N__3497),
            .I(un1_D_UU_040_4));
    InMux I__544 (
            .O(N__3494),
            .I(N__3491));
    LocalMux I__543 (
            .O(N__3491),
            .I(N__3488));
    Span4Mux_v I__542 (
            .O(N__3488),
            .I(N__3485));
    Span4Mux_h I__541 (
            .O(N__3485),
            .I(N__3482));
    Sp12to4 I__540 (
            .O(N__3482),
            .I(N__3479));
    Span12Mux_h I__539 (
            .O(N__3479),
            .I(N__3476));
    Odrv12 I__538 (
            .O(N__3476),
            .I(D_UU_040_in_0));
    IoInMux I__537 (
            .O(N__3473),
            .I(N__3470));
    LocalMux I__536 (
            .O(N__3470),
            .I(N__3466));
    InMux I__535 (
            .O(N__3469),
            .I(N__3463));
    IoSpan4Mux I__534 (
            .O(N__3466),
            .I(N__3460));
    LocalMux I__533 (
            .O(N__3463),
            .I(N__3457));
    IoSpan4Mux I__532 (
            .O(N__3460),
            .I(N__3454));
    Sp12to4 I__531 (
            .O(N__3457),
            .I(N__3451));
    Span4Mux_s2_h I__530 (
            .O(N__3454),
            .I(N__3448));
    Span12Mux_v I__529 (
            .O(N__3451),
            .I(N__3445));
    Sp12to4 I__528 (
            .O(N__3448),
            .I(N__3442));
    Span12Mux_v I__527 (
            .O(N__3445),
            .I(N__3437));
    Span12Mux_h I__526 (
            .O(N__3442),
            .I(N__3437));
    Span12Mux_h I__525 (
            .O(N__3437),
            .I(N__3434));
    Odrv12 I__524 (
            .O(N__3434),
            .I(D_LM_040_in_0));
    IoInMux I__523 (
            .O(N__3431),
            .I(N__3428));
    LocalMux I__522 (
            .O(N__3428),
            .I(N__3425));
    IoSpan4Mux I__521 (
            .O(N__3425),
            .I(N__3422));
    Span4Mux_s2_v I__520 (
            .O(N__3422),
            .I(N__3419));
    Span4Mux_v I__519 (
            .O(N__3419),
            .I(N__3416));
    Odrv4 I__518 (
            .O(N__3416),
            .I(un1_D_UU_040_0));
    IoInMux I__517 (
            .O(N__3413),
            .I(N__3410));
    LocalMux I__516 (
            .O(N__3410),
            .I(N__3407));
    IoSpan4Mux I__515 (
            .O(N__3407),
            .I(N__3404));
    Sp12to4 I__514 (
            .O(N__3404),
            .I(N__3401));
    Span12Mux_s7_h I__513 (
            .O(N__3401),
            .I(N__3398));
    Odrv12 I__512 (
            .O(N__3398),
            .I(un1_D_UM_AMIGA_0));
    InMux I__511 (
            .O(N__3395),
            .I(N__3392));
    LocalMux I__510 (
            .O(N__3392),
            .I(N__3389));
    Span12Mux_h I__509 (
            .O(N__3389),
            .I(N__3386));
    Odrv12 I__508 (
            .O(N__3386),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__507 (
            .O(N__3383),
            .I(N__3380));
    LocalMux I__506 (
            .O(N__3380),
            .I(N__3377));
    Span4Mux_s0_h I__505 (
            .O(N__3377),
            .I(N__3374));
    Span4Mux_h I__504 (
            .O(N__3374),
            .I(N__3371));
    Span4Mux_h I__503 (
            .O(N__3371),
            .I(N__3368));
    Sp12to4 I__502 (
            .O(N__3368),
            .I(N__3365));
    Span12Mux_v I__501 (
            .O(N__3365),
            .I(N__3362));
    Odrv12 I__500 (
            .O(N__3362),
            .I(un1_D_LM_AMIGA_1));
    InMux I__499 (
            .O(N__3359),
            .I(N__3356));
    LocalMux I__498 (
            .O(N__3356),
            .I(N__3353));
    Span4Mux_v I__497 (
            .O(N__3353),
            .I(N__3349));
    InMux I__496 (
            .O(N__3352),
            .I(N__3346));
    Span4Mux_v I__495 (
            .O(N__3349),
            .I(N__3343));
    LocalMux I__494 (
            .O(N__3346),
            .I(N__3340));
    Span4Mux_v I__493 (
            .O(N__3343),
            .I(N__3336));
    Span4Mux_v I__492 (
            .O(N__3340),
            .I(N__3333));
    InMux I__491 (
            .O(N__3339),
            .I(N__3330));
    Sp12to4 I__490 (
            .O(N__3336),
            .I(N__3323));
    Sp12to4 I__489 (
            .O(N__3333),
            .I(N__3323));
    LocalMux I__488 (
            .O(N__3330),
            .I(N__3323));
    Span12Mux_h I__487 (
            .O(N__3323),
            .I(N__3320));
    Odrv12 I__486 (
            .O(N__3320),
            .I(D_UM_AMIGA_in_0));
    InMux I__485 (
            .O(N__3317),
            .I(N__3314));
    LocalMux I__484 (
            .O(N__3314),
            .I(N__3311));
    Odrv4 I__483 (
            .O(N__3311),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    IoInMux I__482 (
            .O(N__3308),
            .I(N__3305));
    LocalMux I__481 (
            .O(N__3305),
            .I(N__3302));
    Span4Mux_s2_h I__480 (
            .O(N__3302),
            .I(N__3299));
    Span4Mux_h I__479 (
            .O(N__3299),
            .I(N__3296));
    Sp12to4 I__478 (
            .O(N__3296),
            .I(N__3293));
    Span12Mux_v I__477 (
            .O(N__3293),
            .I(N__3290));
    Span12Mux_h I__476 (
            .O(N__3290),
            .I(N__3287));
    Odrv12 I__475 (
            .O(N__3287),
            .I(un1_D_UM_AMIGA_1));
    InMux I__474 (
            .O(N__3284),
            .I(N__3281));
    LocalMux I__473 (
            .O(N__3281),
            .I(N__3278));
    Span4Mux_v I__472 (
            .O(N__3278),
            .I(N__3273));
    InMux I__471 (
            .O(N__3277),
            .I(N__3268));
    InMux I__470 (
            .O(N__3276),
            .I(N__3268));
    Sp12to4 I__469 (
            .O(N__3273),
            .I(N__3265));
    LocalMux I__468 (
            .O(N__3268),
            .I(N__3262));
    Span12Mux_h I__467 (
            .O(N__3265),
            .I(N__3259));
    Span12Mux_v I__466 (
            .O(N__3262),
            .I(N__3256));
    Span12Mux_v I__465 (
            .O(N__3259),
            .I(N__3253));
    Span12Mux_h I__464 (
            .O(N__3256),
            .I(N__3250));
    Odrv12 I__463 (
            .O(N__3253),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__462 (
            .O(N__3250),
            .I(D_UM_AMIGA_in_1));
    InMux I__461 (
            .O(N__3245),
            .I(N__3242));
    LocalMux I__460 (
            .O(N__3242),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__459 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__458 (
            .O(N__3236),
            .I(N__3233));
    IoSpan4Mux I__457 (
            .O(N__3233),
            .I(N__3230));
    Span4Mux_s3_h I__456 (
            .O(N__3230),
            .I(N__3227));
    Sp12to4 I__455 (
            .O(N__3227),
            .I(N__3224));
    Span12Mux_s8_h I__454 (
            .O(N__3224),
            .I(N__3221));
    Span12Mux_v I__453 (
            .O(N__3221),
            .I(N__3218));
    Odrv12 I__452 (
            .O(N__3218),
            .I(un1_D_UU_AMIGA_1));
    InMux I__451 (
            .O(N__3215),
            .I(N__3212));
    LocalMux I__450 (
            .O(N__3212),
            .I(N__3209));
    Span12Mux_v I__449 (
            .O(N__3209),
            .I(N__3206));
    Odrv12 I__448 (
            .O(N__3206),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__447 (
            .O(N__3203),
            .I(N__3200));
    LocalMux I__446 (
            .O(N__3200),
            .I(N__3197));
    IoSpan4Mux I__445 (
            .O(N__3197),
            .I(N__3194));
    Span4Mux_s3_h I__444 (
            .O(N__3194),
            .I(N__3191));
    Sp12to4 I__443 (
            .O(N__3191),
            .I(N__3188));
    Span12Mux_s8_h I__442 (
            .O(N__3188),
            .I(N__3185));
    Span12Mux_h I__441 (
            .O(N__3185),
            .I(N__3182));
    Odrv12 I__440 (
            .O(N__3182),
            .I(un1_D_LM_AMIGA_5));
    InMux I__439 (
            .O(N__3179),
            .I(N__3176));
    LocalMux I__438 (
            .O(N__3176),
            .I(N__3173));
    Span12Mux_v I__437 (
            .O(N__3173),
            .I(N__3170));
    Odrv12 I__436 (
            .O(N__3170),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__435 (
            .O(N__3167),
            .I(N__3164));
    LocalMux I__434 (
            .O(N__3164),
            .I(N__3161));
    Span12Mux_s8_h I__433 (
            .O(N__3161),
            .I(N__3158));
    Span12Mux_h I__432 (
            .O(N__3158),
            .I(N__3155));
    Odrv12 I__431 (
            .O(N__3155),
            .I(un1_D_LM_AMIGA_7));
    InMux I__430 (
            .O(N__3152),
            .I(N__3149));
    LocalMux I__429 (
            .O(N__3149),
            .I(N__3146));
    Span4Mux_h I__428 (
            .O(N__3146),
            .I(N__3143));
    Span4Mux_v I__427 (
            .O(N__3143),
            .I(N__3140));
    Sp12to4 I__426 (
            .O(N__3140),
            .I(N__3137));
    Odrv12 I__425 (
            .O(N__3137),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__424 (
            .O(N__3134),
            .I(N__3131));
    LocalMux I__423 (
            .O(N__3131),
            .I(N__3128));
    Span12Mux_s9_h I__422 (
            .O(N__3128),
            .I(N__3125));
    Odrv12 I__421 (
            .O(N__3125),
            .I(un1_D_LM_AMIGA_6));
    IoInMux I__420 (
            .O(N__3122),
            .I(N__3118));
    IoInMux I__419 (
            .O(N__3121),
            .I(N__3115));
    LocalMux I__418 (
            .O(N__3118),
            .I(N__3112));
    LocalMux I__417 (
            .O(N__3115),
            .I(N__3109));
    Span4Mux_s2_v I__416 (
            .O(N__3112),
            .I(N__3106));
    Span4Mux_s2_v I__415 (
            .O(N__3109),
            .I(N__3103));
    Span4Mux_h I__414 (
            .O(N__3106),
            .I(N__3100));
    Span4Mux_h I__413 (
            .O(N__3103),
            .I(N__3097));
    Span4Mux_v I__412 (
            .O(N__3100),
            .I(N__3092));
    Span4Mux_v I__411 (
            .O(N__3097),
            .I(N__3092));
    Odrv4 I__410 (
            .O(N__3092),
            .I(CONSTANT_ONE_NET));
    IoInMux I__409 (
            .O(N__3089),
            .I(N__3086));
    LocalMux I__408 (
            .O(N__3086),
            .I(N__3083));
    IoSpan4Mux I__407 (
            .O(N__3083),
            .I(N__3079));
    InMux I__406 (
            .O(N__3082),
            .I(N__3076));
    Span4Mux_s2_h I__405 (
            .O(N__3079),
            .I(N__3073));
    LocalMux I__404 (
            .O(N__3076),
            .I(N__3070));
    Sp12to4 I__403 (
            .O(N__3073),
            .I(N__3067));
    Span4Mux_v I__402 (
            .O(N__3070),
            .I(N__3064));
    Span12Mux_h I__401 (
            .O(N__3067),
            .I(N__3059));
    Sp12to4 I__400 (
            .O(N__3064),
            .I(N__3059));
    Span12Mux_h I__399 (
            .O(N__3059),
            .I(N__3056));
    Odrv12 I__398 (
            .O(N__3056),
            .I(D_LM_040_in_7));
    InMux I__397 (
            .O(N__3053),
            .I(N__3050));
    LocalMux I__396 (
            .O(N__3050),
            .I(N__3047));
    Span4Mux_v I__395 (
            .O(N__3047),
            .I(N__3044));
    Span4Mux_h I__394 (
            .O(N__3044),
            .I(N__3041));
    Sp12to4 I__393 (
            .O(N__3041),
            .I(N__3038));
    Span12Mux_h I__392 (
            .O(N__3038),
            .I(N__3035));
    Odrv12 I__391 (
            .O(N__3035),
            .I(D_UU_040_in_7));
    IoInMux I__390 (
            .O(N__3032),
            .I(N__3029));
    LocalMux I__389 (
            .O(N__3029),
            .I(N__3026));
    Span4Mux_s3_v I__388 (
            .O(N__3026),
            .I(N__3023));
    Sp12to4 I__387 (
            .O(N__3023),
            .I(N__3020));
    Span12Mux_s11_h I__386 (
            .O(N__3020),
            .I(N__3017));
    Odrv12 I__385 (
            .O(N__3017),
            .I(un1_D_UU_040_7));
    InMux I__384 (
            .O(N__3014),
            .I(N__3011));
    LocalMux I__383 (
            .O(N__3011),
            .I(N__3008));
    Span12Mux_h I__382 (
            .O(N__3008),
            .I(N__3005));
    Odrv12 I__381 (
            .O(N__3005),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__380 (
            .O(N__3002),
            .I(N__2999));
    LocalMux I__379 (
            .O(N__2999),
            .I(N__2996));
    Span4Mux_s0_h I__378 (
            .O(N__2996),
            .I(N__2993));
    Sp12to4 I__377 (
            .O(N__2993),
            .I(N__2990));
    Span12Mux_v I__376 (
            .O(N__2990),
            .I(N__2987));
    Span12Mux_h I__375 (
            .O(N__2987),
            .I(N__2984));
    Odrv12 I__374 (
            .O(N__2984),
            .I(un1_D_LM_AMIGA_3));
    InMux I__373 (
            .O(N__2981),
            .I(N__2978));
    LocalMux I__372 (
            .O(N__2978),
            .I(N__2975));
    Span4Mux_v I__371 (
            .O(N__2975),
            .I(N__2972));
    Sp12to4 I__370 (
            .O(N__2972),
            .I(N__2969));
    Span12Mux_h I__369 (
            .O(N__2969),
            .I(N__2966));
    Odrv12 I__368 (
            .O(N__2966),
            .I(D_UM_040_in_0));
    IoInMux I__367 (
            .O(N__2963),
            .I(N__2959));
    InMux I__366 (
            .O(N__2962),
            .I(N__2956));
    LocalMux I__365 (
            .O(N__2959),
            .I(N__2953));
    LocalMux I__364 (
            .O(N__2956),
            .I(N__2950));
    IoSpan4Mux I__363 (
            .O(N__2953),
            .I(N__2947));
    Span4Mux_v I__362 (
            .O(N__2950),
            .I(N__2944));
    Span4Mux_s2_h I__361 (
            .O(N__2947),
            .I(N__2941));
    Sp12to4 I__360 (
            .O(N__2944),
            .I(N__2938));
    Sp12to4 I__359 (
            .O(N__2941),
            .I(N__2935));
    Span12Mux_v I__358 (
            .O(N__2938),
            .I(N__2930));
    Span12Mux_h I__357 (
            .O(N__2935),
            .I(N__2930));
    Span12Mux_h I__356 (
            .O(N__2930),
            .I(N__2927));
    Odrv12 I__355 (
            .O(N__2927),
            .I(D_LL_040_in_0));
    IoInMux I__354 (
            .O(N__2924),
            .I(N__2921));
    LocalMux I__353 (
            .O(N__2921),
            .I(N__2918));
    Span4Mux_s3_h I__352 (
            .O(N__2918),
            .I(N__2915));
    Sp12to4 I__351 (
            .O(N__2915),
            .I(N__2912));
    Span12Mux_v I__350 (
            .O(N__2912),
            .I(N__2909));
    Odrv12 I__349 (
            .O(N__2909),
            .I(un1_D_UM_040_0));
    InMux I__348 (
            .O(N__2906),
            .I(N__2903));
    LocalMux I__347 (
            .O(N__2903),
            .I(N__2900));
    Span4Mux_v I__346 (
            .O(N__2900),
            .I(N__2897));
    Span4Mux_v I__345 (
            .O(N__2897),
            .I(N__2894));
    Sp12to4 I__344 (
            .O(N__2894),
            .I(N__2891));
    Span12Mux_h I__343 (
            .O(N__2891),
            .I(N__2888));
    Odrv12 I__342 (
            .O(N__2888),
            .I(D_UU_040_in_1));
    IoInMux I__341 (
            .O(N__2885),
            .I(N__2882));
    LocalMux I__340 (
            .O(N__2882),
            .I(N__2878));
    InMux I__339 (
            .O(N__2881),
            .I(N__2875));
    Span4Mux_s3_h I__338 (
            .O(N__2878),
            .I(N__2872));
    LocalMux I__337 (
            .O(N__2875),
            .I(N__2869));
    Span4Mux_h I__336 (
            .O(N__2872),
            .I(N__2866));
    Span4Mux_h I__335 (
            .O(N__2869),
            .I(N__2863));
    Span4Mux_h I__334 (
            .O(N__2866),
            .I(N__2860));
    Sp12to4 I__333 (
            .O(N__2863),
            .I(N__2857));
    Sp12to4 I__332 (
            .O(N__2860),
            .I(N__2852));
    Span12Mux_v I__331 (
            .O(N__2857),
            .I(N__2852));
    Span12Mux_v I__330 (
            .O(N__2852),
            .I(N__2849));
    Span12Mux_h I__329 (
            .O(N__2849),
            .I(N__2846));
    Odrv12 I__328 (
            .O(N__2846),
            .I(D_LM_040_in_1));
    IoInMux I__327 (
            .O(N__2843),
            .I(N__2840));
    LocalMux I__326 (
            .O(N__2840),
            .I(N__2837));
    Span4Mux_s3_h I__325 (
            .O(N__2837),
            .I(N__2834));
    Sp12to4 I__324 (
            .O(N__2834),
            .I(N__2831));
    Span12Mux_s8_v I__323 (
            .O(N__2831),
            .I(N__2828));
    Odrv12 I__322 (
            .O(N__2828),
            .I(un1_D_UU_040_1));
    InMux I__321 (
            .O(N__2825),
            .I(N__2822));
    LocalMux I__320 (
            .O(N__2822),
            .I(N__2819));
    Span4Mux_h I__319 (
            .O(N__2819),
            .I(N__2816));
    Span4Mux_v I__318 (
            .O(N__2816),
            .I(N__2813));
    Odrv4 I__317 (
            .O(N__2813),
            .I(A_040_c_0));
    IoInMux I__316 (
            .O(N__2810),
            .I(N__2807));
    LocalMux I__315 (
            .O(N__2807),
            .I(N__2804));
    Span4Mux_s2_v I__314 (
            .O(N__2804),
            .I(N__2801));
    Span4Mux_v I__313 (
            .O(N__2801),
            .I(N__2798));
    Odrv4 I__312 (
            .O(N__2798),
            .I(A_AMIGA_c_0));
    IoInMux I__311 (
            .O(N__2795),
            .I(N__2792));
    LocalMux I__310 (
            .O(N__2792),
            .I(N__2789));
    Span4Mux_s3_v I__309 (
            .O(N__2789),
            .I(N__2786));
    Odrv4 I__308 (
            .O(N__2786),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__307 (
            .O(N__2783),
            .I(N__2780));
    LocalMux I__306 (
            .O(N__2780),
            .I(N__2777));
    Span4Mux_v I__305 (
            .O(N__2777),
            .I(N__2774));
    Span4Mux_h I__304 (
            .O(N__2774),
            .I(N__2771));
    Span4Mux_h I__303 (
            .O(N__2771),
            .I(N__2768));
    Span4Mux_v I__302 (
            .O(N__2768),
            .I(N__2765));
    Odrv4 I__301 (
            .O(N__2765),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__300 (
            .O(N__2762),
            .I(N__2759));
    LocalMux I__299 (
            .O(N__2759),
            .I(N__2756));
    Span4Mux_s0_h I__298 (
            .O(N__2756),
            .I(N__2753));
    Sp12to4 I__297 (
            .O(N__2753),
            .I(N__2750));
    Span12Mux_s8_v I__296 (
            .O(N__2750),
            .I(N__2747));
    Span12Mux_h I__295 (
            .O(N__2747),
            .I(N__2744));
    Odrv12 I__294 (
            .O(N__2744),
            .I(un1_D_LL_AMIGA_0));
    InMux I__293 (
            .O(N__2741),
            .I(N__2738));
    LocalMux I__292 (
            .O(N__2738),
            .I(N__2735));
    Span4Mux_v I__291 (
            .O(N__2735),
            .I(N__2732));
    Sp12to4 I__290 (
            .O(N__2732),
            .I(N__2729));
    Span12Mux_h I__289 (
            .O(N__2729),
            .I(N__2726));
    Odrv12 I__288 (
            .O(N__2726),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__287 (
            .O(N__2723),
            .I(N__2720));
    LocalMux I__286 (
            .O(N__2720),
            .I(N__2717));
    Span4Mux_s3_h I__285 (
            .O(N__2717),
            .I(N__2714));
    Sp12to4 I__284 (
            .O(N__2714),
            .I(N__2711));
    Span12Mux_s8_v I__283 (
            .O(N__2711),
            .I(N__2708));
    Span12Mux_h I__282 (
            .O(N__2708),
            .I(N__2705));
    Odrv12 I__281 (
            .O(N__2705),
            .I(un1_D_LL_AMIGA_1));
    InMux I__280 (
            .O(N__2702),
            .I(N__2699));
    LocalMux I__279 (
            .O(N__2699),
            .I(N__2696));
    Span12Mux_v I__278 (
            .O(N__2696),
            .I(N__2693));
    Odrv12 I__277 (
            .O(N__2693),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__276 (
            .O(N__2690),
            .I(N__2687));
    LocalMux I__275 (
            .O(N__2687),
            .I(N__2684));
    Span12Mux_s8_h I__274 (
            .O(N__2684),
            .I(N__2681));
    Span12Mux_h I__273 (
            .O(N__2681),
            .I(N__2678));
    Odrv12 I__272 (
            .O(N__2678),
            .I(un1_D_LL_AMIGA_3));
    InMux I__271 (
            .O(N__2675),
            .I(N__2672));
    LocalMux I__270 (
            .O(N__2672),
            .I(N__2669));
    Span4Mux_v I__269 (
            .O(N__2669),
            .I(N__2666));
    Sp12to4 I__268 (
            .O(N__2666),
            .I(N__2663));
    Span12Mux_h I__267 (
            .O(N__2663),
            .I(N__2660));
    Odrv12 I__266 (
            .O(N__2660),
            .I(D_UM_040_in_6));
    IoInMux I__265 (
            .O(N__2657),
            .I(N__2654));
    LocalMux I__264 (
            .O(N__2654),
            .I(N__2651));
    IoSpan4Mux I__263 (
            .O(N__2651),
            .I(N__2647));
    InMux I__262 (
            .O(N__2650),
            .I(N__2644));
    IoSpan4Mux I__261 (
            .O(N__2647),
            .I(N__2641));
    LocalMux I__260 (
            .O(N__2644),
            .I(N__2638));
    Span4Mux_s2_h I__259 (
            .O(N__2641),
            .I(N__2635));
    Span4Mux_v I__258 (
            .O(N__2638),
            .I(N__2632));
    Sp12to4 I__257 (
            .O(N__2635),
            .I(N__2629));
    Sp12to4 I__256 (
            .O(N__2632),
            .I(N__2626));
    Span12Mux_h I__255 (
            .O(N__2629),
            .I(N__2623));
    Span12Mux_h I__254 (
            .O(N__2626),
            .I(N__2620));
    Span12Mux_h I__253 (
            .O(N__2623),
            .I(N__2615));
    Span12Mux_v I__252 (
            .O(N__2620),
            .I(N__2615));
    Odrv12 I__251 (
            .O(N__2615),
            .I(D_LL_040_in_6));
    IoInMux I__250 (
            .O(N__2612),
            .I(N__2609));
    LocalMux I__249 (
            .O(N__2609),
            .I(N__2606));
    Span12Mux_s8_h I__248 (
            .O(N__2606),
            .I(N__2603));
    Span12Mux_v I__247 (
            .O(N__2603),
            .I(N__2600));
    Odrv12 I__246 (
            .O(N__2600),
            .I(un1_D_UM_040_6));
    IoInMux I__245 (
            .O(N__2597),
            .I(N__2594));
    LocalMux I__244 (
            .O(N__2594),
            .I(N__2591));
    Span4Mux_s3_v I__243 (
            .O(N__2591),
            .I(N__2588));
    Span4Mux_h I__242 (
            .O(N__2588),
            .I(N__2585));
    Sp12to4 I__241 (
            .O(N__2585),
            .I(N__2582));
    Odrv12 I__240 (
            .O(N__2582),
            .I(LBENn_c_i));
    InMux I__239 (
            .O(N__2579),
            .I(N__2576));
    LocalMux I__238 (
            .O(N__2576),
            .I(N__2573));
    Span12Mux_v I__237 (
            .O(N__2573),
            .I(N__2570));
    Odrv12 I__236 (
            .O(N__2570),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__235 (
            .O(N__2567),
            .I(N__2564));
    LocalMux I__234 (
            .O(N__2564),
            .I(N__2561));
    IoSpan4Mux I__233 (
            .O(N__2561),
            .I(N__2558));
    IoSpan4Mux I__232 (
            .O(N__2558),
            .I(N__2555));
    Sp12to4 I__231 (
            .O(N__2555),
            .I(N__2552));
    Span12Mux_s9_h I__230 (
            .O(N__2552),
            .I(N__2549));
    Odrv12 I__229 (
            .O(N__2549),
            .I(un1_D_LM_AMIGA_4));
    IoInMux I__228 (
            .O(N__2546),
            .I(N__2543));
    LocalMux I__227 (
            .O(N__2543),
            .I(N__2540));
    Span4Mux_s0_v I__226 (
            .O(N__2540),
            .I(N__2537));
    Sp12to4 I__225 (
            .O(N__2537),
            .I(N__2534));
    Span12Mux_h I__224 (
            .O(N__2534),
            .I(N__2531));
    Span12Mux_v I__223 (
            .O(N__2531),
            .I(N__2528));
    Span12Mux_v I__222 (
            .O(N__2528),
            .I(N__2525));
    Odrv12 I__221 (
            .O(N__2525),
            .I(TAn_in));
    IoInMux I__220 (
            .O(N__2522),
            .I(N__2519));
    LocalMux I__219 (
            .O(N__2519),
            .I(N__2516));
    Span4Mux_s0_h I__218 (
            .O(N__2516),
            .I(N__2513));
    Span4Mux_h I__217 (
            .O(N__2513),
            .I(N__2510));
    Span4Mux_h I__216 (
            .O(N__2510),
            .I(N__2507));
    Sp12to4 I__215 (
            .O(N__2507),
            .I(N__2504));
    Span12Mux_v I__214 (
            .O(N__2504),
            .I(N__2501));
    Span12Mux_v I__213 (
            .O(N__2501),
            .I(N__2498));
    Span12Mux_h I__212 (
            .O(N__2498),
            .I(N__2495));
    Odrv12 I__211 (
            .O(N__2495),
            .I(TCIn_c));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__7753));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2  (
            .in0(N__5050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2825),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_7  (
            .in0(_gnd_net_),
            .in1(N__3625),
            .in2(_gnd_net_),
            .in3(N__5051),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_3_0  (
            .in0(N__6919),
            .in1(N__3359),
            .in2(_gnd_net_),
            .in3(N__2783),
            .lcout(un1_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_3  (
            .in0(N__2741),
            .in1(N__3284),
            .in2(_gnd_net_),
            .in3(N__6917),
            .lcout(un1_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_8_3_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_8_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_8_3_4  (
            .in0(N__6918),
            .in1(N__6053),
            .in2(_gnd_net_),
            .in3(N__2702),
            .lcout(un1_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_7  (
            .in0(N__6898),
            .in1(N__2675),
            .in2(_gnd_net_),
            .in3(N__2650),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BUFENn_obuf_RNO_LC_8_13_3.C_ON=1'b0;
    defparam BUFENn_obuf_RNO_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam BUFENn_obuf_RNO_LC_8_13_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 BUFENn_obuf_RNO_LC_8_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5447),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_5  (
            .in0(N__6899),
            .in1(N__6563),
            .in2(_gnd_net_),
            .in3(N__2579),
            .lcout(un1_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_15_0  (
            .in0(N__6935),
            .in1(N__6727),
            .in2(_gnd_net_),
            .in3(N__3215),
            .lcout(un1_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_8_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_8_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_8_15_2  (
            .in0(N__6937),
            .in1(N__5181),
            .in2(_gnd_net_),
            .in3(N__3179),
            .lcout(un1_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_5  (
            .in0(N__3152),
            .in1(N__4998),
            .in2(_gnd_net_),
            .in3(N__6936),
            .lcout(un1_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_20_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_20_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_20_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_8_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_8_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_8_20_3  (
            .in0(N__3082),
            .in1(N__3053),
            .in2(_gnd_net_),
            .in3(N__6920),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_9_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_9_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_9_11_1  (
            .in0(N__6881),
            .in1(N__6119),
            .in2(_gnd_net_),
            .in3(N__3014),
            .lcout(un1_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_11_5  (
            .in0(N__6880),
            .in1(N__2981),
            .in2(_gnd_net_),
            .in3(N__2962),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_5  (
            .in0(N__6944),
            .in1(N__2906),
            .in2(_gnd_net_),
            .in3(N__2881),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_9_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_9_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_9_20_0  (
            .in0(N__6948),
            .in1(N__3569),
            .in2(_gnd_net_),
            .in3(N__3541),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_6  (
            .in0(N__6947),
            .in1(N__3494),
            .in2(_gnd_net_),
            .in3(N__3469),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_10_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_10_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_10_10_5  (
            .in0(N__7136),
            .in1(N__3317),
            .in2(_gnd_net_),
            .in3(N__3352),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_10_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_10_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_10_10_6  (
            .in0(N__3395),
            .in1(N__3914),
            .in2(_gnd_net_),
            .in3(N__6790),
            .lcout(un1_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_10_11_4 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_10_11_4  (
            .in0(N__5315),
            .in1(N__6481),
            .in2(N__5389),
            .in3(N__4775),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7751),
            .ce(),
            .sr(N__7695));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_10_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_10_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_10_12_7  (
            .in0(N__3339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7748),
            .ce(N__6306),
            .sr(N__6246));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_10_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_10_13_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_10_13_1  (
            .in0(N__3277),
            .in1(N__7187),
            .in2(_gnd_net_),
            .in3(N__3245),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_10_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3276),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7742),
            .ce(N__6288),
            .sr(N__6243));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_14_6  (
            .in0(N__7188),
            .in1(N__3881),
            .in2(_gnd_net_),
            .in3(N__3910),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_14_7  (
            .in0(N__3909),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7740),
            .ce(N__6307),
            .sr(N__6247));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_10_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_10_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_10_20_1  (
            .in0(N__6946),
            .in1(N__3875),
            .in2(_gnd_net_),
            .in3(N__3856),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_10_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_10_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_10_20_6  (
            .in0(N__3802),
            .in1(N__3758),
            .in2(_gnd_net_),
            .in3(N__6945),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_3.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_3.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_3 (
            .in0(N__5428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_11_6_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_11_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_11_6_1  (
            .in0(N__3710),
            .in1(N__7268),
            .in2(_gnd_net_),
            .in3(N__6834),
            .lcout(un1_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_11_6_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_11_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_11_6_3  (
            .in0(N__3671),
            .in1(N__4844),
            .in2(_gnd_net_),
            .in3(N__6833),
            .lcout(un1_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__6435),
            .in2(_gnd_net_),
            .in3(N__3632),
            .lcout(\U111_CYCLE_SM.FLIP_WORD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3  (
            .in0(N__3608),
            .in1(N__5902),
            .in2(_gnd_net_),
            .in3(N__6832),
            .lcout(un1_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_7  (
            .in0(N__4436),
            .in1(N__4943),
            .in2(_gnd_net_),
            .in3(N__6831),
            .lcout(un1_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_11_9_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_11_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5637),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_11_9_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_11_9_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__5638),
            .in2(_gnd_net_),
            .in3(N__4096),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNIDDAN_LC_11_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNIDDAN_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNIDDAN_LC_11_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNIDDAN_LC_11_9_7  (
            .in0(N__7775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5446),
            .lcout(D_UU_AMIGA_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_11_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_11_10_0 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_11_10_0  (
            .in0(N__4759),
            .in1(N__7809),
            .in2(N__7158),
            .in3(N__4463),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7752),
            .ce(),
            .sr(N__7691));
    defparam \U111_CYCLE_SM.TS_EN_LC_11_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_11_10_5 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_11_10_5  (
            .in0(N__4766),
            .in1(N__5015),
            .in2(N__4103),
            .in3(N__4760),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7752),
            .ce(),
            .sr(N__7691));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_11_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_11_10_7 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_11_10_7  (
            .in0(N__6789),
            .in1(N__5313),
            .in2(N__4085),
            .in3(N__6470),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7752),
            .ce(),
            .sr(N__7691));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_11_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_11_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_11_11_1  (
            .in0(N__4073),
            .in1(N__4051),
            .in2(_gnd_net_),
            .in3(N__6791),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_11_11_2.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_11_11_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_11_11_2 (
            .in0(N__7757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_11_3  (
            .in0(N__6436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6500),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCH_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_11_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__5266),
            .in2(_gnd_net_),
            .in3(N__7496),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_123_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_11_5 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_11_5  (
            .in0(N__7805),
            .in1(N__5349),
            .in2(N__4769),
            .in3(N__7443),
            .lcout(\U111_CYCLE_SM.N_121_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNISO2G_3_LC_11_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNISO2G_3_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNISO2G_3_LC_11_11_7 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNISO2G_3_LC_11_11_7  (
            .in0(N__7806),
            .in1(N__7921),
            .in2(_gnd_net_),
            .in3(N__5306),
            .lcout(\U111_CYCLE_SM.un1_CYCLE_STATE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_12_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_12_1  (
            .in0(N__7922),
            .in1(N__7811),
            .in2(N__7872),
            .in3(N__4461),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7743),
            .ce(),
            .sr(N__7684));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIUBHI_LC_11_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIUBHI_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIUBHI_LC_11_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIUBHI_LC_11_12_4  (
            .in0(N__4462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(D_UU_040_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_11_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_11_13_0 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_11_13_0  (
            .in0(N__5657),
            .in1(N__4457),
            .in2(_gnd_net_),
            .in3(N__6328),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81 ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_11_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_11_13_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_11_13_1  (
            .in0(N__6329),
            .in1(_gnd_net_),
            .in2(N__4439),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_11_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5903),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_11_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5524),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_11_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_11_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_11_14_2  (
            .in0(N__4837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_11_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5000),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_11_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5192),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_14_7  (
            .in0(N__4936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7738),
            .ce(N__6302),
            .sr(N__6245));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_11_16_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_11_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_11_16_3  (
            .in0(N__7171),
            .in1(N__5009),
            .in2(_gnd_net_),
            .in3(N__4999),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_16_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_16_4  (
            .in0(N__4935),
            .in1(N__4907),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_11_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_11_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_11_20_1  (
            .in0(N__7192),
            .in1(N__4877),
            .in2(_gnd_net_),
            .in3(N__5511),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_11_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_11_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_11_20_3  (
            .in0(N__7191),
            .in1(N__4853),
            .in2(_gnd_net_),
            .in3(N__4824),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_11_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_11_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_11_20_7  (
            .in0(N__7193),
            .in1(N__5204),
            .in2(_gnd_net_),
            .in3(N__5191),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_0  (
            .in0(N__7406),
            .in1(N__5129),
            .in2(_gnd_net_),
            .in3(N__6915),
            .lcout(un1_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_12_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_12_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_12_3_7  (
            .in0(N__6916),
            .in1(N__6203),
            .in2(_gnd_net_),
            .in3(N__5087),
            .lcout(un1_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_LC_12_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_12_9_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_12_9_7  (
            .in0(N__5035),
            .in1(N__5024),
            .in2(_gnd_net_),
            .in3(N__5314),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7750),
            .ce(),
            .sr(N__7699));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_10_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_10_0  (
            .in0(N__7541),
            .in1(N__5264),
            .in2(_gnd_net_),
            .in3(N__5350),
            .lcout(\U111_CYCLE_SM.N_148 ),
            .ltout(\U111_CYCLE_SM.N_148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_10_1 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_10_1  (
            .in0(N__7585),
            .in1(N__6352),
            .in2(N__5018),
            .in3(N__5639),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_10_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_10_2  (
            .in0(N__5304),
            .in1(N__6463),
            .in2(N__5462),
            .in3(N__7584),
            .lcout(\U111_CYCLE_SM.TS_EN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__5640),
            .in2(_gnd_net_),
            .in3(N__5305),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_10_5  (
            .in0(N__5265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7542),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_10_6 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_10_6  (
            .in0(N__5461),
            .in1(N__5641),
            .in2(N__5450),
            .in3(N__5351),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7744),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNITIC9_0_LC_12_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNITIC9_0_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNITIC9_0_LC_12_11_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNITIC9_0_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__7916),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__5348),
            .in2(_gnd_net_),
            .in3(N__7444),
            .lcout(\U111_CYCLE_SM.N_128_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_11_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_11_2  (
            .in0(N__5432),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5393),
            .lcout(TAn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_11_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_11_3  (
            .in0(N__7543),
            .in1(N__5347),
            .in2(_gnd_net_),
            .in3(N__7582),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_11_4 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_11_4  (
            .in0(N__5655),
            .in1(N__7917),
            .in2(N__5327),
            .in3(N__7808),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_11_5 .LUT_INIT=16'b1111111100011111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_11_5  (
            .in0(N__5267),
            .in1(N__5324),
            .in2(N__5318),
            .in3(N__7418),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7741),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_11_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_11_7  (
            .in0(N__5654),
            .in1(N__6330),
            .in2(_gnd_net_),
            .in3(N__7472),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7741),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_12_0  (
            .in0(N__7544),
            .in1(N__5268),
            .in2(_gnd_net_),
            .in3(N__7441),
            .lcout(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_3 .LUT_INIT=16'b0101110101011111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_3  (
            .in0(N__5269),
            .in1(N__7470),
            .in2(N__7552),
            .in3(N__7559),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_4 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_4  (
            .in0(N__5656),
            .in1(N__6477),
            .in2(N__5591),
            .in3(N__7442),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7739),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5588),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_12_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_12_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_12_12_7  (
            .in0(N__5537),
            .in1(N__5525),
            .in2(_gnd_net_),
            .in3(N__6846),
            .lcout(un1_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_13_6  (
            .in0(N__7398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7737),
            .ce(N__6295),
            .sr(N__6244));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_14_0  (
            .in0(N__7263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_14_1  (
            .in0(N__6562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_12_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_12_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6728),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6052),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_14_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6118),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_6  (
            .in0(N__6193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7736),
            .ce(N__6308),
            .sr(N__6248));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_17_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_17_3  (
            .in0(N__6186),
            .in1(N__6158),
            .in2(_gnd_net_),
            .in3(N__7207),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_17_5  (
            .in0(N__6128),
            .in1(N__6108),
            .in2(_gnd_net_),
            .in3(N__7208),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_18_0  (
            .in0(N__7209),
            .in1(N__6062),
            .in2(_gnd_net_),
            .in3(N__6045),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_12_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_12_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_12_18_7  (
            .in0(N__5981),
            .in1(N__5956),
            .in2(_gnd_net_),
            .in3(N__6949),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_1  (
            .in0(N__5892),
            .in1(N__5855),
            .in2(_gnd_net_),
            .in3(N__7218),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_12_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_12_19_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_12_19_2  (
            .in0(N__6932),
            .in1(N__5819),
            .in2(_gnd_net_),
            .in3(N__5798),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_12_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_12_19_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_12_19_3  (
            .in0(N__5732),
            .in1(N__5701),
            .in2(_gnd_net_),
            .in3(N__6933),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_12_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_12_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_12_20_1  (
            .in0(N__7220),
            .in1(N__6737),
            .in2(_gnd_net_),
            .in3(N__6717),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_4  (
            .in0(N__6655),
            .in1(N__6934),
            .in2(_gnd_net_),
            .in3(N__6614),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_20_7  (
            .in0(N__7219),
            .in1(N__6572),
            .in2(_gnd_net_),
            .in3(N__6549),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_13_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_13_11_0 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_13_11_0  (
            .in0(N__7649),
            .in1(N__7637),
            .in2(N__6359),
            .in3(N__6332),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_13_11_1 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_13_11_1  (
            .in0(N__6379),
            .in1(N__6498),
            .in2(N__6401),
            .in3(N__6358),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_2  (
            .in0(N__6499),
            .in1(N__7471),
            .in2(N__6482),
            .in3(N__6437),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.BURST_LC_13_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_13_11_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_13_11_3  (
            .in0(N__6397),
            .in1(N__6357),
            .in2(N__6380),
            .in3(N__7586),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_13_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_13_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_13_11_4  (
            .in0(N__6353),
            .in1(N__7636),
            .in2(_gnd_net_),
            .in3(N__6331),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_13_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_13_11_6 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_13_11_6  (
            .in0(N__7915),
            .in1(N__7768),
            .in2(N__7873),
            .in3(N__7810),
            .lcout(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7749),
            .ce(),
            .sr(N__7700));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_13_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_13_12_6 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_13_12_6  (
            .in0(N__7648),
            .in1(N__7635),
            .in2(N__7622),
            .in3(N__7583),
            .lcout(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ),
            .ltout(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_13_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_13_12_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_13_12_7  (
            .in0(N__7548),
            .in1(N__7469),
            .in2(N__7448),
            .in3(N__7445),
            .lcout(\U111_CYCLE_SM.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_13_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_13_5  (
            .in0(N__7412),
            .in1(N__7399),
            .in2(_gnd_net_),
            .in3(N__7189),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_14_0  (
            .in0(N__7352),
            .in1(N__6921),
            .in2(_gnd_net_),
            .in3(N__7333),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_14_1  (
            .in0(N__7264),
            .in1(N__7226),
            .in2(_gnd_net_),
            .in3(N__7190),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_13_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_13_20_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_13_20_1  (
            .in0(N__7082),
            .in1(N__6956),
            .in2(_gnd_net_),
            .in3(N__7060),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_13_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_13_20_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_13_20_3  (
            .in0(N__6991),
            .in1(N__6955),
            .in2(_gnd_net_),
            .in3(N__7961),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

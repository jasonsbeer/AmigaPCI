-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 13 2024 16:29:06

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    A : in std_logic_vector(31 downto 1);
    RnW : in std_logic;
    TT1 : in std_logic;
    TICK50 : out std_logic;
    nROMEN : out std_logic;
    nCIACS1 : out std_logic;
    TT0 : in std_logic;
    TICK60 : out std_logic;
    LBENn : in std_logic;
    CLKCIA : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    TSn : in std_logic;
    nBUFEN : out std_logic;
    nREGSPACE : out std_logic;
    nRAMSPACE : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    nCIACS0 : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2369\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_CIA.g0Z0Z_11_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_8\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_CIA.g0Z0Z_10_cascade_\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_CIA.g0Z0Z_2\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\ : std_logic;
signal \A_c_21\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nREGSPACE_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un10_ROMENZ0\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \U409_TICK.TICK603_11_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\ : std_logic;
signal \nBUFEN_c\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS1_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS0_i\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_97_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_97\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un6_ROMENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ROMEN_0\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_347_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \nCIACS0_wire\ : std_logic;
signal \nCIACS1_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \nRAMSPACE_wire\ : std_logic;
signal \nROMEN_wire\ : std_logic;
signal \nBUFEN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \nREGSPACE_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    nCIACS0 <= \nCIACS0_wire\;
    nCIACS1 <= \nCIACS1_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    nRAMSPACE <= \nRAMSPACE_wire\;
    nROMEN <= \nROMEN_wire\;
    nBUFEN <= \nBUFEN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    nREGSPACE <= \nREGSPACE_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4970\,
            RESETB => \N__5222\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6034\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6036\,
            DIN => \N__6035\,
            DOUT => \N__6034\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6036\,
            PADOUT => \N__6035\,
            PADIN => \N__6034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6024\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6026\,
            DIN => \N__6025\,
            DOUT => \N__6024\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6026\,
            PADOUT => \N__6025\,
            PADIN => \N__6024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6015\,
            DIN => \N__6014\,
            DOUT => \N__6013\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6015\,
            PADOUT => \N__6014\,
            PADIN => \N__6013\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4658\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6006\,
            DIN => \N__6005\,
            DOUT => \N__6004\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6006\,
            PADOUT => \N__6005\,
            PADIN => \N__6004\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5997\,
            DIN => \N__5996\,
            DOUT => \N__5995\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5997\,
            PADOUT => \N__5996\,
            PADIN => \N__5995\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5988\,
            DIN => \N__5987\,
            DOUT => \N__5986\,
            PACKAGEPIN => \nCIACS0_wire\
        );

    \nCIACS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5988\,
            PADOUT => \N__5987\,
            PADIN => \N__5986\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5979\,
            DIN => \N__5978\,
            DOUT => \N__5977\,
            PACKAGEPIN => \nCIACS1_wire\
        );

    \nCIACS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5979\,
            PADOUT => \N__5978\,
            PADIN => \N__5977\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3275\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5970\,
            DIN => \N__5969\,
            DOUT => \N__5968\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5970\,
            PADOUT => \N__5969\,
            PADIN => \N__5968\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5961\,
            DIN => \N__5960\,
            DOUT => \N__5959\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5961\,
            PADOUT => \N__5960\,
            PADIN => \N__5959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5952\,
            DIN => \N__5951\,
            DOUT => \N__5950\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5952\,
            PADOUT => \N__5951\,
            PADIN => \N__5950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5943\,
            DIN => \N__5942\,
            DOUT => \N__5941\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__5943\,
            PADOUT => \N__5942\,
            PADIN => \N__5941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5372\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5934\,
            DIN => \N__5933\,
            DOUT => \N__5932\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5934\,
            PADOUT => \N__5933\,
            PADIN => \N__5932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5925\,
            DIN => \N__5924\,
            DOUT => \N__5923\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5925\,
            PADOUT => \N__5924\,
            PADIN => \N__5923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5916\,
            DIN => \N__5915\,
            DOUT => \N__5914\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5916\,
            PADOUT => \N__5915\,
            PADIN => \N__5914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nRAMSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5907\,
            DIN => \N__5906\,
            DOUT => \N__5905\,
            PACKAGEPIN => \nRAMSPACE_wire\
        );

    \nRAMSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5907\,
            PADOUT => \N__5906\,
            PADIN => \N__5905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4799\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nROMEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5898\,
            DIN => \N__5897\,
            DOUT => \N__5896\,
            PACKAGEPIN => \nROMEN_wire\
        );

    \nROMEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5898\,
            PADOUT => \N__5897\,
            PADIN => \N__5896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5889\,
            DIN => \N__5888\,
            DOUT => \N__5887\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5889\,
            PADOUT => \N__5888\,
            PADIN => \N__5887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5880\,
            DIN => \N__5879\,
            DOUT => \N__5878\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5880\,
            PADOUT => \N__5879\,
            PADIN => \N__5878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nBUFEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5871\,
            DIN => \N__5870\,
            DOUT => \N__5869\,
            PACKAGEPIN => \nBUFEN_wire\
        );

    \nBUFEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5871\,
            PADOUT => \N__5870\,
            PADIN => \N__5869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3113\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5862\,
            DIN => \N__5861\,
            DOUT => \N__5860\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5862\,
            PADOUT => \N__5861\,
            PADIN => \N__5860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5853\,
            DIN => \N__5852\,
            DOUT => \N__5851\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5853\,
            PADOUT => \N__5852\,
            PADIN => \N__5851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5844\,
            DIN => \N__5843\,
            DOUT => \N__5842\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5844\,
            PADOUT => \N__5843\,
            PADIN => \N__5842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5835\,
            DIN => \N__5834\,
            DOUT => \N__5833\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5835\,
            PADOUT => \N__5834\,
            PADIN => \N__5833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5826\,
            DIN => \N__5825\,
            DOUT => \N__5824\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5826\,
            PADOUT => \N__5825\,
            PADIN => \N__5824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5817\,
            DIN => \N__5816\,
            DOUT => \N__5815\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5817\,
            PADOUT => \N__5816\,
            PADIN => \N__5815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5808\,
            DIN => \N__5807\,
            DOUT => \N__5806\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5808\,
            PADOUT => \N__5807\,
            PADIN => \N__5806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nREGSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5799\,
            DIN => \N__5798\,
            DOUT => \N__5797\,
            PACKAGEPIN => \nREGSPACE_wire\
        );

    \nREGSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5799\,
            PADOUT => \N__5798\,
            PADIN => \N__5797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5790\,
            DIN => \N__5789\,
            DOUT => \N__5788\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5790\,
            PADOUT => \N__5789\,
            PADIN => \N__5788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4346\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5781\,
            DIN => \N__5780\,
            DOUT => \N__5779\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5781\,
            PADOUT => \N__5780\,
            PADIN => \N__5779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5772\,
            DIN => \N__5771\,
            DOUT => \N__5770\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5772\,
            PADOUT => \N__5771\,
            PADIN => \N__5770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5763\,
            DIN => \N__5762\,
            DOUT => \N__5761\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5763\,
            PADOUT => \N__5762\,
            PADIN => \N__5761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5754\,
            DIN => \N__5753\,
            DOUT => \N__5752\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5754\,
            PADOUT => \N__5753\,
            PADIN => \N__5752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5745\,
            DIN => \N__5744\,
            DOUT => \N__5743\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5745\,
            PADOUT => \N__5744\,
            PADIN => \N__5743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5736\,
            DIN => \N__5735\,
            DOUT => \N__5734\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5736\,
            PADOUT => \N__5735\,
            PADIN => \N__5734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3587\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5727\,
            DIN => \N__5726\,
            DOUT => \N__5725\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5727\,
            PADOUT => \N__5726\,
            PADIN => \N__5725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1319\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5702\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5702\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__5699\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5689\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5684\
        );

    \I__1313\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5684\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5679\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5692\,
            I => \N__5679\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5689\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5684\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5679\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5661\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5661\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5658\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5649\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5649\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5649\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5649\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5658\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__5649\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__5642\,
            I => \N__5637\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5633\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5630\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5625\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5625\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5633\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5630\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5625\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5615\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__5612\,
            I => \N__5608\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5601\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5605\,
            I => \N__5596\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__5604\,
            I => \N__5593\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5601\,
            I => \N__5587\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__5600\,
            I => \N__5584\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__5599\,
            I => \N__5580\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__5596\,
            I => \N__5573\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5570\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5563\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5563\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5563\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__5587\,
            I => \N__5559\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5554\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5554\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5549\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5549\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5546\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5543\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5538\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__5573\,
            I => \N__5532\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5527\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5527\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5524\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__5559\,
            I => \N__5520\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5517\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5514\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5546\,
            I => \N__5509\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5509\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5504\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5504\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5497\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5497\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5497\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5494\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__5532\,
            I => \N__5487\
        );

    \I__1250\ : Span4Mux_v
    port map (
            O => \N__5527\,
            I => \N__5487\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5524\,
            I => \N__5487\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5484\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__5520\,
            I => \N__5469\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__5517\,
            I => \N__5469\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__5514\,
            I => \N__5469\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__5509\,
            I => \N__5469\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5469\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5469\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5469\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__5487\,
            I => \N__5466\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5484\,
            I => \N__5463\
        );

    \I__1238\ : Span4Mux_v
    port map (
            O => \N__5469\,
            I => \N__5460\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__5466\,
            I => \N__5455\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__5463\,
            I => \N__5455\
        );

    \I__1235\ : Sp12to4
    port map (
            O => \N__5460\,
            I => \N__5450\
        );

    \I__1234\ : Sp12to4
    port map (
            O => \N__5455\,
            I => \N__5450\
        );

    \I__1233\ : Span12Mux_h
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__1232\ : Span12Mux_v
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__1231\ : Odrv12
    port map (
            O => \N__5444\,
            I => \RESETn_c\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__1227\ : Sp12to4
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__1226\ : Span12Mux_h
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__1225\ : Span12Mux_v
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__1224\ : Odrv12
    port map (
            O => \N__5423\,
            I => \TACKn_in\
        );

    \I__1223\ : SRMux
    port map (
            O => \N__5420\,
            I => \N__5415\
        );

    \I__1222\ : SRMux
    port map (
            O => \N__5419\,
            I => \N__5412\
        );

    \I__1221\ : SRMux
    port map (
            O => \N__5418\,
            I => \N__5409\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5415\,
            I => \N__5406\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5403\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5409\,
            I => \N__5400\
        );

    \I__1217\ : Span12Mux_h
    port map (
            O => \N__5406\,
            I => \N__5397\
        );

    \I__1216\ : Span4Mux_h
    port map (
            O => \N__5403\,
            I => \N__5394\
        );

    \I__1215\ : Span4Mux_h
    port map (
            O => \N__5400\,
            I => \N__5391\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__5397\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__5394\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__5391\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__5375\,
            I => \TACK_EN_i\
        );

    \I__1207\ : IoInMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__1205\ : IoSpan4Mux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__1204\ : Sp12to4
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__1203\ : Span12Mux_v
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1202\ : Span12Mux_h
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__1201\ : Odrv12
    port map (
            O => \N__5354\,
            I => \N_347_i\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5346\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5342\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5339\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5336\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5332\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5342\,
            I => \N__5327\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5339\,
            I => \N__5327\
        );

    \I__1193\ : Span4Mux_h
    port map (
            O => \N__5336\,
            I => \N__5323\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5319\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5316\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__5327\,
            I => \N__5313\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5310\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__5323\,
            I => \N__5307\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5304\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5319\,
            I => \N__5301\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__5316\,
            I => \N__5298\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__5313\,
            I => \N__5293\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5293\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__5307\,
            I => \N__5288\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5304\,
            I => \N__5288\
        );

    \I__1180\ : Span12Mux_v
    port map (
            O => \N__5301\,
            I => \N__5285\
        );

    \I__1179\ : Span4Mux_v
    port map (
            O => \N__5298\,
            I => \N__5282\
        );

    \I__1178\ : Span4Mux_h
    port map (
            O => \N__5293\,
            I => \N__5279\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__5288\,
            I => \N__5276\
        );

    \I__1176\ : Odrv12
    port map (
            O => \N__5285\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__5282\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__5279\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__5276\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5263\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5260\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5257\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5254\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__5251\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__5248\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__1164\ : IoInMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__1162\ : Span4Mux_s1_v
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__1160\ : Span12Mux_h
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__5225\,
            I => \ROMENm_i\
        );

    \I__1157\ : IoInMux
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__1155\ : Span4Mux_s2_v
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__5210\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5198\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5198\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5198\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__5195\,
            I => \N__5189\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5185\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5178\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5178\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5178\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5175\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5178\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__5168\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__5165\,
            I => \N__5161\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5158\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5139\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5139\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5139\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5136\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5133\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5139\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5133\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__5126\,
            I => \N__5121\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5117\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5114\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5109\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5109\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5109\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5093\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5090\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5085\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5085\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5090\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5085\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5073\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5068\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5068\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5073\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5068\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__5063\,
            I => \N__5057\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5052\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5052\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5047\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5047\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5052\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5047\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__5042\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5032\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5029\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5032\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5029\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__5015\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__5005\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5001\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__5005\,
            I => \N__4998\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4995\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5001\,
            I => \N__4992\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__4998\,
            I => \N__4987\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4987\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__4992\,
            I => \N__4984\
        );

    \I__1078\ : Span12Mux_h
    port map (
            O => \N__4987\,
            I => \N__4981\
        );

    \I__1077\ : Span12Mux_v
    port map (
            O => \N__4984\,
            I => \N__4978\
        );

    \I__1076\ : Span12Mux_v
    port map (
            O => \N__4981\,
            I => \N__4975\
        );

    \I__1075\ : Odrv12
    port map (
            O => \N__4978\,
            I => \TSn_c\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__4975\,
            I => \TSn_c\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__4970\,
            I => \N__4962\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__4969\,
            I => \N__4959\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__4968\,
            I => \N__4956\
        );

    \I__1070\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4953\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__4966\,
            I => \N__4950\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__4965\,
            I => \N__4947\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__4962\,
            I => \N__4944\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4939\
        );

    \I__1065\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4939\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4953\,
            I => \N__4936\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4933\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4930\
        );

    \I__1061\ : IoSpan4Mux
    port map (
            O => \N__4944\,
            I => \N__4927\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4924\
        );

    \I__1059\ : Span4Mux_h
    port map (
            O => \N__4936\,
            I => \N__4917\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__4933\,
            I => \N__4917\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__4930\,
            I => \N__4917\
        );

    \I__1056\ : Span4Mux_s0_v
    port map (
            O => \N__4927\,
            I => \N__4914\
        );

    \I__1055\ : Span4Mux_v
    port map (
            O => \N__4924\,
            I => \N__4911\
        );

    \I__1054\ : Span4Mux_v
    port map (
            O => \N__4917\,
            I => \N__4908\
        );

    \I__1053\ : Sp12to4
    port map (
            O => \N__4914\,
            I => \N__4905\
        );

    \I__1052\ : Sp12to4
    port map (
            O => \N__4911\,
            I => \N__4900\
        );

    \I__1051\ : Sp12to4
    port map (
            O => \N__4908\,
            I => \N__4900\
        );

    \I__1050\ : Span12Mux_v
    port map (
            O => \N__4905\,
            I => \N__4897\
        );

    \I__1049\ : Span12Mux_h
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__1048\ : Span12Mux_v
    port map (
            O => \N__4897\,
            I => \N__4891\
        );

    \I__1047\ : Span12Mux_v
    port map (
            O => \N__4894\,
            I => \N__4888\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__4891\,
            I => \CLK40_IN_c\
        );

    \I__1045\ : Odrv12
    port map (
            O => \N__4888\,
            I => \CLK40_IN_c\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4879\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4876\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4879\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4864\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4861\
        );

    \I__1037\ : Span4Mux_v
    port map (
            O => \N__4864\,
            I => \N__4857\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4861\,
            I => \N__4854\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4851\
        );

    \I__1034\ : Sp12to4
    port map (
            O => \N__4857\,
            I => \N__4846\
        );

    \I__1033\ : Span12Mux_v
    port map (
            O => \N__4854\,
            I => \N__4846\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4851\,
            I => \N__4843\
        );

    \I__1031\ : Span12Mux_v
    port map (
            O => \N__4846\,
            I => \N__4840\
        );

    \I__1030\ : Span12Mux_h
    port map (
            O => \N__4843\,
            I => \N__4837\
        );

    \I__1029\ : Span12Mux_h
    port map (
            O => \N__4840\,
            I => \N__4832\
        );

    \I__1028\ : Span12Mux_v
    port map (
            O => \N__4837\,
            I => \N__4832\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__4832\,
            I => \OVL_c\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4822\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__4825\,
            I => \N__4819\
        );

    \I__1023\ : Span4Mux_v
    port map (
            O => \N__4822\,
            I => \N__4815\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4812\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4809\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__4815\,
            I => \N__4802\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4802\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4802\
        );

    \I__1017\ : Odrv12
    port map (
            O => \N__4802\,
            I => \U409_ADDRESS_DECODE.un6_ROMENZ0\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__1014\ : IoSpan4Mux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__1013\ : Span4Mux_s2_v
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__1012\ : Sp12to4
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__1011\ : Span12Mux_v
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__4781\,
            I => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4774\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4771\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4774\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1005\ : CEMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__4760\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4742\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4742\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4742\
        );

    \I__999\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4742\
        );

    \I__998\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4735\
        );

    \I__997\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4735\
        );

    \I__996\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4735\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4742\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__4730\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__992\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \N__4711\
        );

    \I__989\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4708\
        );

    \I__988\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4699\
        );

    \I__987\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4699\
        );

    \I__986\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4699\
        );

    \I__985\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4699\
        );

    \I__984\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4692\
        );

    \I__983\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4692\
        );

    \I__982\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4692\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4708\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4699\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4692\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__4685\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__977\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4668\
        );

    \I__976\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4668\
        );

    \I__975\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4668\
        );

    \I__974\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4668\
        );

    \I__973\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4663\
        );

    \I__972\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4663\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4668\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4663\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__969\ : IoInMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__967\ : Span4Mux_s0_v
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__966\ : Sp12to4
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__965\ : Span12Mux_h
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__964\ : Span12Mux_v
    port map (
            O => \N__4643\,
            I => \N__4638\
        );

    \I__963\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4635\
        );

    \I__962\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4632\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__4638\,
            I => \CLKCIA_c\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4635\,
            I => \CLKCIA_c\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4632\,
            I => \CLKCIA_c\
        );

    \I__958\ : ClkMux
    port map (
            O => \N__4625\,
            I => \N__4613\
        );

    \I__957\ : ClkMux
    port map (
            O => \N__4624\,
            I => \N__4613\
        );

    \I__956\ : ClkMux
    port map (
            O => \N__4623\,
            I => \N__4613\
        );

    \I__955\ : ClkMux
    port map (
            O => \N__4622\,
            I => \N__4613\
        );

    \I__954\ : GlobalMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__953\ : gio2CtrlBuf
    port map (
            O => \N__4610\,
            I => \CLK28_IN_c_g\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__4607\,
            I => \N__4603\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__4606\,
            I => \N__4599\
        );

    \I__950\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4593\
        );

    \I__949\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4593\
        );

    \I__948\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4588\
        );

    \I__947\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4588\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4593\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4588\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__944\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__943\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4572\
        );

    \I__942\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4572\
        );

    \I__941\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4569\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4577\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4572\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4569\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__937\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4554\
        );

    \I__936\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4554\
        );

    \I__935\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4549\
        );

    \I__934\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4549\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4554\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4549\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__931\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4538\
        );

    \I__930\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4538\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__4535\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__4532\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__926\ : InMux
    port map (
            O => \N__4529\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__925\ : InMux
    port map (
            O => \N__4526\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__924\ : InMux
    port map (
            O => \N__4523\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__4520\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__922\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4514\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__919\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4502\
        );

    \I__918\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4502\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4502\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__4499\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__914\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4488\
        );

    \I__913\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4483\
        );

    \I__912\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4483\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4488\,
            I => \N__4480\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4476\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__4480\,
            I => \N__4473\
        );

    \I__908\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4470\
        );

    \I__907\ : Span4Mux_h
    port map (
            O => \N__4476\,
            I => \N__4467\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__4473\,
            I => \U409_CIA.VMAZ0\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4470\,
            I => \U409_CIA.VMAZ0\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__4467\,
            I => \U409_CIA.VMAZ0\
        );

    \I__903\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4452\
        );

    \I__902\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4452\
        );

    \I__901\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4447\
        );

    \I__900\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4447\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4452\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4447\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__897\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4439\,
            I => \N__4434\
        );

    \I__895\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4431\
        );

    \I__894\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4428\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__4434\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4431\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4428\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__890\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4417\
        );

    \I__889\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4414\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4417\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4414\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__886\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4406\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__4403\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__883\ : IoInMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__881\ : IoSpan4Mux
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__880\ : Span4Mux_s1_v
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__879\ : Sp12to4
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__878\ : Span12Mux_v
    port map (
            O => \N__4385\,
            I => \N__4381\
        );

    \I__877\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4378\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__4381\,
            I => \TACK_OUTn\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4378\,
            I => \TACK_OUTn\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__4373\,
            I => \N__4368\
        );

    \I__873\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4361\
        );

    \I__872\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4361\
        );

    \I__871\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4361\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4361\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__869\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4349\
        );

    \I__868\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4349\
        );

    \I__867\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4349\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4349\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__865\ : IoInMux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__863\ : Span4Mux_s2_v
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__860\ : Sp12to4
    port map (
            O => \N__4331\,
            I => \N__4327\
        );

    \I__859\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4324\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__4327\,
            I => \TICK50_c\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4324\,
            I => \TICK50_c\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__4319\,
            I => \N__4312\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__4318\,
            I => \N__4309\
        );

    \I__854\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4303\
        );

    \I__853\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4300\
        );

    \I__852\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4291\
        );

    \I__851\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4291\
        );

    \I__850\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4291\
        );

    \I__849\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4291\
        );

    \I__848\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4286\
        );

    \I__847\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4286\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4303\,
            I => \U409_TICK.TICK503_10\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4300\,
            I => \U409_TICK.TICK503_10\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4291\,
            I => \U409_TICK.TICK503_10\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4286\,
            I => \U409_TICK.TICK503_10\
        );

    \I__842\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4267\
        );

    \I__841\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4264\
        );

    \I__840\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4255\
        );

    \I__839\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4255\
        );

    \I__838\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4255\
        );

    \I__837\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4255\
        );

    \I__836\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4250\
        );

    \I__835\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4250\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4267\,
            I => \U409_TICK.TICK503_14\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4264\,
            I => \U409_TICK.TICK503_14\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4255\,
            I => \U409_TICK.TICK503_14\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4250\,
            I => \U409_TICK.TICK503_14\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__4241\,
            I => \N__4237\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__4240\,
            I => \N__4234\
        );

    \I__828\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4225\
        );

    \I__827\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4222\
        );

    \I__826\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4215\
        );

    \I__825\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4215\
        );

    \I__824\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4215\
        );

    \I__823\ : InMux
    port map (
            O => \N__4230\,
            I => \N__4208\
        );

    \I__822\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4208\
        );

    \I__821\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4208\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4225\,
            I => \U409_TICK.TICK503_9\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4222\,
            I => \U409_TICK.TICK503_9\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4215\,
            I => \U409_TICK.TICK503_9\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4208\,
            I => \U409_TICK.TICK503_9\
        );

    \I__816\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__814\ : Odrv4
    port map (
            O => \N__4193\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__813\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4186\
        );

    \I__812\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4183\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4186\,
            I => \N__4180\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4183\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__4180\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__808\ : ClkMux
    port map (
            O => \N__4175\,
            I => \N__4142\
        );

    \I__807\ : ClkMux
    port map (
            O => \N__4174\,
            I => \N__4142\
        );

    \I__806\ : ClkMux
    port map (
            O => \N__4173\,
            I => \N__4142\
        );

    \I__805\ : ClkMux
    port map (
            O => \N__4172\,
            I => \N__4142\
        );

    \I__804\ : ClkMux
    port map (
            O => \N__4171\,
            I => \N__4142\
        );

    \I__803\ : ClkMux
    port map (
            O => \N__4170\,
            I => \N__4142\
        );

    \I__802\ : ClkMux
    port map (
            O => \N__4169\,
            I => \N__4142\
        );

    \I__801\ : ClkMux
    port map (
            O => \N__4168\,
            I => \N__4142\
        );

    \I__800\ : ClkMux
    port map (
            O => \N__4167\,
            I => \N__4142\
        );

    \I__799\ : ClkMux
    port map (
            O => \N__4166\,
            I => \N__4142\
        );

    \I__798\ : ClkMux
    port map (
            O => \N__4165\,
            I => \N__4142\
        );

    \I__797\ : GlobalMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__796\ : gio2CtrlBuf
    port map (
            O => \N__4139\,
            I => \CLK6_c_g\
        );

    \I__795\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4130\
        );

    \I__794\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4130\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4130\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__792\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4118\
        );

    \I__791\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4118\
        );

    \I__790\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4118\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4118\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__4115\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__787\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4109\,
            I => \U409_TRANSFER_ACK.N_97\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__4106\,
            I => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\
        );

    \I__784\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4100\,
            I => \U409_TRANSFER_ACK.i6_mux_0\
        );

    \I__782\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4093\
        );

    \I__781\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4090\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4093\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4090\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__778\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4082\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__776\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4076\,
            I => \U409_TRANSFER_ACK.m9_bm\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__4073\,
            I => \U409_TRANSFER_ACK.m9_am_cascade_\
        );

    \I__773\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4063\
        );

    \I__772\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4054\
        );

    \I__771\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4054\
        );

    \I__770\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4054\
        );

    \I__769\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4054\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4063\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4054\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__4049\,
            I => \N__4044\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4048\,
            I => \N__4041\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__4047\,
            I => \N__4037\
        );

    \I__763\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4032\
        );

    \I__762\ : InMux
    port map (
            O => \N__4041\,
            I => \N__4032\
        );

    \I__761\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4029\
        );

    \I__760\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4026\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4032\,
            I => \N__4021\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4029\,
            I => \N__4021\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4026\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__4021\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__754\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4009\
        );

    \I__753\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4006\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4009\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4006\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__750\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3997\
        );

    \I__749\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3994\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3997\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3994\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__746\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3986\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__3983\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3976\
        );

    \I__742\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3973\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3976\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3973\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__739\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3965\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3965\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__737\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__736\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3958\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3955\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__732\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3944\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__730\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3937\
        );

    \I__729\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3934\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3934\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3929\,
            I => \U409_TRANSFER_ACK.N_97_cascade_\
        );

    \I__725\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3922\
        );

    \I__724\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3919\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3922\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3919\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__721\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3910\
        );

    \I__720\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3907\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3910\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3907\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__3902\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__716\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3895\
        );

    \I__715\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3895\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3892\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__3887\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__3884\,
            I => \N__3878\
        );

    \I__710\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3871\
        );

    \I__709\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3871\
        );

    \I__708\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3871\
        );

    \I__707\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3868\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3871\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3868\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__704\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3859\
        );

    \I__703\ : InMux
    port map (
            O => \N__3862\,
            I => \N__3856\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3859\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3856\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__699\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3844\
        );

    \I__698\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3841\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3844\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3841\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__3836\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__694\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3830\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__692\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3823\
        );

    \I__691\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3820\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3823\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3820\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__688\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3811\
        );

    \I__687\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3808\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3811\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3808\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__684\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3799\
        );

    \I__683\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3796\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3799\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3796\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__3791\,
            I => \N__3787\
        );

    \I__679\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3782\
        );

    \I__678\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3782\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3778\
        );

    \I__676\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3775\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__3778\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3775\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__673\ : InMux
    port map (
            O => \N__3770\,
            I => \N__3766\
        );

    \I__672\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3763\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3766\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3763\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__669\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3755\,
            I => \U409_TICK.TICK503_11\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__666\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3746\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__664\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3740\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__662\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__661\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3731\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__659\ : Odrv12
    port map (
            O => \N__3728\,
            I => \CIA_ENABLEm\
        );

    \I__658\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3722\,
            I => \N__3717\
        );

    \I__656\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3712\
        );

    \I__655\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3712\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3717\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3712\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__652\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3701\
        );

    \I__651\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3701\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__3698\,
            I => \N__3694\
        );

    \I__648\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3691\
        );

    \I__647\ : Sp12to4
    port map (
            O => \N__3694\,
            I => \N__3686\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3691\,
            I => \N__3686\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__3686\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \N__3679\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__3682\,
            I => \N__3676\
        );

    \I__642\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3671\
        );

    \I__641\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3671\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3671\,
            I => \N__3667\
        );

    \I__639\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3664\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3667\,
            I => \N__3659\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3664\,
            I => \N__3659\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__634\ : Span4Mux_h
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__3650\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__632\ : SRMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__3641\,
            I => \U409_TRANSFER_ACK.RESETn_c_i\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3638\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__3635\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_\
        );

    \I__627\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3624\
        );

    \I__626\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3624\
        );

    \I__625\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3619\
        );

    \I__624\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3619\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3624\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3619\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__621\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3599\
        );

    \I__620\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3599\
        );

    \I__619\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3599\
        );

    \I__618\ : InMux
    port map (
            O => \N__3611\,
            I => \N__3599\
        );

    \I__617\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3599\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3599\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__615\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3590\
        );

    \I__614\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3590\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3590\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\
        );

    \I__612\ : IoInMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__610\ : Span4Mux_s0_v
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__609\ : Sp12to4
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__608\ : Span12Mux_h
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__607\ : Span12Mux_v
    port map (
            O => \N__3572\,
            I => \N__3568\
        );

    \I__606\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3565\
        );

    \I__605\ : Odrv12
    port map (
            O => \N__3568\,
            I => \TICK60_c\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3565\,
            I => \TICK60_c\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__602\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3554\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__600\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3547\
        );

    \I__599\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3547\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3544\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__596\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3535\
        );

    \I__595\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3535\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3532\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3527\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__591\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3521\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__588\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3512\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__585\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3502\
        );

    \I__584\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3499\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3502\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3499\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__581\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3490\
        );

    \I__580\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3487\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3490\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3487\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__577\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3478\
        );

    \I__576\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3475\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3478\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3475\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__572\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3463\
        );

    \I__571\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3460\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3463\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3460\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__568\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3451\
        );

    \I__567\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3448\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3451\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3448\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__564\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3434\
        );

    \I__563\ : InMux
    port map (
            O => \N__3442\,
            I => \N__3434\
        );

    \I__562\ : InMux
    port map (
            O => \N__3441\,
            I => \N__3434\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3434\,
            I => \N__3427\
        );

    \I__560\ : InMux
    port map (
            O => \N__3433\,
            I => \N__3420\
        );

    \I__559\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3420\
        );

    \I__558\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3420\
        );

    \I__557\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3417\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__3427\,
            I => \U409_TICK.TICK603_10\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3420\,
            I => \U409_TICK.TICK603_10\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3417\,
            I => \U409_TICK.TICK603_10\
        );

    \I__553\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3395\
        );

    \I__552\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3395\
        );

    \I__551\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3395\
        );

    \I__550\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3395\
        );

    \I__549\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3392\
        );

    \I__548\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3387\
        );

    \I__547\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3387\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3395\,
            I => \U409_TICK.TICK603_14\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3392\,
            I => \U409_TICK.TICK603_14\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3387\,
            I => \U409_TICK.TICK603_14\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3380\,
            I => \N__3375\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__3379\,
            I => \N__3368\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__3378\,
            I => \N__3365\
        );

    \I__540\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3362\
        );

    \I__539\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3355\
        );

    \I__538\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3355\
        );

    \I__537\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3355\
        );

    \I__536\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3348\
        );

    \I__535\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3348\
        );

    \I__534\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3348\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3362\,
            I => \U409_TICK.TICK603_9\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3355\,
            I => \U409_TICK.TICK603_9\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3348\,
            I => \U409_TICK.TICK603_9\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3341\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3335\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__527\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3328\
        );

    \I__526\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3328\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3325\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__523\ : InMux
    port map (
            O => \N__3320\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__522\ : InMux
    port map (
            O => \N__3317\,
            I => \bfn_9_6_0_\
        );

    \I__521\ : InMux
    port map (
            O => \N__3314\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__520\ : InMux
    port map (
            O => \N__3311\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__519\ : InMux
    port map (
            O => \N__3308\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__518\ : InMux
    port map (
            O => \N__3305\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__517\ : InMux
    port map (
            O => \N__3302\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__516\ : InMux
    port map (
            O => \N__3299\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__515\ : InMux
    port map (
            O => \N__3296\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__514\ : InMux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__511\ : Sp12to4
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__510\ : Span12Mux_h
    port map (
            O => \N__3281\,
            I => \N__3278\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__3278\,
            I => \A_c_13\
        );

    \I__508\ : IoInMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__506\ : Span4Mux_s1_h
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__505\ : Sp12to4
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__504\ : Span12Mux_s9_v
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__503\ : Span12Mux_h
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__502\ : Odrv12
    port map (
            O => \N__3257\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS1_i\
        );

    \I__501\ : InMux
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__499\ : Span4Mux_v
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__498\ : Sp12to4
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__497\ : Odrv12
    port map (
            O => \N__3242\,
            I => \A_c_12\
        );

    \I__496\ : IoInMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__494\ : Span4Mux_s2_h
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__493\ : Sp12to4
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__492\ : Span12Mux_s9_v
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__491\ : Span12Mux_h
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__490\ : Odrv12
    port map (
            O => \N__3221\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS0_i\
        );

    \I__489\ : InMux
    port map (
            O => \N__3218\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__488\ : InMux
    port map (
            O => \N__3215\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__487\ : InMux
    port map (
            O => \N__3212\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__486\ : InMux
    port map (
            O => \N__3209\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__485\ : InMux
    port map (
            O => \N__3206\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__484\ : InMux
    port map (
            O => \N__3203\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__483\ : InMux
    port map (
            O => \N__3200\,
            I => \bfn_8_9_0_\
        );

    \I__482\ : InMux
    port map (
            O => \N__3197\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__481\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3191\,
            I => \N__3187\
        );

    \I__479\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3184\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__3187\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3184\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__476\ : InMux
    port map (
            O => \N__3179\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__475\ : InMux
    port map (
            O => \N__3176\,
            I => \N__3173\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3173\,
            I => \N__3169\
        );

    \I__473\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3166\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3169\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3166\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__470\ : InMux
    port map (
            O => \N__3161\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__469\ : InMux
    port map (
            O => \N__3158\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__468\ : InMux
    port map (
            O => \N__3155\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__467\ : InMux
    port map (
            O => \N__3152\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__466\ : InMux
    port map (
            O => \N__3149\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__465\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3143\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3143\,
            I => \N__3139\
        );

    \I__463\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__462\ : Span4Mux_h
    port map (
            O => \N__3139\,
            I => \N__3133\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3136\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__3133\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__459\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3121\
        );

    \I__457\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3118\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__3121\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3118\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__454\ : IoInMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3110\,
            I => \N__3107\
        );

    \I__452\ : IoSpan4Mux
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__451\ : IoSpan4Mux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__450\ : Span4Mux_s2_v
    port map (
            O => \N__3101\,
            I => \N__3098\
        );

    \I__449\ : Sp12to4
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__448\ : Span12Mux_v
    port map (
            O => \N__3095\,
            I => \N__3092\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__3092\,
            I => \nBUFEN_c\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__3089\,
            I => \N__3085\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__3088\,
            I => \N__3082\
        );

    \I__444\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3076\
        );

    \I__443\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3076\
        );

    \I__442\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3073\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3076\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3073\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__3068\,
            I => \N__3062\
        );

    \I__438\ : InMux
    port map (
            O => \N__3067\,
            I => \N__3055\
        );

    \I__437\ : InMux
    port map (
            O => \N__3066\,
            I => \N__3055\
        );

    \I__436\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3055\
        );

    \I__435\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3052\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3055\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3052\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__432\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3043\
        );

    \I__431\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3040\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3043\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3040\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__428\ : InMux
    port map (
            O => \N__3035\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__427\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3028\
        );

    \I__426\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3025\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3028\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3025\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__423\ : InMux
    port map (
            O => \N__3020\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__422\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3013\
        );

    \I__421\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3010\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3013\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3010\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__418\ : InMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3002\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__416\ : InMux
    port map (
            O => \N__2999\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__415\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2992\
        );

    \I__414\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2989\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2992\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2989\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__411\ : InMux
    port map (
            O => \N__2984\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__410\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2978\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__408\ : InMux
    port map (
            O => \N__2975\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__407\ : InMux
    port map (
            O => \N__2972\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__406\ : InMux
    port map (
            O => \N__2969\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__405\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2962\
        );

    \I__404\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2959\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2962\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2959\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__401\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2944\
        );

    \I__400\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2944\
        );

    \I__399\ : InMux
    port map (
            O => \N__2952\,
            I => \N__2941\
        );

    \I__398\ : InMux
    port map (
            O => \N__2951\,
            I => \N__2936\
        );

    \I__397\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2936\
        );

    \I__396\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2933\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2944\,
            I => \N__2928\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2928\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2936\,
            I => \N__2925\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2933\,
            I => \N__2922\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__2928\,
            I => \N__2919\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__2925\,
            I => \N__2916\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__2922\,
            I => \N__2913\
        );

    \I__388\ : Sp12to4
    port map (
            O => \N__2919\,
            I => \N__2910\
        );

    \I__387\ : Span4Mux_h
    port map (
            O => \N__2916\,
            I => \N__2907\
        );

    \I__386\ : Span4Mux_h
    port map (
            O => \N__2913\,
            I => \N__2904\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__2910\,
            I => \A_c_23\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__2907\,
            I => \A_c_23\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2904\,
            I => \A_c_23\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__380\ : IoSpan4Mux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__379\ : Span4Mux_s2_v
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__378\ : Sp12to4
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__377\ : Span12Mux_v
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__376\ : Span12Mux_h
    port map (
            O => \N__2879\,
            I => \N__2876\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__2876\,
            I => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\
        );

    \I__374\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2870\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__372\ : Odrv12
    port map (
            O => \N__2867\,
            I => \U409_ADDRESS_DECODE.un10_ROMENZ0\
        );

    \I__371\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2861\,
            I => \U409_TICK.TICK603_8\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__2858\,
            I => \U409_TICK.TICK603_11_cascade_\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__2855\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__367\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2846\
        );

    \I__366\ : InMux
    port map (
            O => \N__2851\,
            I => \N__2846\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__364\ : Span4Mux_h
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__363\ : Span4Mux_v
    port map (
            O => \N__2840\,
            I => \N__2837\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__2837\,
            I => \A_c_29\
        );

    \I__361\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2831\,
            I => \U409_CIA.g0Z0Z_2\
        );

    \I__359\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2822\
        );

    \I__358\ : InMux
    port map (
            O => \N__2827\,
            I => \N__2822\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__355\ : Sp12to4
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__2813\,
            I => \A_c_31\
        );

    \I__353\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2804\
        );

    \I__352\ : InMux
    port map (
            O => \N__2809\,
            I => \N__2804\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__350\ : Span4Mux_v
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__349\ : Sp12to4
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__348\ : Odrv12
    port map (
            O => \N__2795\,
            I => \A_c_30\
        );

    \I__347\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2789\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\
        );

    \I__345\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2780\
        );

    \I__344\ : InMux
    port map (
            O => \N__2785\,
            I => \N__2773\
        );

    \I__343\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2773\
        );

    \I__342\ : InMux
    port map (
            O => \N__2783\,
            I => \N__2773\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2780\,
            I => \N__2770\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2767\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__2770\,
            I => \N__2764\
        );

    \I__338\ : Span12Mux_v
    port map (
            O => \N__2767\,
            I => \N__2761\
        );

    \I__337\ : Sp12to4
    port map (
            O => \N__2764\,
            I => \N__2758\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__2761\,
            I => \A_c_21\
        );

    \I__335\ : Odrv12
    port map (
            O => \N__2758\,
            I => \A_c_21\
        );

    \I__334\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__2747\,
            I => \N__2742\
        );

    \I__331\ : InMux
    port map (
            O => \N__2746\,
            I => \N__2737\
        );

    \I__330\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2737\
        );

    \I__329\ : Sp12to4
    port map (
            O => \N__2742\,
            I => \N__2732\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2737\,
            I => \N__2732\
        );

    \I__327\ : Odrv12
    port map (
            O => \N__2732\,
            I => \A_c_20\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__325\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2720\
        );

    \I__324\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2720\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__322\ : Odrv4
    port map (
            O => \N__2717\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__2714\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\
        );

    \I__320\ : InMux
    port map (
            O => \N__2711\,
            I => \N__2706\
        );

    \I__319\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2701\
        );

    \I__318\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2701\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2706\,
            I => \N__2698\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2701\,
            I => \N__2695\
        );

    \I__315\ : Span4Mux_v
    port map (
            O => \N__2698\,
            I => \N__2692\
        );

    \I__314\ : Span4Mux_h
    port map (
            O => \N__2695\,
            I => \N__2689\
        );

    \I__313\ : Sp12to4
    port map (
            O => \N__2692\,
            I => \N__2686\
        );

    \I__312\ : Span4Mux_v
    port map (
            O => \N__2689\,
            I => \N__2683\
        );

    \I__311\ : Span12Mux_h
    port map (
            O => \N__2686\,
            I => \N__2680\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__2683\,
            I => \N__2677\
        );

    \I__309\ : Span12Mux_v
    port map (
            O => \N__2680\,
            I => \N__2674\
        );

    \I__308\ : Span4Mux_v
    port map (
            O => \N__2677\,
            I => \N__2671\
        );

    \I__307\ : Odrv12
    port map (
            O => \N__2674\,
            I => \A_c_19\
        );

    \I__306\ : Odrv4
    port map (
            O => \N__2671\,
            I => \A_c_19\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__2666\,
            I => \N__2661\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2665\,
            I => \N__2657\
        );

    \I__303\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2653\
        );

    \I__302\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2644\
        );

    \I__301\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2644\
        );

    \I__300\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2644\
        );

    \I__299\ : InMux
    port map (
            O => \N__2656\,
            I => \N__2644\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2653\,
            I => \N__2641\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2644\,
            I => \N__2636\
        );

    \I__296\ : Sp12to4
    port map (
            O => \N__2641\,
            I => \N__2636\
        );

    \I__295\ : Span12Mux_v
    port map (
            O => \N__2636\,
            I => \N__2633\
        );

    \I__294\ : Odrv12
    port map (
            O => \N__2633\,
            I => \A_c_22\
        );

    \I__293\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2627\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2627\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\
        );

    \I__291\ : InMux
    port map (
            O => \N__2624\,
            I => \N__2621\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2621\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__289\ : IoInMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__287\ : Span4Mux_s0_v
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__2609\,
            I => \N__2606\
        );

    \I__285\ : Span4Mux_v
    port map (
            O => \N__2606\,
            I => \N__2603\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__2603\,
            I => \N__2600\
        );

    \I__283\ : Odrv4
    port map (
            O => \N__2600\,
            I => \PORTSIZE_0_i\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__281\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2588\
        );

    \I__280\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2588\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__278\ : Span12Mux_h
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__277\ : Span12Mux_v
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__276\ : Odrv12
    port map (
            O => \N__2579\,
            I => \A_c_18\
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__2576\,
            I => \N__2572\
        );

    \I__274\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2567\
        );

    \I__273\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2567\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__271\ : Span4Mux_v
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__270\ : Span4Mux_h
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__267\ : Odrv4
    port map (
            O => \N__2552\,
            I => \A_c_16\
        );

    \I__266\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2543\
        );

    \I__265\ : InMux
    port map (
            O => \N__2548\,
            I => \N__2543\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__263\ : Span12Mux_s5_h
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__262\ : Span12Mux_v
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__261\ : Odrv12
    port map (
            O => \N__2534\,
            I => \A_c_17\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__2531\,
            I => \U409_CIA.g0Z0Z_11_cascade_\
        );

    \I__259\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__257\ : Odrv4
    port map (
            O => \N__2522\,
            I => \U409_CIA.g0Z0Z_8\
        );

    \I__256\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2516\,
            I => \N__2512\
        );

    \I__254\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2509\
        );

    \I__253\ : Span4Mux_v
    port map (
            O => \N__2512\,
            I => \N__2506\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2509\,
            I => \N__2503\
        );

    \I__251\ : Span4Mux_v
    port map (
            O => \N__2506\,
            I => \N__2498\
        );

    \I__250\ : Span4Mux_v
    port map (
            O => \N__2503\,
            I => \N__2498\
        );

    \I__249\ : Sp12to4
    port map (
            O => \N__2498\,
            I => \N__2495\
        );

    \I__248\ : Odrv12
    port map (
            O => \N__2495\,
            I => \A_c_25\
        );

    \I__247\ : CascadeMux
    port map (
            O => \N__2492\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\
        );

    \I__246\ : InMux
    port map (
            O => \N__2489\,
            I => \N__2483\
        );

    \I__245\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2483\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__243\ : Span4Mux_v
    port map (
            O => \N__2480\,
            I => \N__2477\
        );

    \I__242\ : Sp12to4
    port map (
            O => \N__2477\,
            I => \N__2474\
        );

    \I__241\ : Odrv12
    port map (
            O => \N__2474\,
            I => \A_c_27\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__239\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2462\
        );

    \I__238\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2462\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2462\,
            I => \N__2459\
        );

    \I__236\ : Span4Mux_h
    port map (
            O => \N__2459\,
            I => \N__2456\
        );

    \I__235\ : Span4Mux_v
    port map (
            O => \N__2456\,
            I => \N__2453\
        );

    \I__234\ : Odrv4
    port map (
            O => \N__2453\,
            I => \A_c_24\
        );

    \I__233\ : CascadeMux
    port map (
            O => \N__2450\,
            I => \N__2446\
        );

    \I__232\ : InMux
    port map (
            O => \N__2449\,
            I => \N__2443\
        );

    \I__231\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2440\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2443\,
            I => \N__2435\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2440\,
            I => \N__2435\
        );

    \I__228\ : Span4Mux_v
    port map (
            O => \N__2435\,
            I => \N__2432\
        );

    \I__227\ : Span4Mux_v
    port map (
            O => \N__2432\,
            I => \N__2429\
        );

    \I__226\ : Span4Mux_h
    port map (
            O => \N__2429\,
            I => \N__2426\
        );

    \I__225\ : Odrv4
    port map (
            O => \N__2426\,
            I => \A_c_26\
        );

    \I__224\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2417\
        );

    \I__223\ : InMux
    port map (
            O => \N__2422\,
            I => \N__2417\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2417\,
            I => \N__2414\
        );

    \I__221\ : Span4Mux_v
    port map (
            O => \N__2414\,
            I => \N__2411\
        );

    \I__220\ : Span4Mux_v
    port map (
            O => \N__2411\,
            I => \N__2408\
        );

    \I__219\ : Sp12to4
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__218\ : Odrv12
    port map (
            O => \N__2405\,
            I => \A_c_28\
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__2402\,
            I => \U409_CIA.g0Z0Z_10_cascade_\
        );

    \I__216\ : ClkMux
    port map (
            O => \N__2399\,
            I => \N__2369\
        );

    \I__215\ : ClkMux
    port map (
            O => \N__2398\,
            I => \N__2369\
        );

    \I__214\ : ClkMux
    port map (
            O => \N__2397\,
            I => \N__2369\
        );

    \I__213\ : ClkMux
    port map (
            O => \N__2396\,
            I => \N__2369\
        );

    \I__212\ : ClkMux
    port map (
            O => \N__2395\,
            I => \N__2369\
        );

    \I__211\ : ClkMux
    port map (
            O => \N__2394\,
            I => \N__2369\
        );

    \I__210\ : ClkMux
    port map (
            O => \N__2393\,
            I => \N__2369\
        );

    \I__209\ : ClkMux
    port map (
            O => \N__2392\,
            I => \N__2369\
        );

    \I__208\ : ClkMux
    port map (
            O => \N__2391\,
            I => \N__2369\
        );

    \I__207\ : ClkMux
    port map (
            O => \N__2390\,
            I => \N__2369\
        );

    \I__206\ : GlobalMux
    port map (
            O => \N__2369\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2390\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2397\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2393\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__2391\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__2398\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2396\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__2394\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2392\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__2399\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2395\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2709\,
            in1 => \N__2593\,
            in2 => \N__2576\,
            in3 => \N__2548\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2519\,
            in1 => \N__2710\,
            in2 => \N__2597\,
            in3 => \N__2575\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2753\,
            in1 => \N__2549\,
            in2 => \N__2531\,
            in3 => \N__2528\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5611\,
            in1 => \N__2949\,
            in2 => \_gnd_net_\,
            in3 => \N__2786\,
            lcout => \U409_CIA.g0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2467\,
            in1 => \N__2488\,
            in2 => \N__2450\,
            in3 => \N__2515\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2851\,
            in1 => \N__2422\,
            in2 => \N__2492\,
            in3 => \N__2792\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2828\,
            in1 => \N__2489\,
            in2 => \N__2471\,
            in3 => \N__2449\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2664\,
            in1 => \N__2423\,
            in2 => \N__2402\,
            in3 => \N__2834\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2852\,
            lcout => \U409_CIA.g0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2827\,
            in2 => \_gnd_net_\,
            in3 => \N__2809\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2784\,
            in1 => \N__2660\,
            in2 => \N__2729\,
            in3 => \N__2746\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un6_ROMEN_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__2951\,
            in1 => \_gnd_net_\,
            in2 => \N__2666\,
            in3 => \N__2785\,
            lcout => \U409_ADDRESS_DECODE.un6_ROMENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2745\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2656\,
            in1 => \N__2725\,
            in2 => \N__2714\,
            in3 => \N__5322\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2950\,
            in1 => \N__2711\,
            in2 => \N__2665\,
            in3 => \N__2630\,
            lcout => \U409_ADDRESS_DECODE.un10_ROMENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__2953\,
            in1 => \N__3124\,
            in2 => \N__5612\,
            in3 => \N__2624\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2965\,
            in1 => \N__2954\,
            in2 => \_gnd_net_\,
            in3 => \N__5345\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2966\,
            in1 => \N__2952\,
            in2 => \_gnd_net_\,
            in3 => \N__5326\,
            lcout => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__2873\,
            in2 => \_gnd_net_\,
            in3 => \N__4818\,
            lcout => \U409_ADDRESS_DECODE_un1_ROMEN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__2996\,
            in1 => \N__3017\,
            in2 => \_gnd_net_\,
            in3 => \N__3065\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3431\,
            in1 => \N__3404\,
            in2 => \N__3378\,
            in3 => \N__3005\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3067\,
            in1 => \_gnd_net_\,
            in2 => \N__3089\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3432\,
            in1 => \N__3405\,
            in2 => \N__3379\,
            in3 => \N__2981\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3176\,
            in1 => \N__3047\,
            in2 => \N__3088\,
            in3 => \N__3146\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2864\,
            in1 => \N__3194\,
            in2 => \N__2858\,
            in3 => \N__3032\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3066\,
            in1 => \N__3433\,
            in2 => \N__2855\,
            in3 => \N__3371\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3081\,
            in2 => \N__3068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3046\,
            in2 => \_gnd_net_\,
            in3 => \N__3035\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__4174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3031\,
            in2 => \_gnd_net_\,
            in3 => \N__3020\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__4174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3016\,
            in2 => \_gnd_net_\,
            in3 => \N__2999\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2995\,
            in2 => \_gnd_net_\,
            in3 => \N__2984\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__4174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3538\,
            in2 => \_gnd_net_\,
            in3 => \N__2975\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3466\,
            in2 => \_gnd_net_\,
            in3 => \N__2972\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__4174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3505\,
            in2 => \_gnd_net_\,
            in3 => \N__2969\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3550\,
            in2 => \_gnd_net_\,
            in3 => \N__3200\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3481\,
            in2 => \_gnd_net_\,
            in3 => \N__3197\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__4175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3190\,
            in2 => \_gnd_net_\,
            in3 => \N__3179\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__4175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3172\,
            in2 => \_gnd_net_\,
            in3 => \N__3161\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__4175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3493\,
            in2 => \_gnd_net_\,
            in3 => \N__3158\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__4175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__3155\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3454\,
            in2 => \_gnd_net_\,
            in3 => \N__3152\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3142\,
            in2 => \_gnd_net_\,
            in3 => \N__3149\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__5335\,
            in1 => \N__3128\,
            in2 => \N__4825\,
            in3 => \N__4867\,
            lcout => \nBUFEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3293\,
            in2 => \_gnd_net_\,
            in3 => \N__3737\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3254\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3781\,
            in2 => \N__3884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3802\,
            in2 => \_gnd_net_\,
            in3 => \N__3218\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__4168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3925\,
            in2 => \_gnd_net_\,
            in3 => \N__3215\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__4168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3862\,
            in2 => \_gnd_net_\,
            in3 => \N__3212\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__4168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3826\,
            in2 => \_gnd_net_\,
            in3 => \N__3209\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4012\,
            in2 => \_gnd_net_\,
            in3 => \N__3206\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3847\,
            in2 => \_gnd_net_\,
            in3 => \N__3203\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__4168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3814\,
            in2 => \_gnd_net_\,
            in3 => \N__3320\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__4168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4190\,
            in2 => \_gnd_net_\,
            in3 => \N__3317\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3898\,
            in2 => \_gnd_net_\,
            in3 => \N__3314\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3979\,
            in2 => \_gnd_net_\,
            in3 => \N__3311\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3913\,
            in2 => \_gnd_net_\,
            in3 => \N__3308\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4000\,
            in2 => \_gnd_net_\,
            in3 => \N__3305\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3961\,
            in2 => \_gnd_net_\,
            in3 => \N__3302\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3940\,
            in2 => \_gnd_net_\,
            in3 => \N__3299\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3770\,
            in2 => \_gnd_net_\,
            in3 => \N__3296\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__3430\,
            in1 => \N__3571\,
            in2 => \N__3380\,
            in3 => \N__3406\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3410\,
            in1 => \N__3443\,
            in2 => \N__3560\,
            in3 => \N__3374\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3551\,
            in1 => \N__3539\,
            in2 => \N__3509\,
            in3 => \N__3332\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3408\,
            in1 => \N__3441\,
            in2 => \N__3527\,
            in3 => \N__3524\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3409\,
            in1 => \N__3442\,
            in2 => \N__3518\,
            in3 => \N__3373\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3494\,
            in1 => \N__3482\,
            in2 => \N__3470\,
            in3 => \N__3455\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3407\,
            in1 => \N__3372\,
            in2 => \N__3341\,
            in3 => \N__3338\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__3707\,
            in1 => \N__4492\,
            in2 => \N__3683\,
            in3 => \N__3721\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__3706\,
            in1 => \N__4491\,
            in2 => \N__3682\,
            in3 => \N__3720\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__3725\,
            in1 => \N__3697\,
            in2 => \N__4496\,
            in3 => \N__3670\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__3647\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010011"
        )
    port map (
            in0 => \N__3596\,
            in1 => \N__3630\,
            in2 => \N__4969\,
            in3 => \N__3610\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__3612\,
            in1 => \N__5592\,
            in2 => \N__3638\,
            in3 => \N__4421\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3595\,
            in1 => \N__3629\,
            in2 => \N__4968\,
            in3 => \N__3611\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011001000"
        )
    port map (
            in0 => \N__3613\,
            in1 => \N__5590\,
            in2 => \N__3635\,
            in3 => \N__3631\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__3614\,
            in1 => \N__5591\,
            in2 => \_gnd_net_\,
            in3 => \N__3632\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5349\,
            in1 => \N__5266\,
            in2 => \N__5604\,
            in3 => \N__5004\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3827\,
            in1 => \N__3926\,
            in2 => \_gnd_net_\,
            in3 => \N__3881\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3758\,
            in1 => \N__3914\,
            in2 => \N__3902\,
            in3 => \N__3899\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__4306\,
            in1 => \N__4233\,
            in2 => \N__3887\,
            in3 => \N__3882\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3790\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__3863\,
            in1 => \N__3962\,
            in2 => \N__3851\,
            in3 => \N__3941\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4231\,
            in1 => \N__4270\,
            in2 => \N__3836\,
            in3 => \N__3833\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3815\,
            in1 => \N__3803\,
            in2 => \N__3791\,
            in3 => \N__3769\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4232\,
            in1 => \N__4271\,
            in2 => \N__3752\,
            in3 => \N__4307\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__4229\,
            in2 => \N__4318\,
            in3 => \N__3743\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3980\,
            in1 => \N__4189\,
            in2 => \N__4016\,
            in3 => \N__4001\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__3989\,
            in1 => \N__4272\,
            in2 => \N__3983\,
            in3 => \N__4308\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4274\,
            in1 => \N__4230\,
            in2 => \N__4319\,
            in3 => \N__3968\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4228\,
            in1 => \N__4275\,
            in2 => \N__3950\,
            in3 => \N__4315\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4642\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4127\,
            in1 => \_gnd_net_\,
            in2 => \N__5576\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4066\,
            in1 => \N__4136\,
            in2 => \N__4965\,
            in3 => \N__4126\,
            lcout => \U409_TRANSFER_ACK.N_97\,
            ltout => \U409_TRANSFER_ACK.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__4040\,
            in1 => \N__4437\,
            in2 => \N__3929\,
            in3 => \N__4457\,
            lcout => \U409_TRANSFER_ACK.m9_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4135\,
            in2 => \_gnd_net_\,
            in3 => \N__4125\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100001111"
        )
    port map (
            in0 => \N__4442\,
            in1 => \N__4458\,
            in2 => \N__4115\,
            in3 => \N__4068\,
            lcout => \U409_TRANSFER_ACK.i6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001000"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__4112\,
            in2 => \N__4048\,
            in3 => \N__4097\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5537\,
            in1 => \_gnd_net_\,
            in2 => \N__4106\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__4069\,
            in1 => \N__5536\,
            in2 => \N__4049\,
            in3 => \N__4103\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4882\,
            in2 => \_gnd_net_\,
            in3 => \N__4096\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__4438\,
            in1 => \N__4459\,
            in2 => \N__4047\,
            in3 => \N__4085\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000001010"
        )
    port map (
            in0 => \N__5542\,
            in1 => \N__4079\,
            in2 => \N__4073\,
            in3 => \N__4070\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5541\,
            in2 => \_gnd_net_\,
            in3 => \N__4460\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__4356\,
            in1 => \N__4420\,
            in2 => \N__4373\,
            in3 => \N__4409\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4403\,
            in3 => \N__5579\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011101010"
        )
    port map (
            in0 => \N__4384\,
            in1 => \N__4372\,
            in2 => \N__5600\,
            in3 => \N__4778\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4358\,
            in1 => \_gnd_net_\,
            in2 => \N__5599\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__4371\,
            in2 => \_gnd_net_\,
            in3 => \N__4357\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__4316\,
            in1 => \N__4330\,
            in2 => \N__4241\,
            in3 => \N__4276\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4317\,
            in1 => \N__4277\,
            in2 => \N__4240\,
            in3 => \N__4199\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4677\,
            in2 => \N__4721\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4559\,
            in2 => \_gnd_net_\,
            in3 => \N__4532\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__4624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4751\,
            in2 => \_gnd_net_\,
            in3 => \N__4529\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4581\,
            in2 => \_gnd_net_\,
            in3 => \N__4526\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__4624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4602\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__4753\,
            in1 => \N__4507\,
            in2 => \N__4520\,
            in3 => \N__4714\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101001100"
        )
    port map (
            in0 => \N__4715\,
            in1 => \N__4517\,
            in2 => \N__4511\,
            in3 => \N__4752\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4678\,
            in1 => \N__4582\,
            in2 => \N__4607\,
            in3 => \N__4560\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__4755\,
            in1 => \N__4717\,
            in2 => \_gnd_net_\,
            in3 => \N__4680\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__4479\,
            in1 => \N__4757\,
            in2 => \N__4499\,
            in3 => \N__4544\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4719\,
            in2 => \_gnd_net_\,
            in3 => \N__4681\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4583\,
            in1 => \N__4756\,
            in2 => \N__4606\,
            in3 => \N__4562\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4754\,
            in1 => \N__4716\,
            in2 => \_gnd_net_\,
            in3 => \N__4679\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4641\,
            in2 => \N__4730\,
            in3 => \N__4543\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__4727\,
            in1 => \N__4718\,
            in2 => \N__4685\,
            in3 => \N__4682\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4598\,
            in1 => \N__4580\,
            in2 => \_gnd_net_\,
            in3 => \N__4561\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__5149\,
            in1 => \N__5207\,
            in2 => \N__5195\,
            in3 => \N__5101\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5420\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5205\,
            in1 => \N__5100\,
            in2 => \_gnd_net_\,
            in3 => \N__5148\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5188\,
            in2 => \N__4535\,
            in3 => \N__5062\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5420\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__5078\,
            in2 => \N__5024\,
            in3 => \N__5193\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5420\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5618\,
            in1 => \N__5125\,
            in2 => \_gnd_net_\,
            in3 => \N__5192\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5420\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__4967\,
            in1 => \N__5008\,
            in2 => \N__5165\,
            in3 => \N__5037\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5206\,
            in1 => \_gnd_net_\,
            in2 => \N__5015\,
            in3 => \N__5150\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5420\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__5012\,
            in2 => \N__4966\,
            in3 => \N__5672\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5418\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4883\,
            in1 => \N__5038\,
            in2 => \_gnd_net_\,
            in3 => \N__5164\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5418\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__5641\,
            in2 => \_gnd_net_\,
            in3 => \N__5696\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5418\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__4860\,
            in1 => \N__4829\,
            in2 => \_gnd_net_\,
            in3 => \N__5351\,
            lcout => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__5577\,
            in1 => \N__4777\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__4766\,
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__5578\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5667\,
            in1 => \N__5640\,
            in2 => \N__5126\,
            in3 => \N__5694\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5669\,
            in1 => \N__5695\,
            in2 => \_gnd_net_\,
            in3 => \N__5194\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5419\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5124\,
            in1 => \N__5666\,
            in2 => \N__5063\,
            in3 => \N__5076\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5147\,
            in1 => \N__5099\,
            in2 => \N__5168\,
            in3 => \N__5707\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5146\,
            in1 => \N__5120\,
            in2 => \N__5102\,
            in3 => \N__5077\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5668\,
            in1 => \N__5060\,
            in2 => \N__5042\,
            in3 => \N__5708\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5692\,
            in2 => \_gnd_net_\,
            in3 => \N__5636\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__5693\,
            in1 => \N__5670\,
            in2 => \N__5642\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5441\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5384\,
            lcout => \N_347_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

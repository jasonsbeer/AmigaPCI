// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 25 2025 18:07:05

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    DRA,
    SIZ,
    A,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [9:0] DRA;
    input [1:0] SIZ;
    input [20:0] A;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11804;
    wire N__11803;
    wire N__11802;
    wire N__11795;
    wire N__11794;
    wire N__11793;
    wire N__11786;
    wire N__11785;
    wire N__11784;
    wire N__11777;
    wire N__11776;
    wire N__11775;
    wire N__11768;
    wire N__11767;
    wire N__11766;
    wire N__11759;
    wire N__11758;
    wire N__11757;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11741;
    wire N__11740;
    wire N__11739;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11723;
    wire N__11722;
    wire N__11721;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11687;
    wire N__11686;
    wire N__11685;
    wire N__11678;
    wire N__11677;
    wire N__11676;
    wire N__11669;
    wire N__11668;
    wire N__11667;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11642;
    wire N__11641;
    wire N__11640;
    wire N__11633;
    wire N__11632;
    wire N__11631;
    wire N__11624;
    wire N__11623;
    wire N__11622;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11606;
    wire N__11605;
    wire N__11604;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11588;
    wire N__11587;
    wire N__11586;
    wire N__11579;
    wire N__11578;
    wire N__11577;
    wire N__11570;
    wire N__11569;
    wire N__11568;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11552;
    wire N__11551;
    wire N__11550;
    wire N__11543;
    wire N__11542;
    wire N__11541;
    wire N__11534;
    wire N__11533;
    wire N__11532;
    wire N__11525;
    wire N__11524;
    wire N__11523;
    wire N__11516;
    wire N__11515;
    wire N__11514;
    wire N__11507;
    wire N__11506;
    wire N__11505;
    wire N__11498;
    wire N__11497;
    wire N__11496;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11480;
    wire N__11479;
    wire N__11478;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11453;
    wire N__11452;
    wire N__11451;
    wire N__11444;
    wire N__11443;
    wire N__11442;
    wire N__11435;
    wire N__11434;
    wire N__11433;
    wire N__11426;
    wire N__11425;
    wire N__11424;
    wire N__11417;
    wire N__11416;
    wire N__11415;
    wire N__11408;
    wire N__11407;
    wire N__11406;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11390;
    wire N__11389;
    wire N__11388;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11372;
    wire N__11371;
    wire N__11370;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11354;
    wire N__11353;
    wire N__11352;
    wire N__11345;
    wire N__11344;
    wire N__11343;
    wire N__11336;
    wire N__11335;
    wire N__11334;
    wire N__11327;
    wire N__11326;
    wire N__11325;
    wire N__11318;
    wire N__11317;
    wire N__11316;
    wire N__11309;
    wire N__11308;
    wire N__11307;
    wire N__11300;
    wire N__11299;
    wire N__11298;
    wire N__11291;
    wire N__11290;
    wire N__11289;
    wire N__11282;
    wire N__11281;
    wire N__11280;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11255;
    wire N__11254;
    wire N__11253;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11237;
    wire N__11236;
    wire N__11235;
    wire N__11228;
    wire N__11227;
    wire N__11226;
    wire N__11219;
    wire N__11218;
    wire N__11217;
    wire N__11210;
    wire N__11209;
    wire N__11208;
    wire N__11201;
    wire N__11200;
    wire N__11199;
    wire N__11192;
    wire N__11191;
    wire N__11190;
    wire N__11183;
    wire N__11182;
    wire N__11181;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11156;
    wire N__11155;
    wire N__11154;
    wire N__11147;
    wire N__11146;
    wire N__11145;
    wire N__11138;
    wire N__11137;
    wire N__11136;
    wire N__11129;
    wire N__11128;
    wire N__11127;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11102;
    wire N__11101;
    wire N__11100;
    wire N__11093;
    wire N__11092;
    wire N__11091;
    wire N__11084;
    wire N__11083;
    wire N__11082;
    wire N__11075;
    wire N__11074;
    wire N__11073;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11057;
    wire N__11056;
    wire N__11055;
    wire N__11048;
    wire N__11047;
    wire N__11046;
    wire N__11039;
    wire N__11038;
    wire N__11037;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11021;
    wire N__11020;
    wire N__11019;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10988;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10970;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10954;
    wire N__10949;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10931;
    wire N__10928;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10921;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10904;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10873;
    wire N__10866;
    wire N__10863;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10838;
    wire N__10833;
    wire N__10828;
    wire N__10827;
    wire N__10826;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10805;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10777;
    wire N__10776;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10745;
    wire N__10742;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10714;
    wire N__10713;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10657;
    wire N__10652;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10645;
    wire N__10644;
    wire N__10643;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10633;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10627;
    wire N__10626;
    wire N__10625;
    wire N__10622;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10503;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10462;
    wire N__10459;
    wire N__10458;
    wire N__10457;
    wire N__10456;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10411;
    wire N__10408;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10389;
    wire N__10388;
    wire N__10387;
    wire N__10386;
    wire N__10385;
    wire N__10384;
    wire N__10383;
    wire N__10382;
    wire N__10381;
    wire N__10380;
    wire N__10379;
    wire N__10378;
    wire N__10377;
    wire N__10376;
    wire N__10375;
    wire N__10374;
    wire N__10373;
    wire N__10372;
    wire N__10371;
    wire N__10370;
    wire N__10369;
    wire N__10368;
    wire N__10365;
    wire N__10364;
    wire N__10363;
    wire N__10362;
    wire N__10361;
    wire N__10306;
    wire N__10303;
    wire N__10302;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10290;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10279;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10220;
    wire N__10215;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10194;
    wire N__10193;
    wire N__10190;
    wire N__10189;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10034;
    wire N__10033;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10014;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10002;
    wire N__10001;
    wire N__9998;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9980;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9901;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9893;
    wire N__9890;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9872;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9836;
    wire N__9833;
    wire N__9828;
    wire N__9821;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9809;
    wire N__9808;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9774;
    wire N__9767;
    wire N__9762;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9702;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9456;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9443;
    wire N__9442;
    wire N__9441;
    wire N__9438;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9430;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9408;
    wire N__9403;
    wire N__9398;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9377;
    wire N__9374;
    wire N__9369;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9349;
    wire N__9342;
    wire N__9337;
    wire N__9332;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9310;
    wire N__9301;
    wire N__9300;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9293;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9251;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9233;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9213;
    wire N__9204;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9186;
    wire N__9183;
    wire N__9168;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9108;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9086;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9045;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9036;
    wire N__9033;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8999;
    wire N__8996;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8986;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8975;
    wire N__8968;
    wire N__8965;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8950;
    wire N__8949;
    wire N__8946;
    wire N__8937;
    wire N__8936;
    wire N__8933;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8914;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8893;
    wire N__8892;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8875;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8809;
    wire N__8806;
    wire N__8805;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8785;
    wire N__8780;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8619;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8611;
    wire N__8608;
    wire N__8607;
    wire N__8606;
    wire N__8601;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8575;
    wire N__8566;
    wire N__8565;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8515;
    wire N__8506;
    wire N__8505;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8497;
    wire N__8494;
    wire N__8493;
    wire N__8492;
    wire N__8491;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8460;
    wire N__8455;
    wire N__8454;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8386;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8374;
    wire N__8371;
    wire N__8370;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8298;
    wire N__8295;
    wire N__8290;
    wire N__8287;
    wire N__8286;
    wire N__8285;
    wire N__8282;
    wire N__8277;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8128;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8103;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8082;
    wire N__8079;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8064;
    wire N__8061;
    wire N__8056;
    wire N__8053;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7986;
    wire N__7985;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7964;
    wire N__7961;
    wire N__7960;
    wire N__7957;
    wire N__7950;
    wire N__7945;
    wire N__7942;
    wire N__7937;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7871;
    wire N__7866;
    wire N__7861;
    wire N__7858;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7840;
    wire N__7835;
    wire N__7832;
    wire N__7831;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7800;
    wire N__7795;
    wire N__7794;
    wire N__7793;
    wire N__7792;
    wire N__7791;
    wire N__7790;
    wire N__7787;
    wire N__7780;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7742;
    wire N__7739;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7715;
    wire N__7712;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7688;
    wire N__7683;
    wire N__7680;
    wire N__7673;
    wire N__7670;
    wire N__7665;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7595;
    wire N__7594;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7491;
    wire N__7490;
    wire N__7487;
    wire N__7482;
    wire N__7477;
    wire N__7474;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7468;
    wire N__7467;
    wire N__7466;
    wire N__7463;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7448;
    wire N__7445;
    wire N__7440;
    wire N__7429;
    wire N__7428;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7405;
    wire N__7402;
    wire N__7401;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7378;
    wire N__7377;
    wire N__7376;
    wire N__7373;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7355;
    wire N__7352;
    wire N__7339;
    wire N__7336;
    wire N__7335;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7277;
    wire N__7272;
    wire N__7269;
    wire N__7258;
    wire N__7255;
    wire N__7254;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7237;
    wire N__7234;
    wire N__7225;
    wire N__7224;
    wire N__7223;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7180;
    wire N__7177;
    wire N__7176;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7098;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7086;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7050;
    wire N__7047;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7006;
    wire N__7005;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__6997;
    wire N__6992;
    wire N__6989;
    wire N__6988;
    wire N__6987;
    wire N__6982;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6971;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6951;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6900;
    wire N__6899;
    wire N__6894;
    wire N__6891;
    wire N__6886;
    wire N__6883;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6862;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6847;
    wire N__6844;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6838;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6816;
    wire N__6815;
    wire N__6814;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6798;
    wire N__6791;
    wire N__6788;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6762;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6736;
    wire N__6735;
    wire N__6734;
    wire N__6731;
    wire N__6730;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6658;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6594;
    wire N__6589;
    wire N__6588;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6552;
    wire N__6549;
    wire N__6548;
    wire N__6545;
    wire N__6544;
    wire N__6543;
    wire N__6542;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6525;
    wire N__6522;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6468;
    wire N__6465;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6426;
    wire N__6425;
    wire N__6424;
    wire N__6423;
    wire N__6422;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6316;
    wire N__6313;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6294;
    wire N__6287;
    wire N__6286;
    wire N__6285;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6274;
    wire N__6271;
    wire N__6270;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6232;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6217;
    wire N__6216;
    wire N__6215;
    wire N__6214;
    wire N__6211;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6181;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6160;
    wire N__6155;
    wire N__6148;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6105;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6067;
    wire N__6064;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6052;
    wire N__6049;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6009;
    wire N__6008;
    wire N__6005;
    wire N__6000;
    wire N__5995;
    wire N__5992;
    wire N__5991;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5963;
    wire N__5958;
    wire N__5953;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5832;
    wire N__5829;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5794;
    wire N__5793;
    wire N__5788;
    wire N__5783;
    wire N__5780;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5719;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5707;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5691;
    wire N__5688;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5661;
    wire N__5656;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5629;
    wire N__5626;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5618;
    wire N__5615;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5596;
    wire N__5593;
    wire N__5588;
    wire N__5585;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5506;
    wire N__5505;
    wire N__5502;
    wire N__5501;
    wire N__5500;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5488;
    wire N__5487;
    wire N__5484;
    wire N__5483;
    wire N__5480;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5455;
    wire N__5454;
    wire N__5453;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5441;
    wire N__5440;
    wire N__5435;
    wire N__5430;
    wire N__5423;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5401;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5381;
    wire N__5378;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5355;
    wire N__5350;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5274;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5225;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5200;
    wire N__5197;
    wire N__5196;
    wire N__5195;
    wire N__5192;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5170;
    wire N__5169;
    wire N__5168;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5143;
    wire N__5142;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5116;
    wire N__5115;
    wire N__5110;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5098;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5092;
    wire N__5091;
    wire N__5090;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5035;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5014;
    wire N__5011;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4741;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4621;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4557;
    wire N__4556;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4533;
    wire N__4526;
    wire N__4519;
    wire N__4516;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4489;
    wire N__4488;
    wire N__4487;
    wire N__4486;
    wire N__4481;
    wire N__4476;
    wire N__4471;
    wire N__4470;
    wire N__4467;
    wire N__4466;
    wire N__4465;
    wire N__4460;
    wire N__4455;
    wire N__4450;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4382;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4271;
    wire N__4268;
    wire N__4263;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire A_c_14;
    wire A_c_7;
    wire A_c_16;
    wire A_c_18;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.N_350_cascade_ ;
    wire \U712_CHIP_RAM.N_376_cascade_ ;
    wire \U712_CHIP_RAM.N_280_cascade_ ;
    wire \U712_CHIP_RAM.N_288_cascade_ ;
    wire \U712_CHIP_RAM.N_325_cascade_ ;
    wire \U712_CHIP_RAM.N_308_cascade_ ;
    wire \U712_CHIP_RAM.N_350_0_cascade_ ;
    wire \U712_CHIP_RAM.N_355_cascade_ ;
    wire \U712_CHIP_RAM.N_389_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ;
    wire \U712_CHIP_RAM.N_348_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0 ;
    wire CLK_EN_c;
    wire DBRn_c_i_cascade_;
    wire DBRn_c_i_0;
    wire LATCH_CLK_0_i;
    wire CLK40_PLL_iso_i;
    wire VBENn_c;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_350 ;
    wire \U712_CHIP_RAM.N_283 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0 ;
    wire \U712_CHIP_RAM.N_403 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ;
    wire \U712_CHIP_RAM.N_280 ;
    wire \U712_CHIP_RAM.N_301_cascade_ ;
    wire \U712_CHIP_RAM.N_280_2 ;
    wire \U712_CHIP_RAM.N_192 ;
    wire \U712_CHIP_RAM.N_192_cascade_ ;
    wire \U712_CHIP_RAM.N_215 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_ ;
    wire \U712_CHIP_RAM.N_345 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0 ;
    wire bfn_8_9_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_100 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_400_cascade_ ;
    wire \U712_CHIP_RAM.N_266 ;
    wire \U712_CHIP_RAM.N_304_cascade_ ;
    wire \U712_CHIP_RAM.N_249 ;
    wire \U712_CHIP_RAM.N_355 ;
    wire \U712_CHIP_RAM.N_350_0 ;
    wire \U712_CHIP_RAM.N_291_cascade_ ;
    wire RAMSPACEn_c;
    wire N_246;
    wire REGENn_c;
    wire LATCH_REG;
    wire REG_CPU_CYCLE;
    wire \INVU712_REG_SM.REGENnC_net ;
    wire ASn_c;
    wire C3_c;
    wire \INVU712_REG_SM.ASnC_net ;
    wire A_c_9;
    wire A_c_2;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire A_c_3;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ;
    wire \U712_CHIP_RAM.N_399 ;
    wire \U712_CHIP_RAM.N_399_cascade_ ;
    wire \U712_CHIP_RAM.N_277 ;
    wire \U712_CHIP_RAM.N_277_cascade_ ;
    wire \U712_CHIP_RAM.N_347_cascade_ ;
    wire \U712_CHIP_RAM.N_353 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_347 ;
    wire \U712_CHIP_RAM.N_343_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_391 ;
    wire \U712_CHIP_RAM.N_391_cascade_ ;
    wire \U712_CHIP_RAM.N_387 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ;
    wire \U712_CHIP_RAM.N_352 ;
    wire \U712_CHIP_RAM.N_343 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire AWEn_c;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0 ;
    wire \U712_CHIP_RAM.N_234 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0 ;
    wire WRITE_CYCLE;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ;
    wire \U712_CHIP_RAM.N_292 ;
    wire \U712_CHIP_RAM.N_19 ;
    wire \U712_BYTE_ENABLE.N_185_i ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_5 ;
    wire \INVU712_REG_SM.CYCLE_RUNC_net ;
    wire \U712_REG_SM.N_229_cascade_ ;
    wire \INVU712_REG_SM.STATE_COUNTER_0C_net ;
    wire \U712_REG_SM.LATCH_REG_0_sqmuxa ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_4 ;
    wire \U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_ ;
    wire \U712_REG_SM.REG_CPU_CYCLE_e_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_224 ;
    wire \U712_REG_SM.N_224_cascade_ ;
    wire \U712_REG_SM.N_209_cascade_ ;
    wire \U712_REG_SM.LDSn_7_iv_i_0 ;
    wire \U712_REG_SM.N_297_cascade_ ;
    wire LDSn_c;
    wire \U712_REG_SM.N_295_cascade_ ;
    wire \U712_REG_SM.N_153 ;
    wire UDSn_c;
    wire \INVU712_REG_SM.C3_SYNC_1C_net ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.CYCLE_RUNZ0 ;
    wire TSn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \INVU712_REG_SM.C1_SYNC_0C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ;
    wire \U712_CHIP_RAM.N_136 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_10_8_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire BANK0_c;
    wire A_c_20;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_405 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_405_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_303_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ;
    wire \U712_CHIP_RAM.N_348 ;
    wire \U712_CHIP_RAM.N_186 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.N_198 ;
    wire \U712_CHIP_RAM.N_389 ;
    wire \U712_CHIP_RAM.N_313_cascade_ ;
    wire \U712_CHIP_RAM.N_314 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire LATCH_RAM;
    wire DBR_SYNCZ0Z_1;
    wire DBR_SYNCZ0Z_0;
    wire \U712_BYTE_ENABLE.N_319_cascade_ ;
    wire N_58_i;
    wire \U712_BYTE_ENABLE.N_320 ;
    wire N_56_i;
    wire \U712_BYTE_ENABLE.N_318 ;
    wire \U712_BYTE_ENABLE.N_323_cascade_ ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ;
    wire N_54_i;
    wire DBENn_c;
    wire DMA_CYCLE;
    wire \U712_BYTE_ENABLE.N_315_cascade_ ;
    wire N_60_i;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_3 ;
    wire REG_WRITE_CYCLE;
    wire RnW_c;
    wire \U712_REG_SM.UDSn_7_iv_i_0 ;
    wire \U712_REG_SM.N_245 ;
    wire \U712_REG_SM.un15_0_i_0_0_0 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_6 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_7 ;
    wire \U712_REG_SM.N_209 ;
    wire \U712_REG_SM.N_229 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_1 ;
    wire \INVU712_REG_SM.REG_TACKC_net ;
    wire N_858_i;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_2 ;
    wire \U712_REG_SM.REG_TACK_0_sqmuxa ;
    wire DBRn_c;
    wire \U712_REG_SM.DBR_SYNCZ0Z_0 ;
    wire \U712_REG_SM.DBR_SYNCZ0Z_1 ;
    wire \INVU712_REG_SM.DBR_SYNC_0C_net ;
    wire REG_CYCLE;
    wire DRDENn_c;
    wire N_118_i;
    wire A_c_0;
    wire U712_BYTE_ENABLE_UUBE_i;
    wire LLBEn_c;
    wire N_386;
    wire SIZ_c_0;
    wire A_c_1;
    wire SIZ_c_1;
    wire UMBEn_c;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire CLK40_PLL;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ;
    wire TACK_EN_i_ess;
    wire RASn_c;
    wire WEn_c;
    wire CRCSn_c;
    wire CMA_c_10;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire A_c_6;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire CLK40_PLL_g;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.N_8 ;
    wire RESETn_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire CPU_TACK;
    wire \U712_CYCLE_TERM.N_227_i_0_0_cascade_ ;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.N_227_i_0_en_cascade_ ;
    wire RESETn_c_i;
    wire \U712_CYCLE_TERM.N_227_i_0_en_0 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire CPU_CYCLE;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire CASUn_c;
    wire CASLn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_9;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_3;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_0;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire AGNUS_REV_c;
    wire DRA_c_6;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4051),
            .RESETB(N__8704),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11804),
            .DIN(N__11803),
            .DOUT(N__11802),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11804),
            .PADOUT(N__11803),
            .PADIN(N__11802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7054),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11795),
            .DIN(N__11794),
            .DOUT(N__11793),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11795),
            .PADOUT(N__11794),
            .PADIN(N__11793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11786),
            .DIN(N__11785),
            .DOUT(N__11784),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11786),
            .PADOUT(N__11785),
            .PADIN(N__11784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9604),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11777),
            .DIN(N__11776),
            .DOUT(N__11775),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11777),
            .PADOUT(N__11776),
            .PADIN(N__11775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4801),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11768),
            .DIN(N__11767),
            .DOUT(N__11766),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11768),
            .PADOUT(N__11767),
            .PADIN(N__11766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11759),
            .DIN(N__11758),
            .DOUT(N__11757),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11759),
            .PADOUT(N__11758),
            .PADIN(N__11757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11750),
            .DIN(N__11749),
            .DOUT(N__11748),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11750),
            .PADOUT(N__11749),
            .PADIN(N__11748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11741),
            .DIN(N__11740),
            .DOUT(N__11739),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11741),
            .PADOUT(N__11740),
            .PADIN(N__11739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11732),
            .DIN(N__11731),
            .DOUT(N__11730),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11732),
            .PADOUT(N__11731),
            .PADIN(N__11730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11723),
            .DIN(N__11722),
            .DOUT(N__11721),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11723),
            .PADOUT(N__11722),
            .PADIN(N__11721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11714),
            .DIN(N__11713),
            .DOUT(N__11712),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11714),
            .PADOUT(N__11713),
            .PADIN(N__11712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11705),
            .DIN(N__11704),
            .DOUT(N__11703),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11705),
            .PADOUT(N__11704),
            .PADIN(N__11703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11696),
            .DIN(N__11695),
            .DOUT(N__11694),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11696),
            .PADOUT(N__11695),
            .PADIN(N__11694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11687),
            .DIN(N__11686),
            .DOUT(N__11685),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11687),
            .PADOUT(N__11686),
            .PADIN(N__11685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11678),
            .DIN(N__11677),
            .DOUT(N__11676),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11678),
            .PADOUT(N__11677),
            .PADIN(N__11676),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11669),
            .DIN(N__11668),
            .DOUT(N__11667),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11669),
            .PADOUT(N__11668),
            .PADIN(N__11667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4345),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11660),
            .DIN(N__11659),
            .DOUT(N__11658),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11660),
            .PADOUT(N__11659),
            .PADIN(N__11658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11651),
            .DIN(N__11650),
            .DOUT(N__11649),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11651),
            .PADOUT(N__11650),
            .PADIN(N__11649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11642),
            .DIN(N__11641),
            .DOUT(N__11640),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11642),
            .PADOUT(N__11641),
            .PADIN(N__11640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11633),
            .DIN(N__11632),
            .DOUT(N__11631),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11633),
            .PADOUT(N__11632),
            .PADIN(N__11631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11624),
            .DIN(N__11623),
            .DOUT(N__11622),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11624),
            .PADOUT(N__11623),
            .PADIN(N__11622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8743),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11615),
            .DIN(N__11614),
            .DOUT(N__11613),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11615),
            .PADOUT(N__11614),
            .PADIN(N__11613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11606),
            .DIN(N__11605),
            .DOUT(N__11604),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11606),
            .PADOUT(N__11605),
            .PADIN(N__11604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7903),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11597),
            .DIN(N__11596),
            .DOUT(N__11595),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11597),
            .PADOUT(N__11596),
            .PADIN(N__11595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11588),
            .DIN(N__11587),
            .DOUT(N__11586),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11588),
            .PADOUT(N__11587),
            .PADIN(N__11586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11579),
            .DIN(N__11578),
            .DOUT(N__11577),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11579),
            .PADOUT(N__11578),
            .PADIN(N__11577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11570),
            .DIN(N__11569),
            .DOUT(N__11568),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11570),
            .PADOUT(N__11569),
            .PADIN(N__11568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11561),
            .DIN(N__11560),
            .DOUT(N__11559),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11561),
            .PADOUT(N__11560),
            .PADIN(N__11559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11552),
            .DIN(N__11551),
            .DOUT(N__11550),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11552),
            .PADOUT(N__11551),
            .PADIN(N__11550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4800),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11543),
            .DIN(N__11542),
            .DOUT(N__11541),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11543),
            .PADOUT(N__11542),
            .PADIN(N__11541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11534),
            .DIN(N__11533),
            .DOUT(N__11532),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11534),
            .PADOUT(N__11533),
            .PADIN(N__11532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11525),
            .DIN(N__11524),
            .DOUT(N__11523),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11525),
            .PADOUT(N__11524),
            .PADIN(N__11523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11516),
            .DIN(N__11515),
            .DOUT(N__11514),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11516),
            .PADOUT(N__11515),
            .PADIN(N__11514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11507),
            .DIN(N__11506),
            .DOUT(N__11505),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11507),
            .PADOUT(N__11506),
            .PADIN(N__11505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11498),
            .DIN(N__11497),
            .DOUT(N__11496),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11498),
            .PADOUT(N__11497),
            .PADIN(N__11496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8332),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11489),
            .DIN(N__11488),
            .DOUT(N__11487),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11489),
            .PADOUT(N__11488),
            .PADIN(N__11487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11480),
            .DIN(N__11479),
            .DOUT(N__11478),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11480),
            .PADOUT(N__11479),
            .PADIN(N__11478),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4389),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11471),
            .DIN(N__11470),
            .DOUT(N__11469),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11471),
            .PADOUT(N__11470),
            .PADIN(N__11469),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4183),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11462),
            .DIN(N__11461),
            .DOUT(N__11460),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11462),
            .PADOUT(N__11461),
            .PADIN(N__11460),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11453),
            .DIN(N__11452),
            .DOUT(N__11451),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11453),
            .PADOUT(N__11452),
            .PADIN(N__11451),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4711),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11444),
            .DIN(N__11443),
            .DOUT(N__11442),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11444),
            .PADOUT(N__11443),
            .PADIN(N__11442),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11435),
            .DIN(N__11434),
            .DOUT(N__11433),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11435),
            .PADOUT(N__11434),
            .PADIN(N__11433),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11426),
            .DIN(N__11425),
            .DOUT(N__11424),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11426),
            .PADOUT(N__11425),
            .PADIN(N__11424),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11417),
            .DIN(N__11416),
            .DOUT(N__11415),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11417),
            .PADOUT(N__11416),
            .PADIN(N__11415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11408),
            .DIN(N__11407),
            .DOUT(N__11406),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11408),
            .PADOUT(N__11407),
            .PADIN(N__11406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11399),
            .DIN(N__11398),
            .DOUT(N__11397),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11399),
            .PADOUT(N__11398),
            .PADIN(N__11397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8725),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11390),
            .DIN(N__11389),
            .DOUT(N__11388),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11390),
            .PADOUT(N__11389),
            .PADIN(N__11388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11381),
            .DIN(N__11380),
            .DOUT(N__11379),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11381),
            .PADOUT(N__11380),
            .PADIN(N__11379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4382),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11372),
            .DIN(N__11371),
            .DOUT(N__11370),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11372),
            .PADOUT(N__11371),
            .PADIN(N__11370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9538),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11363),
            .DIN(N__11362),
            .DOUT(N__11361),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11363),
            .PADOUT(N__11362),
            .PADIN(N__11361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11354),
            .DIN(N__11353),
            .DOUT(N__11352),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11354),
            .PADOUT(N__11353),
            .PADIN(N__11352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7078),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11345),
            .DIN(N__11344),
            .DOUT(N__11343),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11345),
            .PADOUT(N__11344),
            .PADIN(N__11343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8254),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11336),
            .DIN(N__11335),
            .DOUT(N__11334),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11336),
            .PADOUT(N__11335),
            .PADIN(N__11334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4765),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11327),
            .DIN(N__11326),
            .DOUT(N__11325),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11327),
            .PADOUT(N__11326),
            .PADIN(N__11325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11318),
            .DIN(N__11317),
            .DOUT(N__11316),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11318),
            .PADOUT(N__11317),
            .PADIN(N__11316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11309),
            .DIN(N__11308),
            .DOUT(N__11307),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11309),
            .PADOUT(N__11308),
            .PADIN(N__11307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7123),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11300),
            .DIN(N__11299),
            .DOUT(N__11298),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11300),
            .PADOUT(N__11299),
            .PADIN(N__11298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8314),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11291),
            .DIN(N__11290),
            .DOUT(N__11289),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11291),
            .PADOUT(N__11290),
            .PADIN(N__11289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11282),
            .DIN(N__11281),
            .DOUT(N__11280),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11282),
            .PADOUT(N__11281),
            .PADIN(N__11280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11273),
            .DIN(N__11272),
            .DOUT(N__11271),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11273),
            .PADOUT(N__11272),
            .PADIN(N__11271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11264),
            .DIN(N__11263),
            .DOUT(N__11262),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11264),
            .PADOUT(N__11263),
            .PADIN(N__11262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11255),
            .DIN(N__11254),
            .DOUT(N__11253),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11255),
            .PADOUT(N__11254),
            .PADIN(N__11253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11246),
            .DIN(N__11245),
            .DOUT(N__11244),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11246),
            .PADOUT(N__11245),
            .PADIN(N__11244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11237),
            .DIN(N__11236),
            .DOUT(N__11235),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11237),
            .PADOUT(N__11236),
            .PADIN(N__11235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8179),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11228),
            .DIN(N__11227),
            .DOUT(N__11226),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11228),
            .PADOUT(N__11227),
            .PADIN(N__11226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8005),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11219),
            .DIN(N__11218),
            .DOUT(N__11217),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11219),
            .PADOUT(N__11218),
            .PADIN(N__11217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11210),
            .DIN(N__11209),
            .DOUT(N__11208),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11210),
            .PADOUT(N__11209),
            .PADIN(N__11208),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6937),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11201),
            .DIN(N__11200),
            .DOUT(N__11199),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11201),
            .PADOUT(N__11200),
            .PADIN(N__11199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7318),
            .DIN0(),
            .DOUT0(N__8413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11192),
            .DIN(N__11191),
            .DOUT(N__11190),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11192),
            .PADOUT(N__11191),
            .PADIN(N__11190),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9475),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11183),
            .DIN(N__11182),
            .DOUT(N__11181),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11183),
            .PADOUT(N__11182),
            .PADIN(N__11181),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11174),
            .DIN(N__11173),
            .DOUT(N__11172),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11174),
            .PADOUT(N__11173),
            .PADIN(N__11172),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11165),
            .DIN(N__11164),
            .DOUT(N__11163),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11165),
            .PADOUT(N__11164),
            .PADIN(N__11163),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11156),
            .DIN(N__11155),
            .DOUT(N__11154),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11156),
            .PADOUT(N__11155),
            .PADIN(N__11154),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11147),
            .DIN(N__11146),
            .DOUT(N__11145),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11147),
            .PADOUT(N__11146),
            .PADIN(N__11145),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11138),
            .DIN(N__11137),
            .DOUT(N__11136),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11138),
            .PADOUT(N__11137),
            .PADIN(N__11136),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11129),
            .DIN(N__11128),
            .DOUT(N__11127),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11129),
            .PADOUT(N__11128),
            .PADIN(N__11127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11120),
            .DIN(N__11119),
            .DOUT(N__11118),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11120),
            .PADOUT(N__11119),
            .PADIN(N__11118),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11111),
            .DIN(N__11110),
            .DOUT(N__11109),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11111),
            .PADOUT(N__11110),
            .PADIN(N__11109),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5983),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11102),
            .DIN(N__11101),
            .DOUT(N__11100),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11102),
            .PADOUT(N__11101),
            .PADIN(N__11100),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11093),
            .DIN(N__11092),
            .DOUT(N__11091),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11093),
            .PADOUT(N__11092),
            .PADIN(N__11091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11084),
            .DIN(N__11083),
            .DOUT(N__11082),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11084),
            .PADOUT(N__11083),
            .PADIN(N__11082),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11075),
            .DIN(N__11074),
            .DOUT(N__11073),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11075),
            .PADOUT(N__11074),
            .PADIN(N__11073),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11066),
            .DIN(N__11065),
            .DOUT(N__11064),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11066),
            .PADOUT(N__11065),
            .PADIN(N__11064),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9565),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11057),
            .DIN(N__11056),
            .DOUT(N__11055),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11057),
            .PADOUT(N__11056),
            .PADIN(N__11055),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11048),
            .DIN(N__11047),
            .DOUT(N__11046),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11048),
            .PADOUT(N__11047),
            .PADIN(N__11046),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11039),
            .DIN(N__11038),
            .DOUT(N__11037),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11039),
            .PADOUT(N__11038),
            .PADIN(N__11037),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4408),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11030),
            .DIN(N__11029),
            .DOUT(N__11028),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11030),
            .PADOUT(N__11029),
            .PADIN(N__11028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11021),
            .DIN(N__11020),
            .DOUT(N__11019),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11021),
            .PADOUT(N__11020),
            .PADIN(N__11019),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4390),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11012),
            .DIN(N__11011),
            .DOUT(N__11010),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11012),
            .PADOUT(N__11011),
            .PADIN(N__11010),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__2674 (
            .O(N__10993),
            .I(N__10989));
    InMux I__2673 (
            .O(N__10992),
            .I(N__10977));
    InMux I__2672 (
            .O(N__10989),
            .I(N__10974));
    InMux I__2671 (
            .O(N__10988),
            .I(N__10971));
    InMux I__2670 (
            .O(N__10987),
            .I(N__10961));
    InMux I__2669 (
            .O(N__10986),
            .I(N__10961));
    InMux I__2668 (
            .O(N__10985),
            .I(N__10961));
    InMux I__2667 (
            .O(N__10984),
            .I(N__10961));
    InMux I__2666 (
            .O(N__10983),
            .I(N__10958));
    InMux I__2665 (
            .O(N__10982),
            .I(N__10955));
    InMux I__2664 (
            .O(N__10981),
            .I(N__10949));
    InMux I__2663 (
            .O(N__10980),
            .I(N__10949));
    LocalMux I__2662 (
            .O(N__10977),
            .I(N__10942));
    LocalMux I__2661 (
            .O(N__10974),
            .I(N__10942));
    LocalMux I__2660 (
            .O(N__10971),
            .I(N__10942));
    InMux I__2659 (
            .O(N__10970),
            .I(N__10939));
    LocalMux I__2658 (
            .O(N__10961),
            .I(N__10936));
    LocalMux I__2657 (
            .O(N__10958),
            .I(N__10931));
    LocalMux I__2656 (
            .O(N__10955),
            .I(N__10931));
    InMux I__2655 (
            .O(N__10954),
            .I(N__10928));
    LocalMux I__2654 (
            .O(N__10949),
            .I(N__10917));
    Span4Mux_v I__2653 (
            .O(N__10942),
            .I(N__10914));
    LocalMux I__2652 (
            .O(N__10939),
            .I(N__10911));
    Span4Mux_v I__2651 (
            .O(N__10936),
            .I(N__10904));
    Span4Mux_h I__2650 (
            .O(N__10931),
            .I(N__10904));
    LocalMux I__2649 (
            .O(N__10928),
            .I(N__10904));
    InMux I__2648 (
            .O(N__10927),
            .I(N__10897));
    InMux I__2647 (
            .O(N__10926),
            .I(N__10897));
    InMux I__2646 (
            .O(N__10925),
            .I(N__10897));
    InMux I__2645 (
            .O(N__10924),
            .I(N__10894));
    InMux I__2644 (
            .O(N__10923),
            .I(N__10891));
    InMux I__2643 (
            .O(N__10922),
            .I(N__10884));
    InMux I__2642 (
            .O(N__10921),
            .I(N__10884));
    InMux I__2641 (
            .O(N__10920),
            .I(N__10884));
    Span4Mux_v I__2640 (
            .O(N__10917),
            .I(N__10881));
    Span4Mux_h I__2639 (
            .O(N__10914),
            .I(N__10878));
    Span4Mux_v I__2638 (
            .O(N__10911),
            .I(N__10873));
    Span4Mux_v I__2637 (
            .O(N__10904),
            .I(N__10873));
    LocalMux I__2636 (
            .O(N__10897),
            .I(N__10866));
    LocalMux I__2635 (
            .O(N__10894),
            .I(N__10866));
    LocalMux I__2634 (
            .O(N__10891),
            .I(N__10866));
    LocalMux I__2633 (
            .O(N__10884),
            .I(N__10863));
    Sp12to4 I__2632 (
            .O(N__10881),
            .I(N__10858));
    Sp12to4 I__2631 (
            .O(N__10878),
            .I(N__10858));
    Sp12to4 I__2630 (
            .O(N__10873),
            .I(N__10855));
    Span12Mux_h I__2629 (
            .O(N__10866),
            .I(N__10852));
    Span12Mux_v I__2628 (
            .O(N__10863),
            .I(N__10849));
    Span12Mux_h I__2627 (
            .O(N__10858),
            .I(N__10846));
    Span12Mux_v I__2626 (
            .O(N__10855),
            .I(N__10843));
    Span12Mux_v I__2625 (
            .O(N__10852),
            .I(N__10838));
    Span12Mux_h I__2624 (
            .O(N__10849),
            .I(N__10838));
    Span12Mux_v I__2623 (
            .O(N__10846),
            .I(N__10833));
    Span12Mux_h I__2622 (
            .O(N__10843),
            .I(N__10833));
    Odrv12 I__2621 (
            .O(N__10838),
            .I(AGNUS_REV_c));
    Odrv12 I__2620 (
            .O(N__10833),
            .I(AGNUS_REV_c));
    InMux I__2619 (
            .O(N__10828),
            .I(N__10823));
    InMux I__2618 (
            .O(N__10827),
            .I(N__10819));
    InMux I__2617 (
            .O(N__10826),
            .I(N__10816));
    LocalMux I__2616 (
            .O(N__10823),
            .I(N__10813));
    InMux I__2615 (
            .O(N__10822),
            .I(N__10810));
    LocalMux I__2614 (
            .O(N__10819),
            .I(N__10805));
    LocalMux I__2613 (
            .O(N__10816),
            .I(N__10805));
    Span4Mux_h I__2612 (
            .O(N__10813),
            .I(N__10800));
    LocalMux I__2611 (
            .O(N__10810),
            .I(N__10800));
    Span4Mux_h I__2610 (
            .O(N__10805),
            .I(N__10797));
    Span4Mux_v I__2609 (
            .O(N__10800),
            .I(N__10794));
    Sp12to4 I__2608 (
            .O(N__10797),
            .I(N__10791));
    Sp12to4 I__2607 (
            .O(N__10794),
            .I(N__10788));
    Span12Mux_v I__2606 (
            .O(N__10791),
            .I(N__10785));
    Span12Mux_h I__2605 (
            .O(N__10788),
            .I(N__10782));
    Odrv12 I__2604 (
            .O(N__10785),
            .I(DRA_c_6));
    Odrv12 I__2603 (
            .O(N__10782),
            .I(DRA_c_6));
    InMux I__2602 (
            .O(N__10777),
            .I(N__10772));
    InMux I__2601 (
            .O(N__10776),
            .I(N__10769));
    InMux I__2600 (
            .O(N__10775),
            .I(N__10766));
    LocalMux I__2599 (
            .O(N__10772),
            .I(N__10762));
    LocalMux I__2598 (
            .O(N__10769),
            .I(N__10759));
    LocalMux I__2597 (
            .O(N__10766),
            .I(N__10756));
    CascadeMux I__2596 (
            .O(N__10765),
            .I(N__10753));
    Span4Mux_v I__2595 (
            .O(N__10762),
            .I(N__10750));
    Span4Mux_v I__2594 (
            .O(N__10759),
            .I(N__10745));
    Span4Mux_v I__2593 (
            .O(N__10756),
            .I(N__10745));
    InMux I__2592 (
            .O(N__10753),
            .I(N__10742));
    Sp12to4 I__2591 (
            .O(N__10750),
            .I(N__10735));
    Sp12to4 I__2590 (
            .O(N__10745),
            .I(N__10735));
    LocalMux I__2589 (
            .O(N__10742),
            .I(N__10735));
    Span12Mux_h I__2588 (
            .O(N__10735),
            .I(N__10732));
    Odrv12 I__2587 (
            .O(N__10732),
            .I(DRA_c_7));
    InMux I__2586 (
            .O(N__10729),
            .I(N__10726));
    LocalMux I__2585 (
            .O(N__10726),
            .I(N__10723));
    Span4Mux_v I__2584 (
            .O(N__10723),
            .I(N__10720));
    Odrv4 I__2583 (
            .O(N__10720),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    ClkMux I__2582 (
            .O(N__10717),
            .I(N__10702));
    ClkMux I__2581 (
            .O(N__10716),
            .I(N__10702));
    ClkMux I__2580 (
            .O(N__10715),
            .I(N__10702));
    ClkMux I__2579 (
            .O(N__10714),
            .I(N__10702));
    ClkMux I__2578 (
            .O(N__10713),
            .I(N__10702));
    GlobalMux I__2577 (
            .O(N__10702),
            .I(N__10699));
    gio2CtrlBuf I__2576 (
            .O(N__10699),
            .I(C3_c_g));
    CEMux I__2575 (
            .O(N__10696),
            .I(N__10669));
    CEMux I__2574 (
            .O(N__10695),
            .I(N__10669));
    CEMux I__2573 (
            .O(N__10694),
            .I(N__10669));
    CEMux I__2572 (
            .O(N__10693),
            .I(N__10669));
    CEMux I__2571 (
            .O(N__10692),
            .I(N__10669));
    CEMux I__2570 (
            .O(N__10691),
            .I(N__10669));
    CEMux I__2569 (
            .O(N__10690),
            .I(N__10669));
    CEMux I__2568 (
            .O(N__10689),
            .I(N__10669));
    CEMux I__2567 (
            .O(N__10688),
            .I(N__10669));
    GlobalMux I__2566 (
            .O(N__10669),
            .I(N__10666));
    gio2CtrlBuf I__2565 (
            .O(N__10666),
            .I(DBRn_c_i_0_g));
    InMux I__2564 (
            .O(N__10663),
            .I(N__10657));
    InMux I__2563 (
            .O(N__10662),
            .I(N__10652));
    InMux I__2562 (
            .O(N__10661),
            .I(N__10652));
    InMux I__2561 (
            .O(N__10660),
            .I(N__10649));
    LocalMux I__2560 (
            .O(N__10657),
            .I(N__10636));
    LocalMux I__2559 (
            .O(N__10652),
            .I(N__10629));
    LocalMux I__2558 (
            .O(N__10649),
            .I(N__10622));
    SRMux I__2557 (
            .O(N__10648),
            .I(N__10516));
    SRMux I__2556 (
            .O(N__10647),
            .I(N__10516));
    SRMux I__2555 (
            .O(N__10646),
            .I(N__10516));
    SRMux I__2554 (
            .O(N__10645),
            .I(N__10516));
    SRMux I__2553 (
            .O(N__10644),
            .I(N__10516));
    SRMux I__2552 (
            .O(N__10643),
            .I(N__10516));
    SRMux I__2551 (
            .O(N__10642),
            .I(N__10516));
    SRMux I__2550 (
            .O(N__10641),
            .I(N__10516));
    SRMux I__2549 (
            .O(N__10640),
            .I(N__10516));
    SRMux I__2548 (
            .O(N__10639),
            .I(N__10516));
    Glb2LocalMux I__2547 (
            .O(N__10636),
            .I(N__10516));
    SRMux I__2546 (
            .O(N__10635),
            .I(N__10516));
    SRMux I__2545 (
            .O(N__10634),
            .I(N__10516));
    SRMux I__2544 (
            .O(N__10633),
            .I(N__10516));
    SRMux I__2543 (
            .O(N__10632),
            .I(N__10516));
    Glb2LocalMux I__2542 (
            .O(N__10629),
            .I(N__10516));
    SRMux I__2541 (
            .O(N__10628),
            .I(N__10516));
    SRMux I__2540 (
            .O(N__10627),
            .I(N__10516));
    SRMux I__2539 (
            .O(N__10626),
            .I(N__10516));
    SRMux I__2538 (
            .O(N__10625),
            .I(N__10516));
    Glb2LocalMux I__2537 (
            .O(N__10622),
            .I(N__10516));
    SRMux I__2536 (
            .O(N__10621),
            .I(N__10516));
    SRMux I__2535 (
            .O(N__10620),
            .I(N__10516));
    SRMux I__2534 (
            .O(N__10619),
            .I(N__10516));
    SRMux I__2533 (
            .O(N__10618),
            .I(N__10516));
    SRMux I__2532 (
            .O(N__10617),
            .I(N__10516));
    SRMux I__2531 (
            .O(N__10616),
            .I(N__10516));
    SRMux I__2530 (
            .O(N__10615),
            .I(N__10516));
    SRMux I__2529 (
            .O(N__10614),
            .I(N__10516));
    SRMux I__2528 (
            .O(N__10613),
            .I(N__10516));
    SRMux I__2527 (
            .O(N__10612),
            .I(N__10516));
    SRMux I__2526 (
            .O(N__10611),
            .I(N__10516));
    SRMux I__2525 (
            .O(N__10610),
            .I(N__10516));
    SRMux I__2524 (
            .O(N__10609),
            .I(N__10516));
    SRMux I__2523 (
            .O(N__10608),
            .I(N__10516));
    SRMux I__2522 (
            .O(N__10607),
            .I(N__10516));
    SRMux I__2521 (
            .O(N__10606),
            .I(N__10516));
    SRMux I__2520 (
            .O(N__10605),
            .I(N__10516));
    SRMux I__2519 (
            .O(N__10604),
            .I(N__10516));
    SRMux I__2518 (
            .O(N__10603),
            .I(N__10516));
    SRMux I__2517 (
            .O(N__10602),
            .I(N__10516));
    SRMux I__2516 (
            .O(N__10601),
            .I(N__10516));
    GlobalMux I__2515 (
            .O(N__10516),
            .I(N__10513));
    gio2CtrlBuf I__2514 (
            .O(N__10513),
            .I(RESETn_c_i_g));
    InMux I__2513 (
            .O(N__10510),
            .I(N__10503));
    InMux I__2512 (
            .O(N__10509),
            .I(N__10503));
    InMux I__2511 (
            .O(N__10508),
            .I(N__10499));
    LocalMux I__2510 (
            .O(N__10503),
            .I(N__10496));
    InMux I__2509 (
            .O(N__10502),
            .I(N__10493));
    LocalMux I__2508 (
            .O(N__10499),
            .I(N__10490));
    Span4Mux_v I__2507 (
            .O(N__10496),
            .I(N__10485));
    LocalMux I__2506 (
            .O(N__10493),
            .I(N__10485));
    Span4Mux_v I__2505 (
            .O(N__10490),
            .I(N__10482));
    Span4Mux_v I__2504 (
            .O(N__10485),
            .I(N__10479));
    Sp12to4 I__2503 (
            .O(N__10482),
            .I(N__10476));
    Span4Mux_v I__2502 (
            .O(N__10479),
            .I(N__10473));
    Span12Mux_h I__2501 (
            .O(N__10476),
            .I(N__10470));
    Sp12to4 I__2500 (
            .O(N__10473),
            .I(N__10467));
    Span12Mux_v I__2499 (
            .O(N__10470),
            .I(N__10462));
    Span12Mux_h I__2498 (
            .O(N__10467),
            .I(N__10462));
    Odrv12 I__2497 (
            .O(N__10462),
            .I(CASUn_c));
    InMux I__2496 (
            .O(N__10459),
            .I(N__10451));
    InMux I__2495 (
            .O(N__10458),
            .I(N__10451));
    InMux I__2494 (
            .O(N__10457),
            .I(N__10448));
    InMux I__2493 (
            .O(N__10456),
            .I(N__10445));
    LocalMux I__2492 (
            .O(N__10451),
            .I(N__10442));
    LocalMux I__2491 (
            .O(N__10448),
            .I(N__10439));
    LocalMux I__2490 (
            .O(N__10445),
            .I(N__10436));
    Span4Mux_h I__2489 (
            .O(N__10442),
            .I(N__10431));
    Span4Mux_v I__2488 (
            .O(N__10439),
            .I(N__10431));
    Span4Mux_v I__2487 (
            .O(N__10436),
            .I(N__10428));
    Sp12to4 I__2486 (
            .O(N__10431),
            .I(N__10425));
    Span4Mux_v I__2485 (
            .O(N__10428),
            .I(N__10422));
    Span12Mux_h I__2484 (
            .O(N__10425),
            .I(N__10419));
    Sp12to4 I__2483 (
            .O(N__10422),
            .I(N__10416));
    Span12Mux_v I__2482 (
            .O(N__10419),
            .I(N__10411));
    Span12Mux_h I__2481 (
            .O(N__10416),
            .I(N__10411));
    Odrv12 I__2480 (
            .O(N__10411),
            .I(CASLn_c));
    InMux I__2479 (
            .O(N__10408),
            .I(N__10404));
    InMux I__2478 (
            .O(N__10407),
            .I(N__10401));
    LocalMux I__2477 (
            .O(N__10404),
            .I(N__10396));
    LocalMux I__2476 (
            .O(N__10401),
            .I(N__10396));
    Odrv12 I__2475 (
            .O(N__10396),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__2474 (
            .O(N__10393),
            .I(N__10390));
    LocalMux I__2473 (
            .O(N__10390),
            .I(N__10365));
    ClkMux I__2472 (
            .O(N__10389),
            .I(N__10306));
    ClkMux I__2471 (
            .O(N__10388),
            .I(N__10306));
    ClkMux I__2470 (
            .O(N__10387),
            .I(N__10306));
    ClkMux I__2469 (
            .O(N__10386),
            .I(N__10306));
    ClkMux I__2468 (
            .O(N__10385),
            .I(N__10306));
    ClkMux I__2467 (
            .O(N__10384),
            .I(N__10306));
    ClkMux I__2466 (
            .O(N__10383),
            .I(N__10306));
    ClkMux I__2465 (
            .O(N__10382),
            .I(N__10306));
    ClkMux I__2464 (
            .O(N__10381),
            .I(N__10306));
    ClkMux I__2463 (
            .O(N__10380),
            .I(N__10306));
    ClkMux I__2462 (
            .O(N__10379),
            .I(N__10306));
    ClkMux I__2461 (
            .O(N__10378),
            .I(N__10306));
    ClkMux I__2460 (
            .O(N__10377),
            .I(N__10306));
    ClkMux I__2459 (
            .O(N__10376),
            .I(N__10306));
    ClkMux I__2458 (
            .O(N__10375),
            .I(N__10306));
    ClkMux I__2457 (
            .O(N__10374),
            .I(N__10306));
    ClkMux I__2456 (
            .O(N__10373),
            .I(N__10306));
    ClkMux I__2455 (
            .O(N__10372),
            .I(N__10306));
    ClkMux I__2454 (
            .O(N__10371),
            .I(N__10306));
    ClkMux I__2453 (
            .O(N__10370),
            .I(N__10306));
    ClkMux I__2452 (
            .O(N__10369),
            .I(N__10306));
    ClkMux I__2451 (
            .O(N__10368),
            .I(N__10306));
    Glb2LocalMux I__2450 (
            .O(N__10365),
            .I(N__10306));
    ClkMux I__2449 (
            .O(N__10364),
            .I(N__10306));
    ClkMux I__2448 (
            .O(N__10363),
            .I(N__10306));
    ClkMux I__2447 (
            .O(N__10362),
            .I(N__10306));
    ClkMux I__2446 (
            .O(N__10361),
            .I(N__10306));
    GlobalMux I__2445 (
            .O(N__10306),
            .I(CLK80_PLL));
    InMux I__2444 (
            .O(N__10303),
            .I(N__10297));
    InMux I__2443 (
            .O(N__10302),
            .I(N__10297));
    LocalMux I__2442 (
            .O(N__10297),
            .I(N__10294));
    Odrv12 I__2441 (
            .O(N__10294),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2440 (
            .O(N__10291),
            .I(N__10286));
    InMux I__2439 (
            .O(N__10290),
            .I(N__10283));
    InMux I__2438 (
            .O(N__10289),
            .I(N__10280));
    LocalMux I__2437 (
            .O(N__10286),
            .I(N__10272));
    LocalMux I__2436 (
            .O(N__10283),
            .I(N__10272));
    LocalMux I__2435 (
            .O(N__10280),
            .I(N__10272));
    InMux I__2434 (
            .O(N__10279),
            .I(N__10269));
    Span4Mux_v I__2433 (
            .O(N__10272),
            .I(N__10266));
    LocalMux I__2432 (
            .O(N__10269),
            .I(N__10263));
    Sp12to4 I__2431 (
            .O(N__10266),
            .I(N__10260));
    Span12Mux_v I__2430 (
            .O(N__10263),
            .I(N__10257));
    Span12Mux_h I__2429 (
            .O(N__10260),
            .I(N__10254));
    Span12Mux_h I__2428 (
            .O(N__10257),
            .I(N__10249));
    Span12Mux_v I__2427 (
            .O(N__10254),
            .I(N__10249));
    Odrv12 I__2426 (
            .O(N__10249),
            .I(DRA_c_2));
    CascadeMux I__2425 (
            .O(N__10246),
            .I(N__10243));
    InMux I__2424 (
            .O(N__10243),
            .I(N__10240));
    LocalMux I__2423 (
            .O(N__10240),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2422 (
            .O(N__10237),
            .I(N__10234));
    LocalMux I__2421 (
            .O(N__10234),
            .I(N__10228));
    InMux I__2420 (
            .O(N__10233),
            .I(N__10225));
    InMux I__2419 (
            .O(N__10232),
            .I(N__10220));
    InMux I__2418 (
            .O(N__10231),
            .I(N__10220));
    Span4Mux_h I__2417 (
            .O(N__10228),
            .I(N__10215));
    LocalMux I__2416 (
            .O(N__10225),
            .I(N__10215));
    LocalMux I__2415 (
            .O(N__10220),
            .I(N__10210));
    Sp12to4 I__2414 (
            .O(N__10215),
            .I(N__10210));
    Span12Mux_v I__2413 (
            .O(N__10210),
            .I(N__10207));
    Span12Mux_h I__2412 (
            .O(N__10207),
            .I(N__10204));
    Odrv12 I__2411 (
            .O(N__10204),
            .I(DRA_c_5));
    InMux I__2410 (
            .O(N__10201),
            .I(N__10198));
    LocalMux I__2409 (
            .O(N__10198),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2408 (
            .O(N__10195),
            .I(N__10190));
    InMux I__2407 (
            .O(N__10194),
            .I(N__10184));
    InMux I__2406 (
            .O(N__10193),
            .I(N__10184));
    LocalMux I__2405 (
            .O(N__10190),
            .I(N__10181));
    InMux I__2404 (
            .O(N__10189),
            .I(N__10178));
    LocalMux I__2403 (
            .O(N__10184),
            .I(N__10175));
    Span4Mux_v I__2402 (
            .O(N__10181),
            .I(N__10172));
    LocalMux I__2401 (
            .O(N__10178),
            .I(N__10169));
    Span4Mux_v I__2400 (
            .O(N__10175),
            .I(N__10166));
    Sp12to4 I__2399 (
            .O(N__10172),
            .I(N__10163));
    Span12Mux_v I__2398 (
            .O(N__10169),
            .I(N__10158));
    Sp12to4 I__2397 (
            .O(N__10166),
            .I(N__10158));
    Span12Mux_h I__2396 (
            .O(N__10163),
            .I(N__10155));
    Span12Mux_h I__2395 (
            .O(N__10158),
            .I(N__10152));
    Odrv12 I__2394 (
            .O(N__10155),
            .I(DRA_c_8));
    Odrv12 I__2393 (
            .O(N__10152),
            .I(DRA_c_8));
    InMux I__2392 (
            .O(N__10147),
            .I(N__10144));
    LocalMux I__2391 (
            .O(N__10144),
            .I(N__10141));
    Odrv4 I__2390 (
            .O(N__10141),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    CascadeMux I__2389 (
            .O(N__10138),
            .I(N__10133));
    InMux I__2388 (
            .O(N__10137),
            .I(N__10130));
    InMux I__2387 (
            .O(N__10136),
            .I(N__10127));
    InMux I__2386 (
            .O(N__10133),
            .I(N__10124));
    LocalMux I__2385 (
            .O(N__10130),
            .I(N__10121));
    LocalMux I__2384 (
            .O(N__10127),
            .I(N__10117));
    LocalMux I__2383 (
            .O(N__10124),
            .I(N__10114));
    Span4Mux_h I__2382 (
            .O(N__10121),
            .I(N__10111));
    InMux I__2381 (
            .O(N__10120),
            .I(N__10108));
    Span4Mux_v I__2380 (
            .O(N__10117),
            .I(N__10103));
    Span4Mux_h I__2379 (
            .O(N__10114),
            .I(N__10103));
    Span4Mux_v I__2378 (
            .O(N__10111),
            .I(N__10100));
    LocalMux I__2377 (
            .O(N__10108),
            .I(N__10097));
    Sp12to4 I__2376 (
            .O(N__10103),
            .I(N__10094));
    Sp12to4 I__2375 (
            .O(N__10100),
            .I(N__10089));
    Span12Mux_v I__2374 (
            .O(N__10097),
            .I(N__10089));
    Span12Mux_v I__2373 (
            .O(N__10094),
            .I(N__10086));
    Span12Mux_h I__2372 (
            .O(N__10089),
            .I(N__10083));
    Span12Mux_h I__2371 (
            .O(N__10086),
            .I(N__10078));
    Span12Mux_v I__2370 (
            .O(N__10083),
            .I(N__10078));
    Odrv12 I__2369 (
            .O(N__10078),
            .I(DRA_c_9));
    InMux I__2368 (
            .O(N__10075),
            .I(N__10072));
    LocalMux I__2367 (
            .O(N__10072),
            .I(N__10069));
    Span12Mux_h I__2366 (
            .O(N__10069),
            .I(N__10066));
    Odrv12 I__2365 (
            .O(N__10066),
            .I(RAS0n_c));
    CascadeMux I__2364 (
            .O(N__10063),
            .I(N__10060));
    InMux I__2363 (
            .O(N__10060),
            .I(N__10057));
    LocalMux I__2362 (
            .O(N__10057),
            .I(N__10054));
    Span4Mux_v I__2361 (
            .O(N__10054),
            .I(N__10051));
    Odrv4 I__2360 (
            .O(N__10051),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2359 (
            .O(N__10048),
            .I(N__10044));
    InMux I__2358 (
            .O(N__10047),
            .I(N__10041));
    LocalMux I__2357 (
            .O(N__10044),
            .I(N__10038));
    LocalMux I__2356 (
            .O(N__10041),
            .I(N__10035));
    Span4Mux_v I__2355 (
            .O(N__10038),
            .I(N__10028));
    Span4Mux_v I__2354 (
            .O(N__10035),
            .I(N__10028));
    InMux I__2353 (
            .O(N__10034),
            .I(N__10025));
    InMux I__2352 (
            .O(N__10033),
            .I(N__10022));
    Span4Mux_v I__2351 (
            .O(N__10028),
            .I(N__10019));
    LocalMux I__2350 (
            .O(N__10025),
            .I(N__10014));
    LocalMux I__2349 (
            .O(N__10022),
            .I(N__10014));
    Sp12to4 I__2348 (
            .O(N__10019),
            .I(N__10009));
    Span12Mux_v I__2347 (
            .O(N__10014),
            .I(N__10009));
    Span12Mux_h I__2346 (
            .O(N__10009),
            .I(N__10006));
    Odrv12 I__2345 (
            .O(N__10006),
            .I(DRA_c_3));
    InMux I__2344 (
            .O(N__10003),
            .I(N__9998));
    InMux I__2343 (
            .O(N__10002),
            .I(N__9994));
    InMux I__2342 (
            .O(N__10001),
            .I(N__9991));
    LocalMux I__2341 (
            .O(N__9998),
            .I(N__9988));
    InMux I__2340 (
            .O(N__9997),
            .I(N__9985));
    LocalMux I__2339 (
            .O(N__9994),
            .I(N__9980));
    LocalMux I__2338 (
            .O(N__9991),
            .I(N__9980));
    Span4Mux_h I__2337 (
            .O(N__9988),
            .I(N__9975));
    LocalMux I__2336 (
            .O(N__9985),
            .I(N__9975));
    Span4Mux_v I__2335 (
            .O(N__9980),
            .I(N__9972));
    Span4Mux_v I__2334 (
            .O(N__9975),
            .I(N__9969));
    Span4Mux_v I__2333 (
            .O(N__9972),
            .I(N__9966));
    Span4Mux_v I__2332 (
            .O(N__9969),
            .I(N__9963));
    Sp12to4 I__2331 (
            .O(N__9966),
            .I(N__9960));
    Sp12to4 I__2330 (
            .O(N__9963),
            .I(N__9957));
    Span12Mux_h I__2329 (
            .O(N__9960),
            .I(N__9954));
    Span12Mux_h I__2328 (
            .O(N__9957),
            .I(N__9951));
    Odrv12 I__2327 (
            .O(N__9954),
            .I(DRA_c_4));
    Odrv12 I__2326 (
            .O(N__9951),
            .I(DRA_c_4));
    CascadeMux I__2325 (
            .O(N__9946),
            .I(N__9943));
    InMux I__2324 (
            .O(N__9943),
            .I(N__9940));
    LocalMux I__2323 (
            .O(N__9940),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2322 (
            .O(N__9937),
            .I(N__9934));
    LocalMux I__2321 (
            .O(N__9934),
            .I(N__9931));
    Span4Mux_v I__2320 (
            .O(N__9931),
            .I(N__9927));
    InMux I__2319 (
            .O(N__9930),
            .I(N__9924));
    Sp12to4 I__2318 (
            .O(N__9927),
            .I(N__9921));
    LocalMux I__2317 (
            .O(N__9924),
            .I(N__9918));
    Span12Mux_h I__2316 (
            .O(N__9921),
            .I(N__9915));
    Span12Mux_h I__2315 (
            .O(N__9918),
            .I(N__9912));
    Span12Mux_v I__2314 (
            .O(N__9915),
            .I(N__9909));
    Span12Mux_v I__2313 (
            .O(N__9912),
            .I(N__9906));
    Odrv12 I__2312 (
            .O(N__9909),
            .I(DRA_c_0));
    Odrv12 I__2311 (
            .O(N__9906),
            .I(DRA_c_0));
    InMux I__2310 (
            .O(N__9901),
            .I(N__9897));
    InMux I__2309 (
            .O(N__9900),
            .I(N__9894));
    LocalMux I__2308 (
            .O(N__9897),
            .I(N__9890));
    LocalMux I__2307 (
            .O(N__9894),
            .I(N__9886));
    InMux I__2306 (
            .O(N__9893),
            .I(N__9883));
    Span4Mux_v I__2305 (
            .O(N__9890),
            .I(N__9880));
    InMux I__2304 (
            .O(N__9889),
            .I(N__9877));
    Span4Mux_v I__2303 (
            .O(N__9886),
            .I(N__9872));
    LocalMux I__2302 (
            .O(N__9883),
            .I(N__9872));
    Sp12to4 I__2301 (
            .O(N__9880),
            .I(N__9867));
    LocalMux I__2300 (
            .O(N__9877),
            .I(N__9867));
    Sp12to4 I__2299 (
            .O(N__9872),
            .I(N__9864));
    Span12Mux_h I__2298 (
            .O(N__9867),
            .I(N__9861));
    Span12Mux_v I__2297 (
            .O(N__9864),
            .I(N__9858));
    Span12Mux_v I__2296 (
            .O(N__9861),
            .I(N__9855));
    Span12Mux_h I__2295 (
            .O(N__9858),
            .I(N__9852));
    Odrv12 I__2294 (
            .O(N__9855),
            .I(DRA_c_1));
    Odrv12 I__2293 (
            .O(N__9852),
            .I(DRA_c_1));
    InMux I__2292 (
            .O(N__9847),
            .I(N__9844));
    LocalMux I__2291 (
            .O(N__9844),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    CascadeMux I__2290 (
            .O(N__9841),
            .I(N__9833));
    InMux I__2289 (
            .O(N__9840),
            .I(N__9828));
    InMux I__2288 (
            .O(N__9839),
            .I(N__9828));
    InMux I__2287 (
            .O(N__9838),
            .I(N__9821));
    InMux I__2286 (
            .O(N__9837),
            .I(N__9821));
    InMux I__2285 (
            .O(N__9836),
            .I(N__9821));
    InMux I__2284 (
            .O(N__9833),
            .I(N__9818));
    LocalMux I__2283 (
            .O(N__9828),
            .I(N__9809));
    LocalMux I__2282 (
            .O(N__9821),
            .I(N__9809));
    LocalMux I__2281 (
            .O(N__9818),
            .I(N__9809));
    InMux I__2280 (
            .O(N__9817),
            .I(N__9803));
    InMux I__2279 (
            .O(N__9816),
            .I(N__9803));
    Span4Mux_v I__2278 (
            .O(N__9809),
            .I(N__9800));
    InMux I__2277 (
            .O(N__9808),
            .I(N__9797));
    LocalMux I__2276 (
            .O(N__9803),
            .I(N__9794));
    Odrv4 I__2275 (
            .O(N__9800),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2274 (
            .O(N__9797),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2273 (
            .O(N__9794),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__2272 (
            .O(N__9787),
            .I(N__9784));
    LocalMux I__2271 (
            .O(N__9784),
            .I(N__9781));
    Odrv12 I__2270 (
            .O(N__9781),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__2269 (
            .O(N__9778),
            .I(N__9767));
    InMux I__2268 (
            .O(N__9777),
            .I(N__9767));
    InMux I__2267 (
            .O(N__9776),
            .I(N__9767));
    InMux I__2266 (
            .O(N__9775),
            .I(N__9762));
    InMux I__2265 (
            .O(N__9774),
            .I(N__9762));
    LocalMux I__2264 (
            .O(N__9767),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2263 (
            .O(N__9762),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    IoInMux I__2262 (
            .O(N__9757),
            .I(N__9754));
    LocalMux I__2261 (
            .O(N__9754),
            .I(N__9751));
    Span4Mux_s2_h I__2260 (
            .O(N__9751),
            .I(N__9748));
    Sp12to4 I__2259 (
            .O(N__9748),
            .I(N__9745));
    Span12Mux_v I__2258 (
            .O(N__9745),
            .I(N__9742));
    Span12Mux_h I__2257 (
            .O(N__9742),
            .I(N__9739));
    Odrv12 I__2256 (
            .O(N__9739),
            .I(CMA_c_3));
    CEMux I__2255 (
            .O(N__9736),
            .I(N__9732));
    CEMux I__2254 (
            .O(N__9735),
            .I(N__9729));
    LocalMux I__2253 (
            .O(N__9732),
            .I(N__9722));
    LocalMux I__2252 (
            .O(N__9729),
            .I(N__9719));
    CEMux I__2251 (
            .O(N__9728),
            .I(N__9716));
    CEMux I__2250 (
            .O(N__9727),
            .I(N__9713));
    CEMux I__2249 (
            .O(N__9726),
            .I(N__9710));
    CEMux I__2248 (
            .O(N__9725),
            .I(N__9707));
    Span4Mux_h I__2247 (
            .O(N__9722),
            .I(N__9702));
    Span4Mux_h I__2246 (
            .O(N__9719),
            .I(N__9702));
    LocalMux I__2245 (
            .O(N__9716),
            .I(N__9697));
    LocalMux I__2244 (
            .O(N__9713),
            .I(N__9697));
    LocalMux I__2243 (
            .O(N__9710),
            .I(N__9694));
    LocalMux I__2242 (
            .O(N__9707),
            .I(N__9691));
    Odrv4 I__2241 (
            .O(N__9702),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2240 (
            .O(N__9697),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2239 (
            .O(N__9694),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2238 (
            .O(N__9691),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2237 (
            .O(N__9682),
            .I(N__9679));
    LocalMux I__2236 (
            .O(N__9679),
            .I(N__9676));
    Span4Mux_h I__2235 (
            .O(N__9676),
            .I(N__9673));
    Odrv4 I__2234 (
            .O(N__9673),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__2233 (
            .O(N__9670),
            .I(N__9667));
    InMux I__2232 (
            .O(N__9667),
            .I(N__9664));
    LocalMux I__2231 (
            .O(N__9664),
            .I(N__9661));
    Odrv4 I__2230 (
            .O(N__9661),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2229 (
            .O(N__9658),
            .I(N__9655));
    LocalMux I__2228 (
            .O(N__9655),
            .I(N__9652));
    Span4Mux_v I__2227 (
            .O(N__9652),
            .I(N__9649));
    Odrv4 I__2226 (
            .O(N__9649),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2225 (
            .O(N__9646),
            .I(N__9643));
    LocalMux I__2224 (
            .O(N__9643),
            .I(N__9640));
    Odrv4 I__2223 (
            .O(N__9640),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2222 (
            .O(N__9637),
            .I(N__9634));
    LocalMux I__2221 (
            .O(N__9634),
            .I(N__9631));
    Odrv4 I__2220 (
            .O(N__9631),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2219 (
            .O(N__9628),
            .I(N__9625));
    LocalMux I__2218 (
            .O(N__9625),
            .I(N__9622));
    Span4Mux_h I__2217 (
            .O(N__9622),
            .I(N__9619));
    Odrv4 I__2216 (
            .O(N__9619),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2215 (
            .O(N__9616),
            .I(N__9613));
    LocalMux I__2214 (
            .O(N__9613),
            .I(N__9610));
    Span4Mux_h I__2213 (
            .O(N__9610),
            .I(N__9607));
    Odrv4 I__2212 (
            .O(N__9607),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    IoInMux I__2211 (
            .O(N__9604),
            .I(N__9601));
    LocalMux I__2210 (
            .O(N__9601),
            .I(N__9598));
    Span4Mux_s2_v I__2209 (
            .O(N__9598),
            .I(N__9595));
    Span4Mux_v I__2208 (
            .O(N__9595),
            .I(N__9592));
    Sp12to4 I__2207 (
            .O(N__9592),
            .I(N__9589));
    Span12Mux_h I__2206 (
            .O(N__9589),
            .I(N__9586));
    Odrv12 I__2205 (
            .O(N__9586),
            .I(CASn_c));
    CascadeMux I__2204 (
            .O(N__9583),
            .I(N__9580));
    InMux I__2203 (
            .O(N__9580),
            .I(N__9577));
    LocalMux I__2202 (
            .O(N__9577),
            .I(N__9574));
    Span4Mux_h I__2201 (
            .O(N__9574),
            .I(N__9571));
    Odrv4 I__2200 (
            .O(N__9571),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    CascadeMux I__2199 (
            .O(N__9568),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ));
    IoInMux I__2198 (
            .O(N__9565),
            .I(N__9562));
    LocalMux I__2197 (
            .O(N__9562),
            .I(N__9559));
    Span4Mux_s3_h I__2196 (
            .O(N__9559),
            .I(N__9556));
    Sp12to4 I__2195 (
            .O(N__9556),
            .I(N__9553));
    Span12Mux_s10_v I__2194 (
            .O(N__9553),
            .I(N__9550));
    Span12Mux_h I__2193 (
            .O(N__9550),
            .I(N__9547));
    Odrv12 I__2192 (
            .O(N__9547),
            .I(CMA_c_6));
    InMux I__2191 (
            .O(N__9544),
            .I(N__9541));
    LocalMux I__2190 (
            .O(N__9541),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__2189 (
            .O(N__9538),
            .I(N__9535));
    LocalMux I__2188 (
            .O(N__9535),
            .I(N__9532));
    IoSpan4Mux I__2187 (
            .O(N__9532),
            .I(N__9529));
    Span4Mux_s2_h I__2186 (
            .O(N__9529),
            .I(N__9526));
    Sp12to4 I__2185 (
            .O(N__9526),
            .I(N__9523));
    Span12Mux_h I__2184 (
            .O(N__9523),
            .I(N__9520));
    Odrv12 I__2183 (
            .O(N__9520),
            .I(CMA_c_4));
    InMux I__2182 (
            .O(N__9517),
            .I(N__9514));
    LocalMux I__2181 (
            .O(N__9514),
            .I(N__9511));
    Span4Mux_h I__2180 (
            .O(N__9511),
            .I(N__9508));
    Odrv4 I__2179 (
            .O(N__9508),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__2178 (
            .O(N__9505),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ));
    IoInMux I__2177 (
            .O(N__9502),
            .I(N__9499));
    LocalMux I__2176 (
            .O(N__9499),
            .I(N__9496));
    IoSpan4Mux I__2175 (
            .O(N__9496),
            .I(N__9493));
    Span4Mux_s2_h I__2174 (
            .O(N__9493),
            .I(N__9490));
    Sp12to4 I__2173 (
            .O(N__9490),
            .I(N__9487));
    Span12Mux_h I__2172 (
            .O(N__9487),
            .I(N__9484));
    Odrv12 I__2171 (
            .O(N__9484),
            .I(CMA_c_7));
    InMux I__2170 (
            .O(N__9481),
            .I(N__9478));
    LocalMux I__2169 (
            .O(N__9478),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__2168 (
            .O(N__9475),
            .I(N__9472));
    LocalMux I__2167 (
            .O(N__9472),
            .I(N__9469));
    IoSpan4Mux I__2166 (
            .O(N__9469),
            .I(N__9466));
    Span4Mux_s2_v I__2165 (
            .O(N__9466),
            .I(N__9463));
    Sp12to4 I__2164 (
            .O(N__9463),
            .I(N__9460));
    Odrv12 I__2163 (
            .O(N__9460),
            .I(CMA_c_2));
    InMux I__2162 (
            .O(N__9457),
            .I(N__9443));
    InMux I__2161 (
            .O(N__9456),
            .I(N__9443));
    CascadeMux I__2160 (
            .O(N__9455),
            .I(N__9438));
    CascadeMux I__2159 (
            .O(N__9454),
            .I(N__9434));
    CascadeMux I__2158 (
            .O(N__9453),
            .I(N__9431));
    InMux I__2157 (
            .O(N__9452),
            .I(N__9425));
    InMux I__2156 (
            .O(N__9451),
            .I(N__9425));
    InMux I__2155 (
            .O(N__9450),
            .I(N__9420));
    InMux I__2154 (
            .O(N__9449),
            .I(N__9417));
    InMux I__2153 (
            .O(N__9448),
            .I(N__9414));
    LocalMux I__2152 (
            .O(N__9443),
            .I(N__9408));
    InMux I__2151 (
            .O(N__9442),
            .I(N__9403));
    InMux I__2150 (
            .O(N__9441),
            .I(N__9403));
    InMux I__2149 (
            .O(N__9438),
            .I(N__9398));
    InMux I__2148 (
            .O(N__9437),
            .I(N__9398));
    InMux I__2147 (
            .O(N__9434),
            .I(N__9393));
    InMux I__2146 (
            .O(N__9431),
            .I(N__9393));
    InMux I__2145 (
            .O(N__9430),
            .I(N__9390));
    LocalMux I__2144 (
            .O(N__9425),
            .I(N__9387));
    InMux I__2143 (
            .O(N__9424),
            .I(N__9384));
    InMux I__2142 (
            .O(N__9423),
            .I(N__9381));
    LocalMux I__2141 (
            .O(N__9420),
            .I(N__9374));
    LocalMux I__2140 (
            .O(N__9417),
            .I(N__9369));
    LocalMux I__2139 (
            .O(N__9414),
            .I(N__9369));
    InMux I__2138 (
            .O(N__9413),
            .I(N__9364));
    InMux I__2137 (
            .O(N__9412),
            .I(N__9364));
    InMux I__2136 (
            .O(N__9411),
            .I(N__9361));
    Span4Mux_v I__2135 (
            .O(N__9408),
            .I(N__9358));
    LocalMux I__2134 (
            .O(N__9403),
            .I(N__9349));
    LocalMux I__2133 (
            .O(N__9398),
            .I(N__9349));
    LocalMux I__2132 (
            .O(N__9393),
            .I(N__9349));
    LocalMux I__2131 (
            .O(N__9390),
            .I(N__9349));
    Span4Mux_h I__2130 (
            .O(N__9387),
            .I(N__9342));
    LocalMux I__2129 (
            .O(N__9384),
            .I(N__9342));
    LocalMux I__2128 (
            .O(N__9381),
            .I(N__9342));
    InMux I__2127 (
            .O(N__9380),
            .I(N__9337));
    InMux I__2126 (
            .O(N__9379),
            .I(N__9337));
    InMux I__2125 (
            .O(N__9378),
            .I(N__9332));
    InMux I__2124 (
            .O(N__9377),
            .I(N__9332));
    Span4Mux_v I__2123 (
            .O(N__9374),
            .I(N__9323));
    Span4Mux_h I__2122 (
            .O(N__9369),
            .I(N__9323));
    LocalMux I__2121 (
            .O(N__9364),
            .I(N__9323));
    LocalMux I__2120 (
            .O(N__9361),
            .I(N__9323));
    Span4Mux_v I__2119 (
            .O(N__9358),
            .I(N__9320));
    Span4Mux_h I__2118 (
            .O(N__9349),
            .I(N__9317));
    Span4Mux_h I__2117 (
            .O(N__9342),
            .I(N__9310));
    LocalMux I__2116 (
            .O(N__9337),
            .I(N__9310));
    LocalMux I__2115 (
            .O(N__9332),
            .I(N__9310));
    Odrv4 I__2114 (
            .O(N__9323),
            .I(CPU_CYCLE));
    Odrv4 I__2113 (
            .O(N__9320),
            .I(CPU_CYCLE));
    Odrv4 I__2112 (
            .O(N__9317),
            .I(CPU_CYCLE));
    Odrv4 I__2111 (
            .O(N__9310),
            .I(CPU_CYCLE));
    CascadeMux I__2110 (
            .O(N__9301),
            .I(N__9293));
    InMux I__2109 (
            .O(N__9300),
            .I(N__9288));
    InMux I__2108 (
            .O(N__9299),
            .I(N__9288));
    CascadeMux I__2107 (
            .O(N__9298),
            .I(N__9285));
    InMux I__2106 (
            .O(N__9297),
            .I(N__9282));
    InMux I__2105 (
            .O(N__9296),
            .I(N__9278));
    InMux I__2104 (
            .O(N__9293),
            .I(N__9275));
    LocalMux I__2103 (
            .O(N__9288),
            .I(N__9272));
    InMux I__2102 (
            .O(N__9285),
            .I(N__9269));
    LocalMux I__2101 (
            .O(N__9282),
            .I(N__9266));
    CascadeMux I__2100 (
            .O(N__9281),
            .I(N__9263));
    LocalMux I__2099 (
            .O(N__9278),
            .I(N__9256));
    LocalMux I__2098 (
            .O(N__9275),
            .I(N__9256));
    Span4Mux_h I__2097 (
            .O(N__9272),
            .I(N__9240));
    LocalMux I__2096 (
            .O(N__9269),
            .I(N__9240));
    Span4Mux_v I__2095 (
            .O(N__9266),
            .I(N__9233));
    InMux I__2094 (
            .O(N__9263),
            .I(N__9228));
    InMux I__2093 (
            .O(N__9262),
            .I(N__9228));
    InMux I__2092 (
            .O(N__9261),
            .I(N__9225));
    Span4Mux_v I__2091 (
            .O(N__9256),
            .I(N__9222));
    InMux I__2090 (
            .O(N__9255),
            .I(N__9213));
    InMux I__2089 (
            .O(N__9254),
            .I(N__9213));
    InMux I__2088 (
            .O(N__9253),
            .I(N__9213));
    InMux I__2087 (
            .O(N__9252),
            .I(N__9213));
    InMux I__2086 (
            .O(N__9251),
            .I(N__9204));
    InMux I__2085 (
            .O(N__9250),
            .I(N__9204));
    InMux I__2084 (
            .O(N__9249),
            .I(N__9204));
    InMux I__2083 (
            .O(N__9248),
            .I(N__9204));
    InMux I__2082 (
            .O(N__9247),
            .I(N__9199));
    InMux I__2081 (
            .O(N__9246),
            .I(N__9199));
    InMux I__2080 (
            .O(N__9245),
            .I(N__9196));
    Span4Mux_h I__2079 (
            .O(N__9240),
            .I(N__9193));
    InMux I__2078 (
            .O(N__9239),
            .I(N__9186));
    InMux I__2077 (
            .O(N__9238),
            .I(N__9186));
    InMux I__2076 (
            .O(N__9237),
            .I(N__9186));
    InMux I__2075 (
            .O(N__9236),
            .I(N__9183));
    Sp12to4 I__2074 (
            .O(N__9233),
            .I(N__9168));
    LocalMux I__2073 (
            .O(N__9228),
            .I(N__9168));
    LocalMux I__2072 (
            .O(N__9225),
            .I(N__9168));
    Sp12to4 I__2071 (
            .O(N__9222),
            .I(N__9168));
    LocalMux I__2070 (
            .O(N__9213),
            .I(N__9168));
    LocalMux I__2069 (
            .O(N__9204),
            .I(N__9168));
    LocalMux I__2068 (
            .O(N__9199),
            .I(N__9168));
    LocalMux I__2067 (
            .O(N__9196),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2066 (
            .O(N__9193),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2065 (
            .O(N__9186),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2064 (
            .O(N__9183),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2063 (
            .O(N__9168),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__2062 (
            .O(N__9157),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_ ));
    InMux I__2061 (
            .O(N__9154),
            .I(N__9151));
    LocalMux I__2060 (
            .O(N__9151),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__2059 (
            .O(N__9148),
            .I(N__9145));
    LocalMux I__2058 (
            .O(N__9145),
            .I(N__9142));
    Span4Mux_s3_v I__2057 (
            .O(N__9142),
            .I(N__9139));
    Span4Mux_v I__2056 (
            .O(N__9139),
            .I(N__9136));
    Span4Mux_v I__2055 (
            .O(N__9136),
            .I(N__9133));
    Span4Mux_h I__2054 (
            .O(N__9133),
            .I(N__9130));
    Odrv4 I__2053 (
            .O(N__9130),
            .I(CMA_c_0));
    CascadeMux I__2052 (
            .O(N__9127),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ));
    InMux I__2051 (
            .O(N__9124),
            .I(N__9121));
    LocalMux I__2050 (
            .O(N__9121),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2049 (
            .O(N__9118),
            .I(N__9115));
    LocalMux I__2048 (
            .O(N__9115),
            .I(N__9112));
    Odrv4 I__2047 (
            .O(N__9112),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2046 (
            .O(N__9109),
            .I(N__9103));
    InMux I__2045 (
            .O(N__9108),
            .I(N__9103));
    LocalMux I__2044 (
            .O(N__9103),
            .I(N__9100));
    Span4Mux_v I__2043 (
            .O(N__9100),
            .I(N__9097));
    Odrv4 I__2042 (
            .O(N__9097),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2041 (
            .O(N__9094),
            .I(N__9090));
    InMux I__2040 (
            .O(N__9093),
            .I(N__9087));
    LocalMux I__2039 (
            .O(N__9090),
            .I(N__9082));
    LocalMux I__2038 (
            .O(N__9087),
            .I(N__9073));
    ClkMux I__2037 (
            .O(N__9086),
            .I(N__9052));
    ClkMux I__2036 (
            .O(N__9085),
            .I(N__9052));
    Glb2LocalMux I__2035 (
            .O(N__9082),
            .I(N__9052));
    ClkMux I__2034 (
            .O(N__9081),
            .I(N__9052));
    ClkMux I__2033 (
            .O(N__9080),
            .I(N__9052));
    ClkMux I__2032 (
            .O(N__9079),
            .I(N__9052));
    ClkMux I__2031 (
            .O(N__9078),
            .I(N__9052));
    ClkMux I__2030 (
            .O(N__9077),
            .I(N__9052));
    ClkMux I__2029 (
            .O(N__9076),
            .I(N__9052));
    Glb2LocalMux I__2028 (
            .O(N__9073),
            .I(N__9052));
    GlobalMux I__2027 (
            .O(N__9052),
            .I(N__9049));
    gio2CtrlBuf I__2026 (
            .O(N__9049),
            .I(CLK40_PLL_g));
    InMux I__2025 (
            .O(N__9046),
            .I(N__9040));
    InMux I__2024 (
            .O(N__9045),
            .I(N__9040));
    LocalMux I__2023 (
            .O(N__9040),
            .I(N__9033));
    InMux I__2022 (
            .O(N__9039),
            .I(N__9028));
    InMux I__2021 (
            .O(N__9038),
            .I(N__9028));
    InMux I__2020 (
            .O(N__9037),
            .I(N__9025));
    InMux I__2019 (
            .O(N__9036),
            .I(N__9022));
    Odrv4 I__2018 (
            .O(N__9033),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2017 (
            .O(N__9028),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2016 (
            .O(N__9025),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2015 (
            .O(N__9022),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__2014 (
            .O(N__9013),
            .I(N__9010));
    InMux I__2013 (
            .O(N__9010),
            .I(N__9007));
    LocalMux I__2012 (
            .O(N__9007),
            .I(\U712_CYCLE_TERM.N_8 ));
    CascadeMux I__2011 (
            .O(N__9004),
            .I(N__9000));
    CascadeMux I__2010 (
            .O(N__9003),
            .I(N__8996));
    InMux I__2009 (
            .O(N__9000),
            .I(N__8986));
    InMux I__2008 (
            .O(N__8999),
            .I(N__8986));
    InMux I__2007 (
            .O(N__8996),
            .I(N__8981));
    InMux I__2006 (
            .O(N__8995),
            .I(N__8981));
    InMux I__2005 (
            .O(N__8994),
            .I(N__8978));
    InMux I__2004 (
            .O(N__8993),
            .I(N__8968));
    InMux I__2003 (
            .O(N__8992),
            .I(N__8968));
    InMux I__2002 (
            .O(N__8991),
            .I(N__8968));
    LocalMux I__2001 (
            .O(N__8986),
            .I(N__8965));
    LocalMux I__2000 (
            .O(N__8981),
            .I(N__8960));
    LocalMux I__1999 (
            .O(N__8978),
            .I(N__8960));
    InMux I__1998 (
            .O(N__8977),
            .I(N__8957));
    InMux I__1997 (
            .O(N__8976),
            .I(N__8954));
    InMux I__1996 (
            .O(N__8975),
            .I(N__8951));
    LocalMux I__1995 (
            .O(N__8968),
            .I(N__8946));
    Span4Mux_v I__1994 (
            .O(N__8965),
            .I(N__8937));
    Span4Mux_h I__1993 (
            .O(N__8960),
            .I(N__8937));
    LocalMux I__1992 (
            .O(N__8957),
            .I(N__8937));
    LocalMux I__1991 (
            .O(N__8954),
            .I(N__8937));
    LocalMux I__1990 (
            .O(N__8951),
            .I(N__8933));
    InMux I__1989 (
            .O(N__8950),
            .I(N__8928));
    InMux I__1988 (
            .O(N__8949),
            .I(N__8928));
    Span4Mux_v I__1987 (
            .O(N__8946),
            .I(N__8925));
    Span4Mux_v I__1986 (
            .O(N__8937),
            .I(N__8922));
    InMux I__1985 (
            .O(N__8936),
            .I(N__8919));
    Sp12to4 I__1984 (
            .O(N__8933),
            .I(N__8914));
    LocalMux I__1983 (
            .O(N__8928),
            .I(N__8914));
    Sp12to4 I__1982 (
            .O(N__8925),
            .I(N__8907));
    Sp12to4 I__1981 (
            .O(N__8922),
            .I(N__8907));
    LocalMux I__1980 (
            .O(N__8919),
            .I(N__8907));
    Span12Mux_v I__1979 (
            .O(N__8914),
            .I(N__8904));
    Span12Mux_h I__1978 (
            .O(N__8907),
            .I(N__8901));
    Span12Mux_h I__1977 (
            .O(N__8904),
            .I(N__8898));
    Odrv12 I__1976 (
            .O(N__8901),
            .I(RESETn_c));
    Odrv12 I__1975 (
            .O(N__8898),
            .I(RESETn_c));
    InMux I__1974 (
            .O(N__8893),
            .I(N__8888));
    InMux I__1973 (
            .O(N__8892),
            .I(N__8885));
    InMux I__1972 (
            .O(N__8891),
            .I(N__8882));
    LocalMux I__1971 (
            .O(N__8888),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1970 (
            .O(N__8885),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1969 (
            .O(N__8882),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1968 (
            .O(N__8875),
            .I(N__8871));
    InMux I__1967 (
            .O(N__8874),
            .I(N__8868));
    LocalMux I__1966 (
            .O(N__8871),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1965 (
            .O(N__8868),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__1964 (
            .O(N__8863),
            .I(N__8858));
    CascadeMux I__1963 (
            .O(N__8862),
            .I(N__8855));
    InMux I__1962 (
            .O(N__8861),
            .I(N__8851));
    InMux I__1961 (
            .O(N__8858),
            .I(N__8848));
    InMux I__1960 (
            .O(N__8855),
            .I(N__8845));
    InMux I__1959 (
            .O(N__8854),
            .I(N__8842));
    LocalMux I__1958 (
            .O(N__8851),
            .I(N__8838));
    LocalMux I__1957 (
            .O(N__8848),
            .I(N__8835));
    LocalMux I__1956 (
            .O(N__8845),
            .I(N__8830));
    LocalMux I__1955 (
            .O(N__8842),
            .I(N__8830));
    InMux I__1954 (
            .O(N__8841),
            .I(N__8827));
    Span4Mux_h I__1953 (
            .O(N__8838),
            .I(N__8824));
    Span4Mux_h I__1952 (
            .O(N__8835),
            .I(N__8821));
    Span4Mux_h I__1951 (
            .O(N__8830),
            .I(N__8818));
    LocalMux I__1950 (
            .O(N__8827),
            .I(CPU_TACK));
    Odrv4 I__1949 (
            .O(N__8824),
            .I(CPU_TACK));
    Odrv4 I__1948 (
            .O(N__8821),
            .I(CPU_TACK));
    Odrv4 I__1947 (
            .O(N__8818),
            .I(CPU_TACK));
    CascadeMux I__1946 (
            .O(N__8809),
            .I(\U712_CYCLE_TERM.N_227_i_0_0_cascade_ ));
    CascadeMux I__1945 (
            .O(N__8806),
            .I(N__8801));
    InMux I__1944 (
            .O(N__8805),
            .I(N__8796));
    InMux I__1943 (
            .O(N__8804),
            .I(N__8793));
    InMux I__1942 (
            .O(N__8801),
            .I(N__8790));
    InMux I__1941 (
            .O(N__8800),
            .I(N__8785));
    InMux I__1940 (
            .O(N__8799),
            .I(N__8785));
    LocalMux I__1939 (
            .O(N__8796),
            .I(N__8780));
    LocalMux I__1938 (
            .O(N__8793),
            .I(N__8780));
    LocalMux I__1937 (
            .O(N__8790),
            .I(REG_TACK));
    LocalMux I__1936 (
            .O(N__8785),
            .I(REG_TACK));
    Odrv4 I__1935 (
            .O(N__8780),
            .I(REG_TACK));
    CascadeMux I__1934 (
            .O(N__8773),
            .I(\U712_CYCLE_TERM.N_227_i_0_en_cascade_ ));
    IoInMux I__1933 (
            .O(N__8770),
            .I(N__8767));
    LocalMux I__1932 (
            .O(N__8767),
            .I(N__8764));
    Span12Mux_s1_v I__1931 (
            .O(N__8764),
            .I(N__8760));
    InMux I__1930 (
            .O(N__8763),
            .I(N__8757));
    Odrv12 I__1929 (
            .O(N__8760),
            .I(RESETn_c_i));
    LocalMux I__1928 (
            .O(N__8757),
            .I(RESETn_c_i));
    CEMux I__1927 (
            .O(N__8752),
            .I(N__8749));
    LocalMux I__1926 (
            .O(N__8749),
            .I(N__8746));
    Odrv4 I__1925 (
            .O(N__8746),
            .I(\U712_CYCLE_TERM.N_227_i_0_en_0 ));
    IoInMux I__1924 (
            .O(N__8743),
            .I(N__8740));
    LocalMux I__1923 (
            .O(N__8740),
            .I(N__8737));
    Span4Mux_s2_v I__1922 (
            .O(N__8737),
            .I(N__8734));
    Sp12to4 I__1921 (
            .O(N__8734),
            .I(N__8731));
    Span12Mux_h I__1920 (
            .O(N__8731),
            .I(N__8728));
    Odrv12 I__1919 (
            .O(N__8728),
            .I(CRCSn_c));
    IoInMux I__1918 (
            .O(N__8725),
            .I(N__8722));
    LocalMux I__1917 (
            .O(N__8722),
            .I(N__8719));
    Span4Mux_s2_v I__1916 (
            .O(N__8719),
            .I(N__8716));
    Span4Mux_v I__1915 (
            .O(N__8716),
            .I(N__8713));
    Span4Mux_v I__1914 (
            .O(N__8713),
            .I(N__8710));
    Span4Mux_h I__1913 (
            .O(N__8710),
            .I(N__8707));
    Odrv4 I__1912 (
            .O(N__8707),
            .I(CMA_c_10));
    IoInMux I__1911 (
            .O(N__8704),
            .I(N__8700));
    InMux I__1910 (
            .O(N__8703),
            .I(N__8697));
    LocalMux I__1909 (
            .O(N__8700),
            .I(N__8694));
    LocalMux I__1908 (
            .O(N__8697),
            .I(N__8691));
    Span12Mux_s11_v I__1907 (
            .O(N__8694),
            .I(N__8688));
    Span4Mux_h I__1906 (
            .O(N__8691),
            .I(N__8685));
    Odrv12 I__1905 (
            .O(N__8688),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1904 (
            .O(N__8685),
            .I(CONSTANT_ONE_NET));
    InMux I__1903 (
            .O(N__8680),
            .I(N__8677));
    LocalMux I__1902 (
            .O(N__8677),
            .I(N__8674));
    Odrv12 I__1901 (
            .O(N__8674),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1900 (
            .O(N__8671),
            .I(N__8668));
    LocalMux I__1899 (
            .O(N__8668),
            .I(N__8665));
    Span4Mux_v I__1898 (
            .O(N__8665),
            .I(N__8662));
    Span4Mux_v I__1897 (
            .O(N__8662),
            .I(N__8659));
    Sp12to4 I__1896 (
            .O(N__8659),
            .I(N__8656));
    Span12Mux_h I__1895 (
            .O(N__8656),
            .I(N__8653));
    Odrv12 I__1894 (
            .O(N__8653),
            .I(A_c_6));
    InMux I__1893 (
            .O(N__8650),
            .I(N__8647));
    LocalMux I__1892 (
            .O(N__8647),
            .I(N__8644));
    Span12Mux_v I__1891 (
            .O(N__8644),
            .I(N__8641));
    Span12Mux_h I__1890 (
            .O(N__8641),
            .I(N__8638));
    Odrv12 I__1889 (
            .O(N__8638),
            .I(A_c_13));
    CascadeMux I__1888 (
            .O(N__8635),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    CascadeMux I__1887 (
            .O(N__8632),
            .I(N__8629));
    InMux I__1886 (
            .O(N__8629),
            .I(N__8626));
    LocalMux I__1885 (
            .O(N__8626),
            .I(N__8623));
    Odrv12 I__1884 (
            .O(N__8623),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1883 (
            .O(N__8620),
            .I(N__8615));
    InMux I__1882 (
            .O(N__8619),
            .I(N__8612));
    InMux I__1881 (
            .O(N__8618),
            .I(N__8608));
    LocalMux I__1880 (
            .O(N__8615),
            .I(N__8601));
    LocalMux I__1879 (
            .O(N__8612),
            .I(N__8601));
    InMux I__1878 (
            .O(N__8611),
            .I(N__8597));
    LocalMux I__1877 (
            .O(N__8608),
            .I(N__8594));
    InMux I__1876 (
            .O(N__8607),
            .I(N__8591));
    InMux I__1875 (
            .O(N__8606),
            .I(N__8588));
    Span4Mux_v I__1874 (
            .O(N__8601),
            .I(N__8585));
    InMux I__1873 (
            .O(N__8600),
            .I(N__8582));
    LocalMux I__1872 (
            .O(N__8597),
            .I(N__8575));
    Span4Mux_h I__1871 (
            .O(N__8594),
            .I(N__8575));
    LocalMux I__1870 (
            .O(N__8591),
            .I(N__8575));
    LocalMux I__1869 (
            .O(N__8588),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1868 (
            .O(N__8585),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__1867 (
            .O(N__8582),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__1866 (
            .O(N__8575),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    CascadeMux I__1865 (
            .O(N__8566),
            .I(N__8561));
    InMux I__1864 (
            .O(N__8565),
            .I(N__8558));
    CascadeMux I__1863 (
            .O(N__8564),
            .I(N__8555));
    InMux I__1862 (
            .O(N__8561),
            .I(N__8551));
    LocalMux I__1861 (
            .O(N__8558),
            .I(N__8548));
    InMux I__1860 (
            .O(N__8555),
            .I(N__8545));
    CascadeMux I__1859 (
            .O(N__8554),
            .I(N__8542));
    LocalMux I__1858 (
            .O(N__8551),
            .I(N__8538));
    Span4Mux_h I__1857 (
            .O(N__8548),
            .I(N__8535));
    LocalMux I__1856 (
            .O(N__8545),
            .I(N__8532));
    InMux I__1855 (
            .O(N__8542),
            .I(N__8529));
    InMux I__1854 (
            .O(N__8541),
            .I(N__8526));
    Span12Mux_h I__1853 (
            .O(N__8538),
            .I(N__8523));
    Span4Mux_h I__1852 (
            .O(N__8535),
            .I(N__8520));
    Span4Mux_h I__1851 (
            .O(N__8532),
            .I(N__8515));
    LocalMux I__1850 (
            .O(N__8529),
            .I(N__8515));
    LocalMux I__1849 (
            .O(N__8526),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv12 I__1848 (
            .O(N__8523),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1847 (
            .O(N__8520),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1846 (
            .O(N__8515),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__1845 (
            .O(N__8506),
            .I(N__8501));
    InMux I__1844 (
            .O(N__8505),
            .I(N__8498));
    InMux I__1843 (
            .O(N__8504),
            .I(N__8494));
    LocalMux I__1842 (
            .O(N__8501),
            .I(N__8486));
    LocalMux I__1841 (
            .O(N__8498),
            .I(N__8486));
    InMux I__1840 (
            .O(N__8497),
            .I(N__8483));
    LocalMux I__1839 (
            .O(N__8494),
            .I(N__8480));
    InMux I__1838 (
            .O(N__8493),
            .I(N__8475));
    InMux I__1837 (
            .O(N__8492),
            .I(N__8475));
    InMux I__1836 (
            .O(N__8491),
            .I(N__8472));
    Span4Mux_v I__1835 (
            .O(N__8486),
            .I(N__8469));
    LocalMux I__1834 (
            .O(N__8483),
            .I(N__8460));
    Span4Mux_h I__1833 (
            .O(N__8480),
            .I(N__8460));
    LocalMux I__1832 (
            .O(N__8475),
            .I(N__8460));
    LocalMux I__1831 (
            .O(N__8472),
            .I(N__8460));
    Odrv4 I__1830 (
            .O(N__8469),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__1829 (
            .O(N__8460),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    CascadeMux I__1828 (
            .O(N__8455),
            .I(N__8450));
    IoInMux I__1827 (
            .O(N__8454),
            .I(N__8447));
    InMux I__1826 (
            .O(N__8453),
            .I(N__8442));
    InMux I__1825 (
            .O(N__8450),
            .I(N__8442));
    LocalMux I__1824 (
            .O(N__8447),
            .I(N__8439));
    LocalMux I__1823 (
            .O(N__8442),
            .I(N__8436));
    Span12Mux_s3_h I__1822 (
            .O(N__8439),
            .I(N__8433));
    Span4Mux_h I__1821 (
            .O(N__8436),
            .I(N__8430));
    Span12Mux_v I__1820 (
            .O(N__8433),
            .I(N__8427));
    Sp12to4 I__1819 (
            .O(N__8430),
            .I(N__8424));
    Span12Mux_h I__1818 (
            .O(N__8427),
            .I(N__8421));
    Span12Mux_v I__1817 (
            .O(N__8424),
            .I(N__8418));
    Odrv12 I__1816 (
            .O(N__8421),
            .I(CLK40_PLL));
    Odrv12 I__1815 (
            .O(N__8418),
            .I(CLK40_PLL));
    IoInMux I__1814 (
            .O(N__8413),
            .I(N__8410));
    LocalMux I__1813 (
            .O(N__8410),
            .I(N__8407));
    IoSpan4Mux I__1812 (
            .O(N__8407),
            .I(N__8404));
    Span4Mux_s2_h I__1811 (
            .O(N__8404),
            .I(N__8401));
    Sp12to4 I__1810 (
            .O(N__8401),
            .I(N__8398));
    Span12Mux_h I__1809 (
            .O(N__8398),
            .I(N__8394));
    InMux I__1808 (
            .O(N__8397),
            .I(N__8391));
    Odrv12 I__1807 (
            .O(N__8394),
            .I(TACK_OUTn));
    LocalMux I__1806 (
            .O(N__8391),
            .I(TACK_OUTn));
    InMux I__1805 (
            .O(N__8386),
            .I(N__8382));
    InMux I__1804 (
            .O(N__8385),
            .I(N__8379));
    LocalMux I__1803 (
            .O(N__8382),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__1802 (
            .O(N__8379),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1801 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__1800 (
            .O(N__8371),
            .I(N__8366));
    InMux I__1799 (
            .O(N__8370),
            .I(N__8363));
    InMux I__1798 (
            .O(N__8369),
            .I(N__8360));
    Odrv12 I__1797 (
            .O(N__8366),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1796 (
            .O(N__8363),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1795 (
            .O(N__8360),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1794 (
            .O(N__8353),
            .I(N__8350));
    LocalMux I__1793 (
            .O(N__8350),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__1792 (
            .O(N__8347),
            .I(N__8344));
    InMux I__1791 (
            .O(N__8344),
            .I(N__8341));
    LocalMux I__1790 (
            .O(N__8341),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ));
    InMux I__1789 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__1788 (
            .O(N__8335),
            .I(TACK_EN_i_ess));
    IoInMux I__1787 (
            .O(N__8332),
            .I(N__8329));
    LocalMux I__1786 (
            .O(N__8329),
            .I(N__8326));
    IoSpan4Mux I__1785 (
            .O(N__8326),
            .I(N__8323));
    Sp12to4 I__1784 (
            .O(N__8323),
            .I(N__8320));
    Span12Mux_s9_v I__1783 (
            .O(N__8320),
            .I(N__8317));
    Odrv12 I__1782 (
            .O(N__8317),
            .I(RASn_c));
    IoInMux I__1781 (
            .O(N__8314),
            .I(N__8311));
    LocalMux I__1780 (
            .O(N__8311),
            .I(N__8308));
    Span12Mux_s4_h I__1779 (
            .O(N__8308),
            .I(N__8305));
    Span12Mux_h I__1778 (
            .O(N__8305),
            .I(N__8302));
    Odrv12 I__1777 (
            .O(N__8302),
            .I(WEn_c));
    CascadeMux I__1776 (
            .O(N__8299),
            .I(N__8295));
    InMux I__1775 (
            .O(N__8298),
            .I(N__8290));
    InMux I__1774 (
            .O(N__8295),
            .I(N__8290));
    LocalMux I__1773 (
            .O(N__8290),
            .I(N__8287));
    Span4Mux_v I__1772 (
            .O(N__8287),
            .I(N__8282));
    InMux I__1771 (
            .O(N__8286),
            .I(N__8277));
    InMux I__1770 (
            .O(N__8285),
            .I(N__8277));
    Odrv4 I__1769 (
            .O(N__8282),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1768 (
            .O(N__8277),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1767 (
            .O(N__8272),
            .I(N__8269));
    LocalMux I__1766 (
            .O(N__8269),
            .I(N__8266));
    Sp12to4 I__1765 (
            .O(N__8266),
            .I(N__8263));
    Span12Mux_v I__1764 (
            .O(N__8263),
            .I(N__8260));
    Span12Mux_h I__1763 (
            .O(N__8260),
            .I(N__8257));
    Odrv12 I__1762 (
            .O(N__8257),
            .I(A_c_19));
    IoInMux I__1761 (
            .O(N__8254),
            .I(N__8251));
    LocalMux I__1760 (
            .O(N__8251),
            .I(N__8248));
    Span12Mux_s5_h I__1759 (
            .O(N__8248),
            .I(N__8245));
    Span12Mux_h I__1758 (
            .O(N__8245),
            .I(N__8242));
    Odrv12 I__1757 (
            .O(N__8242),
            .I(CMA_c_9));
    InMux I__1756 (
            .O(N__8239),
            .I(N__8236));
    LocalMux I__1755 (
            .O(N__8236),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1754 (
            .O(N__8233),
            .I(N__8230));
    LocalMux I__1753 (
            .O(N__8230),
            .I(N__8227));
    IoSpan4Mux I__1752 (
            .O(N__8227),
            .I(N__8224));
    Span4Mux_s3_h I__1751 (
            .O(N__8224),
            .I(N__8221));
    Sp12to4 I__1750 (
            .O(N__8221),
            .I(N__8218));
    Span12Mux_h I__1749 (
            .O(N__8218),
            .I(N__8215));
    Odrv12 I__1748 (
            .O(N__8215),
            .I(CMA_c_5));
    InMux I__1747 (
            .O(N__8212),
            .I(N__8209));
    LocalMux I__1746 (
            .O(N__8209),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1745 (
            .O(N__8206),
            .I(N__8203));
    LocalMux I__1744 (
            .O(N__8203),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1743 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__1742 (
            .O(N__8197),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__1741 (
            .O(N__8194),
            .I(N__8191));
    InMux I__1740 (
            .O(N__8191),
            .I(N__8188));
    LocalMux I__1739 (
            .O(N__8188),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__1738 (
            .O(N__8185),
            .I(N__8182));
    LocalMux I__1737 (
            .O(N__8182),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1736 (
            .O(N__8179),
            .I(N__8176));
    LocalMux I__1735 (
            .O(N__8176),
            .I(N__8173));
    Span4Mux_s3_v I__1734 (
            .O(N__8173),
            .I(N__8170));
    Span4Mux_v I__1733 (
            .O(N__8170),
            .I(N__8167));
    Span4Mux_v I__1732 (
            .O(N__8167),
            .I(N__8164));
    Odrv4 I__1731 (
            .O(N__8164),
            .I(CMA_c_1));
    InMux I__1730 (
            .O(N__8161),
            .I(N__8158));
    LocalMux I__1729 (
            .O(N__8158),
            .I(N__8155));
    Odrv4 I__1728 (
            .O(N__8155),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1727 (
            .O(N__8152),
            .I(N__8149));
    LocalMux I__1726 (
            .O(N__8149),
            .I(N__8146));
    Span4Mux_v I__1725 (
            .O(N__8146),
            .I(N__8143));
    Odrv4 I__1724 (
            .O(N__8143),
            .I(DBRn_c_i));
    InMux I__1723 (
            .O(N__8140),
            .I(N__8136));
    InMux I__1722 (
            .O(N__8139),
            .I(N__8133));
    LocalMux I__1721 (
            .O(N__8136),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    LocalMux I__1720 (
            .O(N__8133),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__1719 (
            .O(N__8128),
            .I(N__8124));
    InMux I__1718 (
            .O(N__8127),
            .I(N__8121));
    LocalMux I__1717 (
            .O(N__8124),
            .I(N__8117));
    LocalMux I__1716 (
            .O(N__8121),
            .I(N__8114));
    InMux I__1715 (
            .O(N__8120),
            .I(N__8111));
    Span4Mux_v I__1714 (
            .O(N__8117),
            .I(N__8108));
    Span4Mux_v I__1713 (
            .O(N__8114),
            .I(N__8103));
    LocalMux I__1712 (
            .O(N__8111),
            .I(N__8103));
    Span4Mux_v I__1711 (
            .O(N__8108),
            .I(N__8098));
    Span4Mux_v I__1710 (
            .O(N__8103),
            .I(N__8098));
    Sp12to4 I__1709 (
            .O(N__8098),
            .I(N__8095));
    Span12Mux_h I__1708 (
            .O(N__8095),
            .I(N__8092));
    Odrv12 I__1707 (
            .O(N__8092),
            .I(DBRn_c));
    InMux I__1706 (
            .O(N__8089),
            .I(N__8086));
    LocalMux I__1705 (
            .O(N__8086),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_0 ));
    InMux I__1704 (
            .O(N__8083),
            .I(N__8079));
    InMux I__1703 (
            .O(N__8082),
            .I(N__8075));
    LocalMux I__1702 (
            .O(N__8079),
            .I(N__8072));
    CascadeMux I__1701 (
            .O(N__8078),
            .I(N__8069));
    LocalMux I__1700 (
            .O(N__8075),
            .I(N__8064));
    Span4Mux_h I__1699 (
            .O(N__8072),
            .I(N__8064));
    InMux I__1698 (
            .O(N__8069),
            .I(N__8061));
    Odrv4 I__1697 (
            .O(N__8064),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    LocalMux I__1696 (
            .O(N__8061),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    InMux I__1695 (
            .O(N__8056),
            .I(N__8053));
    LocalMux I__1694 (
            .O(N__8053),
            .I(N__8049));
    InMux I__1693 (
            .O(N__8052),
            .I(N__8046));
    Span4Mux_v I__1692 (
            .O(N__8049),
            .I(N__8042));
    LocalMux I__1691 (
            .O(N__8046),
            .I(N__8039));
    InMux I__1690 (
            .O(N__8045),
            .I(N__8036));
    Odrv4 I__1689 (
            .O(N__8042),
            .I(REG_CYCLE));
    Odrv4 I__1688 (
            .O(N__8039),
            .I(REG_CYCLE));
    LocalMux I__1687 (
            .O(N__8036),
            .I(REG_CYCLE));
    IoInMux I__1686 (
            .O(N__8029),
            .I(N__8026));
    LocalMux I__1685 (
            .O(N__8026),
            .I(N__8023));
    Span4Mux_s0_v I__1684 (
            .O(N__8023),
            .I(N__8020));
    Span4Mux_v I__1683 (
            .O(N__8020),
            .I(N__8017));
    Span4Mux_v I__1682 (
            .O(N__8017),
            .I(N__8014));
    Sp12to4 I__1681 (
            .O(N__8014),
            .I(N__8011));
    Span12Mux_s11_h I__1680 (
            .O(N__8011),
            .I(N__8008));
    Odrv12 I__1679 (
            .O(N__8008),
            .I(DRDENn_c));
    IoInMux I__1678 (
            .O(N__8005),
            .I(N__8002));
    LocalMux I__1677 (
            .O(N__8002),
            .I(N__7999));
    IoSpan4Mux I__1676 (
            .O(N__7999),
            .I(N__7996));
    Span4Mux_s3_v I__1675 (
            .O(N__7996),
            .I(N__7993));
    Span4Mux_v I__1674 (
            .O(N__7993),
            .I(N__7990));
    Odrv4 I__1673 (
            .O(N__7990),
            .I(N_118_i));
    InMux I__1672 (
            .O(N__7987),
            .I(N__7978));
    InMux I__1671 (
            .O(N__7986),
            .I(N__7975));
    InMux I__1670 (
            .O(N__7985),
            .I(N__7972));
    InMux I__1669 (
            .O(N__7984),
            .I(N__7969));
    InMux I__1668 (
            .O(N__7983),
            .I(N__7964));
    InMux I__1667 (
            .O(N__7982),
            .I(N__7964));
    InMux I__1666 (
            .O(N__7981),
            .I(N__7961));
    LocalMux I__1665 (
            .O(N__7978),
            .I(N__7957));
    LocalMux I__1664 (
            .O(N__7975),
            .I(N__7950));
    LocalMux I__1663 (
            .O(N__7972),
            .I(N__7950));
    LocalMux I__1662 (
            .O(N__7969),
            .I(N__7950));
    LocalMux I__1661 (
            .O(N__7964),
            .I(N__7945));
    LocalMux I__1660 (
            .O(N__7961),
            .I(N__7945));
    InMux I__1659 (
            .O(N__7960),
            .I(N__7942));
    Span4Mux_v I__1658 (
            .O(N__7957),
            .I(N__7937));
    Span4Mux_v I__1657 (
            .O(N__7950),
            .I(N__7937));
    Span4Mux_h I__1656 (
            .O(N__7945),
            .I(N__7932));
    LocalMux I__1655 (
            .O(N__7942),
            .I(N__7932));
    Span4Mux_h I__1654 (
            .O(N__7937),
            .I(N__7929));
    Span4Mux_v I__1653 (
            .O(N__7932),
            .I(N__7926));
    Sp12to4 I__1652 (
            .O(N__7929),
            .I(N__7921));
    Sp12to4 I__1651 (
            .O(N__7926),
            .I(N__7921));
    Odrv12 I__1650 (
            .O(N__7921),
            .I(A_c_0));
    IoInMux I__1649 (
            .O(N__7918),
            .I(N__7915));
    LocalMux I__1648 (
            .O(N__7915),
            .I(N__7912));
    Span4Mux_s3_v I__1647 (
            .O(N__7912),
            .I(N__7909));
    Span4Mux_h I__1646 (
            .O(N__7909),
            .I(N__7906));
    Odrv4 I__1645 (
            .O(N__7906),
            .I(U712_BYTE_ENABLE_UUBE_i));
    IoInMux I__1644 (
            .O(N__7903),
            .I(N__7900));
    LocalMux I__1643 (
            .O(N__7900),
            .I(N__7897));
    Span4Mux_s2_v I__1642 (
            .O(N__7897),
            .I(N__7894));
    Span4Mux_h I__1641 (
            .O(N__7894),
            .I(N__7891));
    Span4Mux_v I__1640 (
            .O(N__7891),
            .I(N__7888));
    Odrv4 I__1639 (
            .O(N__7888),
            .I(LLBEn_c));
    InMux I__1638 (
            .O(N__7885),
            .I(N__7881));
    InMux I__1637 (
            .O(N__7884),
            .I(N__7878));
    LocalMux I__1636 (
            .O(N__7881),
            .I(N__7871));
    LocalMux I__1635 (
            .O(N__7878),
            .I(N__7871));
    InMux I__1634 (
            .O(N__7877),
            .I(N__7866));
    InMux I__1633 (
            .O(N__7876),
            .I(N__7866));
    Span4Mux_v I__1632 (
            .O(N__7871),
            .I(N__7861));
    LocalMux I__1631 (
            .O(N__7866),
            .I(N__7861));
    Odrv4 I__1630 (
            .O(N__7861),
            .I(N_386));
    CascadeMux I__1629 (
            .O(N__7858),
            .I(N__7854));
    InMux I__1628 (
            .O(N__7857),
            .I(N__7851));
    InMux I__1627 (
            .O(N__7854),
            .I(N__7848));
    LocalMux I__1626 (
            .O(N__7851),
            .I(N__7840));
    LocalMux I__1625 (
            .O(N__7848),
            .I(N__7840));
    InMux I__1624 (
            .O(N__7847),
            .I(N__7835));
    InMux I__1623 (
            .O(N__7846),
            .I(N__7835));
    InMux I__1622 (
            .O(N__7845),
            .I(N__7832));
    Span4Mux_v I__1621 (
            .O(N__7840),
            .I(N__7826));
    LocalMux I__1620 (
            .O(N__7835),
            .I(N__7826));
    LocalMux I__1619 (
            .O(N__7832),
            .I(N__7823));
    InMux I__1618 (
            .O(N__7831),
            .I(N__7820));
    Span4Mux_h I__1617 (
            .O(N__7826),
            .I(N__7817));
    Span12Mux_h I__1616 (
            .O(N__7823),
            .I(N__7814));
    LocalMux I__1615 (
            .O(N__7820),
            .I(N__7811));
    Span4Mux_v I__1614 (
            .O(N__7817),
            .I(N__7808));
    Span12Mux_v I__1613 (
            .O(N__7814),
            .I(N__7805));
    Span12Mux_v I__1612 (
            .O(N__7811),
            .I(N__7800));
    Sp12to4 I__1611 (
            .O(N__7808),
            .I(N__7800));
    Odrv12 I__1610 (
            .O(N__7805),
            .I(SIZ_c_0));
    Odrv12 I__1609 (
            .O(N__7800),
            .I(SIZ_c_0));
    InMux I__1608 (
            .O(N__7795),
            .I(N__7787));
    InMux I__1607 (
            .O(N__7794),
            .I(N__7780));
    InMux I__1606 (
            .O(N__7793),
            .I(N__7780));
    InMux I__1605 (
            .O(N__7792),
            .I(N__7780));
    CascadeMux I__1604 (
            .O(N__7791),
            .I(N__7776));
    CascadeMux I__1603 (
            .O(N__7790),
            .I(N__7773));
    LocalMux I__1602 (
            .O(N__7787),
            .I(N__7770));
    LocalMux I__1601 (
            .O(N__7780),
            .I(N__7767));
    InMux I__1600 (
            .O(N__7779),
            .I(N__7760));
    InMux I__1599 (
            .O(N__7776),
            .I(N__7760));
    InMux I__1598 (
            .O(N__7773),
            .I(N__7760));
    Span4Mux_v I__1597 (
            .O(N__7770),
            .I(N__7757));
    Span4Mux_v I__1596 (
            .O(N__7767),
            .I(N__7754));
    LocalMux I__1595 (
            .O(N__7760),
            .I(N__7751));
    Span4Mux_v I__1594 (
            .O(N__7757),
            .I(N__7747));
    Span4Mux_v I__1593 (
            .O(N__7754),
            .I(N__7742));
    Span4Mux_v I__1592 (
            .O(N__7751),
            .I(N__7742));
    InMux I__1591 (
            .O(N__7750),
            .I(N__7739));
    Sp12to4 I__1590 (
            .O(N__7747),
            .I(N__7732));
    Sp12to4 I__1589 (
            .O(N__7742),
            .I(N__7732));
    LocalMux I__1588 (
            .O(N__7739),
            .I(N__7732));
    Span12Mux_h I__1587 (
            .O(N__7732),
            .I(N__7729));
    Odrv12 I__1586 (
            .O(N__7729),
            .I(A_c_1));
    InMux I__1585 (
            .O(N__7726),
            .I(N__7723));
    LocalMux I__1584 (
            .O(N__7723),
            .I(N__7719));
    InMux I__1583 (
            .O(N__7722),
            .I(N__7716));
    Span4Mux_v I__1582 (
            .O(N__7719),
            .I(N__7712));
    LocalMux I__1581 (
            .O(N__7716),
            .I(N__7705));
    InMux I__1580 (
            .O(N__7715),
            .I(N__7702));
    Span4Mux_v I__1579 (
            .O(N__7712),
            .I(N__7699));
    InMux I__1578 (
            .O(N__7711),
            .I(N__7696));
    InMux I__1577 (
            .O(N__7710),
            .I(N__7693));
    InMux I__1576 (
            .O(N__7709),
            .I(N__7688));
    InMux I__1575 (
            .O(N__7708),
            .I(N__7688));
    Sp12to4 I__1574 (
            .O(N__7705),
            .I(N__7683));
    LocalMux I__1573 (
            .O(N__7702),
            .I(N__7683));
    Span4Mux_v I__1572 (
            .O(N__7699),
            .I(N__7680));
    LocalMux I__1571 (
            .O(N__7696),
            .I(N__7673));
    LocalMux I__1570 (
            .O(N__7693),
            .I(N__7673));
    LocalMux I__1569 (
            .O(N__7688),
            .I(N__7673));
    Span12Mux_h I__1568 (
            .O(N__7683),
            .I(N__7670));
    Sp12to4 I__1567 (
            .O(N__7680),
            .I(N__7665));
    Span12Mux_v I__1566 (
            .O(N__7673),
            .I(N__7665));
    Span12Mux_v I__1565 (
            .O(N__7670),
            .I(N__7660));
    Span12Mux_h I__1564 (
            .O(N__7665),
            .I(N__7660));
    Odrv12 I__1563 (
            .O(N__7660),
            .I(SIZ_c_1));
    IoInMux I__1562 (
            .O(N__7657),
            .I(N__7654));
    LocalMux I__1561 (
            .O(N__7654),
            .I(N__7651));
    Span4Mux_s2_v I__1560 (
            .O(N__7651),
            .I(N__7648));
    Span4Mux_v I__1559 (
            .O(N__7648),
            .I(N__7645));
    Sp12to4 I__1558 (
            .O(N__7645),
            .I(N__7642));
    Odrv12 I__1557 (
            .O(N__7642),
            .I(UMBEn_c));
    InMux I__1556 (
            .O(N__7639),
            .I(N__7636));
    LocalMux I__1555 (
            .O(N__7636),
            .I(N__7633));
    Sp12to4 I__1554 (
            .O(N__7633),
            .I(N__7630));
    Span12Mux_v I__1553 (
            .O(N__7630),
            .I(N__7627));
    Span12Mux_h I__1552 (
            .O(N__7627),
            .I(N__7624));
    Odrv12 I__1551 (
            .O(N__7624),
            .I(A_c_17));
    IoInMux I__1550 (
            .O(N__7621),
            .I(N__7618));
    LocalMux I__1549 (
            .O(N__7618),
            .I(N__7615));
    IoSpan4Mux I__1548 (
            .O(N__7615),
            .I(N__7612));
    Span4Mux_s3_h I__1547 (
            .O(N__7612),
            .I(N__7609));
    Sp12to4 I__1546 (
            .O(N__7609),
            .I(N__7606));
    Span12Mux_h I__1545 (
            .O(N__7606),
            .I(N__7603));
    Odrv12 I__1544 (
            .O(N__7603),
            .I(CMA_c_8));
    CascadeMux I__1543 (
            .O(N__7600),
            .I(N__7596));
    InMux I__1542 (
            .O(N__7599),
            .I(N__7590));
    InMux I__1541 (
            .O(N__7596),
            .I(N__7587));
    InMux I__1540 (
            .O(N__7595),
            .I(N__7584));
    InMux I__1539 (
            .O(N__7594),
            .I(N__7581));
    InMux I__1538 (
            .O(N__7593),
            .I(N__7578));
    LocalMux I__1537 (
            .O(N__7590),
            .I(REG_WRITE_CYCLE));
    LocalMux I__1536 (
            .O(N__7587),
            .I(REG_WRITE_CYCLE));
    LocalMux I__1535 (
            .O(N__7584),
            .I(REG_WRITE_CYCLE));
    LocalMux I__1534 (
            .O(N__7581),
            .I(REG_WRITE_CYCLE));
    LocalMux I__1533 (
            .O(N__7578),
            .I(REG_WRITE_CYCLE));
    InMux I__1532 (
            .O(N__7567),
            .I(N__7563));
    InMux I__1531 (
            .O(N__7566),
            .I(N__7559));
    LocalMux I__1530 (
            .O(N__7563),
            .I(N__7556));
    InMux I__1529 (
            .O(N__7562),
            .I(N__7552));
    LocalMux I__1528 (
            .O(N__7559),
            .I(N__7549));
    Span4Mux_v I__1527 (
            .O(N__7556),
            .I(N__7546));
    InMux I__1526 (
            .O(N__7555),
            .I(N__7543));
    LocalMux I__1525 (
            .O(N__7552),
            .I(N__7540));
    Sp12to4 I__1524 (
            .O(N__7549),
            .I(N__7533));
    Sp12to4 I__1523 (
            .O(N__7546),
            .I(N__7533));
    LocalMux I__1522 (
            .O(N__7543),
            .I(N__7533));
    Span4Mux_v I__1521 (
            .O(N__7540),
            .I(N__7530));
    Span12Mux_h I__1520 (
            .O(N__7533),
            .I(N__7527));
    Sp12to4 I__1519 (
            .O(N__7530),
            .I(N__7524));
    Span12Mux_v I__1518 (
            .O(N__7527),
            .I(N__7521));
    Span12Mux_h I__1517 (
            .O(N__7524),
            .I(N__7518));
    Odrv12 I__1516 (
            .O(N__7521),
            .I(RnW_c));
    Odrv12 I__1515 (
            .O(N__7518),
            .I(RnW_c));
    InMux I__1514 (
            .O(N__7513),
            .I(N__7510));
    LocalMux I__1513 (
            .O(N__7510),
            .I(N__7507));
    Odrv4 I__1512 (
            .O(N__7507),
            .I(\U712_REG_SM.UDSn_7_iv_i_0 ));
    InMux I__1511 (
            .O(N__7504),
            .I(N__7501));
    LocalMux I__1510 (
            .O(N__7501),
            .I(\U712_REG_SM.N_245 ));
    InMux I__1509 (
            .O(N__7498),
            .I(N__7495));
    LocalMux I__1508 (
            .O(N__7495),
            .I(\U712_REG_SM.un15_0_i_0_0_0 ));
    InMux I__1507 (
            .O(N__7492),
            .I(N__7487));
    InMux I__1506 (
            .O(N__7491),
            .I(N__7482));
    InMux I__1505 (
            .O(N__7490),
            .I(N__7482));
    LocalMux I__1504 (
            .O(N__7487),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    LocalMux I__1503 (
            .O(N__7482),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    CascadeMux I__1502 (
            .O(N__7477),
            .I(N__7474));
    InMux I__1501 (
            .O(N__7474),
            .I(N__7468));
    CascadeMux I__1500 (
            .O(N__7473),
            .I(N__7463));
    CascadeMux I__1499 (
            .O(N__7472),
            .I(N__7459));
    InMux I__1498 (
            .O(N__7471),
            .I(N__7456));
    LocalMux I__1497 (
            .O(N__7468),
            .I(N__7453));
    InMux I__1496 (
            .O(N__7467),
            .I(N__7448));
    InMux I__1495 (
            .O(N__7466),
            .I(N__7448));
    InMux I__1494 (
            .O(N__7463),
            .I(N__7445));
    InMux I__1493 (
            .O(N__7462),
            .I(N__7440));
    InMux I__1492 (
            .O(N__7459),
            .I(N__7440));
    LocalMux I__1491 (
            .O(N__7456),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    Odrv4 I__1490 (
            .O(N__7453),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1489 (
            .O(N__7448),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1488 (
            .O(N__7445),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1487 (
            .O(N__7440),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    CascadeMux I__1486 (
            .O(N__7429),
            .I(N__7424));
    InMux I__1485 (
            .O(N__7428),
            .I(N__7421));
    InMux I__1484 (
            .O(N__7427),
            .I(N__7418));
    InMux I__1483 (
            .O(N__7424),
            .I(N__7415));
    LocalMux I__1482 (
            .O(N__7421),
            .I(N__7412));
    LocalMux I__1481 (
            .O(N__7418),
            .I(\U712_REG_SM.N_209 ));
    LocalMux I__1480 (
            .O(N__7415),
            .I(\U712_REG_SM.N_209 ));
    Odrv4 I__1479 (
            .O(N__7412),
            .I(\U712_REG_SM.N_209 ));
    CascadeMux I__1478 (
            .O(N__7405),
            .I(N__7402));
    InMux I__1477 (
            .O(N__7402),
            .I(N__7397));
    InMux I__1476 (
            .O(N__7401),
            .I(N__7394));
    InMux I__1475 (
            .O(N__7400),
            .I(N__7391));
    LocalMux I__1474 (
            .O(N__7397),
            .I(\U712_REG_SM.N_229 ));
    LocalMux I__1473 (
            .O(N__7394),
            .I(\U712_REG_SM.N_229 ));
    LocalMux I__1472 (
            .O(N__7391),
            .I(\U712_REG_SM.N_229 ));
    CascadeMux I__1471 (
            .O(N__7384),
            .I(N__7378));
    CascadeMux I__1470 (
            .O(N__7383),
            .I(N__7373));
    InMux I__1469 (
            .O(N__7382),
            .I(N__7369));
    InMux I__1468 (
            .O(N__7381),
            .I(N__7366));
    InMux I__1467 (
            .O(N__7378),
            .I(N__7363));
    InMux I__1466 (
            .O(N__7377),
            .I(N__7360));
    InMux I__1465 (
            .O(N__7376),
            .I(N__7355));
    InMux I__1464 (
            .O(N__7373),
            .I(N__7355));
    InMux I__1463 (
            .O(N__7372),
            .I(N__7352));
    LocalMux I__1462 (
            .O(N__7369),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1461 (
            .O(N__7366),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1460 (
            .O(N__7363),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1459 (
            .O(N__7360),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1458 (
            .O(N__7355),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1457 (
            .O(N__7352),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    InMux I__1456 (
            .O(N__7339),
            .I(N__7336));
    LocalMux I__1455 (
            .O(N__7336),
            .I(N__7331));
    InMux I__1454 (
            .O(N__7335),
            .I(N__7328));
    InMux I__1453 (
            .O(N__7334),
            .I(N__7325));
    Odrv4 I__1452 (
            .O(N__7331),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1451 (
            .O(N__7328),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1450 (
            .O(N__7325),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    IoInMux I__1449 (
            .O(N__7318),
            .I(N__7315));
    LocalMux I__1448 (
            .O(N__7315),
            .I(N__7312));
    Span4Mux_s1_h I__1447 (
            .O(N__7312),
            .I(N__7309));
    Sp12to4 I__1446 (
            .O(N__7309),
            .I(N__7306));
    Span12Mux_v I__1445 (
            .O(N__7306),
            .I(N__7303));
    Span12Mux_h I__1444 (
            .O(N__7303),
            .I(N__7300));
    Odrv12 I__1443 (
            .O(N__7300),
            .I(N_858_i));
    CascadeMux I__1442 (
            .O(N__7297),
            .I(N__7294));
    InMux I__1441 (
            .O(N__7294),
            .I(N__7285));
    InMux I__1440 (
            .O(N__7293),
            .I(N__7282));
    InMux I__1439 (
            .O(N__7292),
            .I(N__7277));
    InMux I__1438 (
            .O(N__7291),
            .I(N__7277));
    InMux I__1437 (
            .O(N__7290),
            .I(N__7272));
    InMux I__1436 (
            .O(N__7289),
            .I(N__7272));
    InMux I__1435 (
            .O(N__7288),
            .I(N__7269));
    LocalMux I__1434 (
            .O(N__7285),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1433 (
            .O(N__7282),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1432 (
            .O(N__7277),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1431 (
            .O(N__7272),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1430 (
            .O(N__7269),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__1429 (
            .O(N__7258),
            .I(N__7255));
    InMux I__1428 (
            .O(N__7255),
            .I(N__7247));
    InMux I__1427 (
            .O(N__7254),
            .I(N__7242));
    InMux I__1426 (
            .O(N__7253),
            .I(N__7242));
    InMux I__1425 (
            .O(N__7252),
            .I(N__7237));
    InMux I__1424 (
            .O(N__7251),
            .I(N__7237));
    InMux I__1423 (
            .O(N__7250),
            .I(N__7234));
    LocalMux I__1422 (
            .O(N__7247),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1421 (
            .O(N__7242),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1420 (
            .O(N__7237),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1419 (
            .O(N__7234),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1418 (
            .O(N__7225),
            .I(N__7220));
    CascadeMux I__1417 (
            .O(N__7224),
            .I(N__7213));
    InMux I__1416 (
            .O(N__7223),
            .I(N__7210));
    InMux I__1415 (
            .O(N__7220),
            .I(N__7207));
    InMux I__1414 (
            .O(N__7219),
            .I(N__7204));
    InMux I__1413 (
            .O(N__7218),
            .I(N__7197));
    InMux I__1412 (
            .O(N__7217),
            .I(N__7197));
    InMux I__1411 (
            .O(N__7216),
            .I(N__7197));
    InMux I__1410 (
            .O(N__7213),
            .I(N__7194));
    LocalMux I__1409 (
            .O(N__7210),
            .I(N__7191));
    LocalMux I__1408 (
            .O(N__7207),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1407 (
            .O(N__7204),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1406 (
            .O(N__7197),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1405 (
            .O(N__7194),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    Odrv4 I__1404 (
            .O(N__7191),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    InMux I__1403 (
            .O(N__7180),
            .I(N__7177));
    LocalMux I__1402 (
            .O(N__7177),
            .I(N__7172));
    InMux I__1401 (
            .O(N__7176),
            .I(N__7169));
    InMux I__1400 (
            .O(N__7175),
            .I(N__7166));
    Odrv4 I__1399 (
            .O(N__7172),
            .I(\U712_REG_SM.REG_TACK_0_sqmuxa ));
    LocalMux I__1398 (
            .O(N__7169),
            .I(\U712_REG_SM.REG_TACK_0_sqmuxa ));
    LocalMux I__1397 (
            .O(N__7166),
            .I(\U712_REG_SM.REG_TACK_0_sqmuxa ));
    CascadeMux I__1396 (
            .O(N__7159),
            .I(\U712_BYTE_ENABLE.N_319_cascade_ ));
    IoInMux I__1395 (
            .O(N__7156),
            .I(N__7153));
    LocalMux I__1394 (
            .O(N__7153),
            .I(N__7150));
    IoSpan4Mux I__1393 (
            .O(N__7150),
            .I(N__7147));
    Span4Mux_s2_h I__1392 (
            .O(N__7147),
            .I(N__7144));
    Span4Mux_h I__1391 (
            .O(N__7144),
            .I(N__7141));
    Sp12to4 I__1390 (
            .O(N__7141),
            .I(N__7138));
    Span12Mux_h I__1389 (
            .O(N__7138),
            .I(N__7135));
    Span12Mux_v I__1388 (
            .O(N__7135),
            .I(N__7132));
    Odrv12 I__1387 (
            .O(N__7132),
            .I(N_58_i));
    InMux I__1386 (
            .O(N__7129),
            .I(N__7126));
    LocalMux I__1385 (
            .O(N__7126),
            .I(\U712_BYTE_ENABLE.N_320 ));
    IoInMux I__1384 (
            .O(N__7123),
            .I(N__7120));
    LocalMux I__1383 (
            .O(N__7120),
            .I(N__7117));
    Span4Mux_s3_h I__1382 (
            .O(N__7117),
            .I(N__7114));
    Span4Mux_v I__1381 (
            .O(N__7114),
            .I(N__7111));
    Sp12to4 I__1380 (
            .O(N__7111),
            .I(N__7108));
    Span12Mux_h I__1379 (
            .O(N__7108),
            .I(N__7105));
    Span12Mux_v I__1378 (
            .O(N__7105),
            .I(N__7102));
    Odrv12 I__1377 (
            .O(N__7102),
            .I(N_56_i));
    InMux I__1376 (
            .O(N__7099),
            .I(N__7093));
    InMux I__1375 (
            .O(N__7098),
            .I(N__7093));
    LocalMux I__1374 (
            .O(N__7093),
            .I(\U712_BYTE_ENABLE.N_318 ));
    CascadeMux I__1373 (
            .O(N__7090),
            .I(\U712_BYTE_ENABLE.N_323_cascade_ ));
    InMux I__1372 (
            .O(N__7087),
            .I(N__7081));
    InMux I__1371 (
            .O(N__7086),
            .I(N__7081));
    LocalMux I__1370 (
            .O(N__7081),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ));
    IoInMux I__1369 (
            .O(N__7078),
            .I(N__7075));
    LocalMux I__1368 (
            .O(N__7075),
            .I(N__7072));
    Span4Mux_s1_v I__1367 (
            .O(N__7072),
            .I(N__7069));
    Span4Mux_v I__1366 (
            .O(N__7069),
            .I(N__7066));
    Span4Mux_v I__1365 (
            .O(N__7066),
            .I(N__7063));
    Span4Mux_v I__1364 (
            .O(N__7063),
            .I(N__7060));
    Span4Mux_v I__1363 (
            .O(N__7060),
            .I(N__7057));
    Odrv4 I__1362 (
            .O(N__7057),
            .I(N_54_i));
    IoInMux I__1361 (
            .O(N__7054),
            .I(N__7051));
    LocalMux I__1360 (
            .O(N__7051),
            .I(N__7047));
    CascadeMux I__1359 (
            .O(N__7050),
            .I(N__7041));
    IoSpan4Mux I__1358 (
            .O(N__7047),
            .I(N__7038));
    InMux I__1357 (
            .O(N__7046),
            .I(N__7029));
    InMux I__1356 (
            .O(N__7045),
            .I(N__7029));
    InMux I__1355 (
            .O(N__7044),
            .I(N__7029));
    InMux I__1354 (
            .O(N__7041),
            .I(N__7029));
    Sp12to4 I__1353 (
            .O(N__7038),
            .I(N__7026));
    LocalMux I__1352 (
            .O(N__7029),
            .I(N__7023));
    Span12Mux_s7_v I__1351 (
            .O(N__7026),
            .I(N__7019));
    Span4Mux_h I__1350 (
            .O(N__7023),
            .I(N__7016));
    InMux I__1349 (
            .O(N__7022),
            .I(N__7013));
    Odrv12 I__1348 (
            .O(N__7019),
            .I(DBENn_c));
    Odrv4 I__1347 (
            .O(N__7016),
            .I(DBENn_c));
    LocalMux I__1346 (
            .O(N__7013),
            .I(DBENn_c));
    InMux I__1345 (
            .O(N__7006),
            .I(N__6997));
    InMux I__1344 (
            .O(N__7005),
            .I(N__6997));
    InMux I__1343 (
            .O(N__7004),
            .I(N__6992));
    InMux I__1342 (
            .O(N__7003),
            .I(N__6992));
    InMux I__1341 (
            .O(N__7002),
            .I(N__6989));
    LocalMux I__1340 (
            .O(N__6997),
            .I(N__6982));
    LocalMux I__1339 (
            .O(N__6992),
            .I(N__6982));
    LocalMux I__1338 (
            .O(N__6989),
            .I(N__6978));
    InMux I__1337 (
            .O(N__6988),
            .I(N__6975));
    CascadeMux I__1336 (
            .O(N__6987),
            .I(N__6972));
    Span4Mux_h I__1335 (
            .O(N__6982),
            .I(N__6967));
    InMux I__1334 (
            .O(N__6981),
            .I(N__6964));
    Span4Mux_v I__1333 (
            .O(N__6978),
            .I(N__6961));
    LocalMux I__1332 (
            .O(N__6975),
            .I(N__6958));
    InMux I__1331 (
            .O(N__6972),
            .I(N__6951));
    InMux I__1330 (
            .O(N__6971),
            .I(N__6951));
    InMux I__1329 (
            .O(N__6970),
            .I(N__6951));
    Odrv4 I__1328 (
            .O(N__6967),
            .I(DMA_CYCLE));
    LocalMux I__1327 (
            .O(N__6964),
            .I(DMA_CYCLE));
    Odrv4 I__1326 (
            .O(N__6961),
            .I(DMA_CYCLE));
    Odrv4 I__1325 (
            .O(N__6958),
            .I(DMA_CYCLE));
    LocalMux I__1324 (
            .O(N__6951),
            .I(DMA_CYCLE));
    CascadeMux I__1323 (
            .O(N__6940),
            .I(\U712_BYTE_ENABLE.N_315_cascade_ ));
    IoInMux I__1322 (
            .O(N__6937),
            .I(N__6934));
    LocalMux I__1321 (
            .O(N__6934),
            .I(N__6931));
    IoSpan4Mux I__1320 (
            .O(N__6931),
            .I(N__6928));
    Sp12to4 I__1319 (
            .O(N__6928),
            .I(N__6925));
    Span12Mux_s9_h I__1318 (
            .O(N__6925),
            .I(N__6922));
    Span12Mux_v I__1317 (
            .O(N__6922),
            .I(N__6919));
    Odrv12 I__1316 (
            .O(N__6919),
            .I(N_60_i));
    CascadeMux I__1315 (
            .O(N__6916),
            .I(N__6913));
    InMux I__1314 (
            .O(N__6913),
            .I(N__6910));
    LocalMux I__1313 (
            .O(N__6910),
            .I(N__6907));
    Span12Mux_h I__1312 (
            .O(N__6907),
            .I(N__6904));
    Odrv12 I__1311 (
            .O(N__6904),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__1310 (
            .O(N__6901),
            .I(N__6894));
    InMux I__1309 (
            .O(N__6900),
            .I(N__6894));
    InMux I__1308 (
            .O(N__6899),
            .I(N__6891));
    LocalMux I__1307 (
            .O(N__6894),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    LocalMux I__1306 (
            .O(N__6891),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    InMux I__1305 (
            .O(N__6886),
            .I(N__6883));
    LocalMux I__1304 (
            .O(N__6883),
            .I(N__6878));
    InMux I__1303 (
            .O(N__6882),
            .I(N__6875));
    InMux I__1302 (
            .O(N__6881),
            .I(N__6872));
    Span4Mux_h I__1301 (
            .O(N__6878),
            .I(N__6869));
    LocalMux I__1300 (
            .O(N__6875),
            .I(\U712_CHIP_RAM.N_348 ));
    LocalMux I__1299 (
            .O(N__6872),
            .I(\U712_CHIP_RAM.N_348 ));
    Odrv4 I__1298 (
            .O(N__6869),
            .I(\U712_CHIP_RAM.N_348 ));
    InMux I__1297 (
            .O(N__6862),
            .I(N__6858));
    InMux I__1296 (
            .O(N__6861),
            .I(N__6855));
    LocalMux I__1295 (
            .O(N__6858),
            .I(N__6852));
    LocalMux I__1294 (
            .O(N__6855),
            .I(\U712_CHIP_RAM.N_186 ));
    Odrv4 I__1293 (
            .O(N__6852),
            .I(\U712_CHIP_RAM.N_186 ));
    CascadeMux I__1292 (
            .O(N__6847),
            .I(N__6844));
    InMux I__1291 (
            .O(N__6844),
            .I(N__6838));
    CascadeMux I__1290 (
            .O(N__6843),
            .I(N__6832));
    InMux I__1289 (
            .O(N__6842),
            .I(N__6829));
    InMux I__1288 (
            .O(N__6841),
            .I(N__6826));
    LocalMux I__1287 (
            .O(N__6838),
            .I(N__6823));
    InMux I__1286 (
            .O(N__6837),
            .I(N__6820));
    CascadeMux I__1285 (
            .O(N__6836),
            .I(N__6817));
    InMux I__1284 (
            .O(N__6835),
            .I(N__6809));
    InMux I__1283 (
            .O(N__6832),
            .I(N__6809));
    LocalMux I__1282 (
            .O(N__6829),
            .I(N__6806));
    LocalMux I__1281 (
            .O(N__6826),
            .I(N__6803));
    Span4Mux_v I__1280 (
            .O(N__6823),
            .I(N__6798));
    LocalMux I__1279 (
            .O(N__6820),
            .I(N__6798));
    InMux I__1278 (
            .O(N__6817),
            .I(N__6791));
    InMux I__1277 (
            .O(N__6816),
            .I(N__6791));
    InMux I__1276 (
            .O(N__6815),
            .I(N__6791));
    InMux I__1275 (
            .O(N__6814),
            .I(N__6788));
    LocalMux I__1274 (
            .O(N__6809),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1273 (
            .O(N__6806),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1272 (
            .O(N__6803),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1271 (
            .O(N__6798),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1270 (
            .O(N__6791),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1269 (
            .O(N__6788),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    InMux I__1268 (
            .O(N__6775),
            .I(N__6770));
    InMux I__1267 (
            .O(N__6774),
            .I(N__6767));
    InMux I__1266 (
            .O(N__6773),
            .I(N__6762));
    LocalMux I__1265 (
            .O(N__6770),
            .I(N__6757));
    LocalMux I__1264 (
            .O(N__6767),
            .I(N__6757));
    InMux I__1263 (
            .O(N__6766),
            .I(N__6754));
    InMux I__1262 (
            .O(N__6765),
            .I(N__6751));
    LocalMux I__1261 (
            .O(N__6762),
            .I(N__6748));
    Span4Mux_h I__1260 (
            .O(N__6757),
            .I(N__6745));
    LocalMux I__1259 (
            .O(N__6754),
            .I(\U712_CHIP_RAM.N_198 ));
    LocalMux I__1258 (
            .O(N__6751),
            .I(\U712_CHIP_RAM.N_198 ));
    Odrv4 I__1257 (
            .O(N__6748),
            .I(\U712_CHIP_RAM.N_198 ));
    Odrv4 I__1256 (
            .O(N__6745),
            .I(\U712_CHIP_RAM.N_198 ));
    InMux I__1255 (
            .O(N__6736),
            .I(N__6731));
    InMux I__1254 (
            .O(N__6735),
            .I(N__6725));
    InMux I__1253 (
            .O(N__6734),
            .I(N__6725));
    LocalMux I__1252 (
            .O(N__6731),
            .I(N__6722));
    InMux I__1251 (
            .O(N__6730),
            .I(N__6719));
    LocalMux I__1250 (
            .O(N__6725),
            .I(N__6716));
    Span4Mux_h I__1249 (
            .O(N__6722),
            .I(N__6713));
    LocalMux I__1248 (
            .O(N__6719),
            .I(N__6710));
    Span4Mux_h I__1247 (
            .O(N__6716),
            .I(N__6707));
    Odrv4 I__1246 (
            .O(N__6713),
            .I(\U712_CHIP_RAM.N_389 ));
    Odrv4 I__1245 (
            .O(N__6710),
            .I(\U712_CHIP_RAM.N_389 ));
    Odrv4 I__1244 (
            .O(N__6707),
            .I(\U712_CHIP_RAM.N_389 ));
    CascadeMux I__1243 (
            .O(N__6700),
            .I(\U712_CHIP_RAM.N_313_cascade_ ));
    InMux I__1242 (
            .O(N__6697),
            .I(N__6694));
    LocalMux I__1241 (
            .O(N__6694),
            .I(\U712_CHIP_RAM.N_314 ));
    CascadeMux I__1240 (
            .O(N__6691),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ));
    CEMux I__1239 (
            .O(N__6688),
            .I(N__6685));
    LocalMux I__1238 (
            .O(N__6685),
            .I(N__6682));
    Span4Mux_h I__1237 (
            .O(N__6682),
            .I(N__6679));
    Span4Mux_h I__1236 (
            .O(N__6679),
            .I(N__6676));
    Odrv4 I__1235 (
            .O(N__6676),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ));
    InMux I__1234 (
            .O(N__6673),
            .I(N__6669));
    InMux I__1233 (
            .O(N__6672),
            .I(N__6666));
    LocalMux I__1232 (
            .O(N__6669),
            .I(N__6663));
    LocalMux I__1231 (
            .O(N__6666),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    Odrv4 I__1230 (
            .O(N__6663),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1229 (
            .O(N__6658),
            .I(N__6654));
    InMux I__1228 (
            .O(N__6657),
            .I(N__6651));
    LocalMux I__1227 (
            .O(N__6654),
            .I(N__6648));
    LocalMux I__1226 (
            .O(N__6651),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv4 I__1225 (
            .O(N__6648),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__1224 (
            .O(N__6643),
            .I(N__6640));
    InMux I__1223 (
            .O(N__6640),
            .I(N__6637));
    LocalMux I__1222 (
            .O(N__6637),
            .I(N__6633));
    InMux I__1221 (
            .O(N__6636),
            .I(N__6630));
    Odrv4 I__1220 (
            .O(N__6633),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1219 (
            .O(N__6630),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1218 (
            .O(N__6625),
            .I(N__6622));
    LocalMux I__1217 (
            .O(N__6622),
            .I(N__6619));
    Odrv4 I__1216 (
            .O(N__6619),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__1215 (
            .O(N__6616),
            .I(N__6610));
    InMux I__1214 (
            .O(N__6615),
            .I(N__6607));
    InMux I__1213 (
            .O(N__6614),
            .I(N__6604));
    InMux I__1212 (
            .O(N__6613),
            .I(N__6601));
    InMux I__1211 (
            .O(N__6610),
            .I(N__6598));
    LocalMux I__1210 (
            .O(N__6607),
            .I(N__6595));
    LocalMux I__1209 (
            .O(N__6604),
            .I(N__6589));
    LocalMux I__1208 (
            .O(N__6601),
            .I(N__6589));
    LocalMux I__1207 (
            .O(N__6598),
            .I(N__6583));
    Span4Mux_v I__1206 (
            .O(N__6595),
            .I(N__6583));
    InMux I__1205 (
            .O(N__6594),
            .I(N__6580));
    Span4Mux_h I__1204 (
            .O(N__6589),
            .I(N__6577));
    InMux I__1203 (
            .O(N__6588),
            .I(N__6574));
    Odrv4 I__1202 (
            .O(N__6583),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1201 (
            .O(N__6580),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1200 (
            .O(N__6577),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1199 (
            .O(N__6574),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1198 (
            .O(N__6565),
            .I(N__6562));
    LocalMux I__1197 (
            .O(N__6562),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ));
    CascadeMux I__1196 (
            .O(N__6559),
            .I(N__6556));
    InMux I__1195 (
            .O(N__6556),
            .I(N__6553));
    LocalMux I__1194 (
            .O(N__6553),
            .I(N__6549));
    CascadeMux I__1193 (
            .O(N__6552),
            .I(N__6545));
    Span4Mux_h I__1192 (
            .O(N__6549),
            .I(N__6538));
    InMux I__1191 (
            .O(N__6548),
            .I(N__6535));
    InMux I__1190 (
            .O(N__6545),
            .I(N__6530));
    InMux I__1189 (
            .O(N__6544),
            .I(N__6530));
    InMux I__1188 (
            .O(N__6543),
            .I(N__6525));
    InMux I__1187 (
            .O(N__6542),
            .I(N__6525));
    InMux I__1186 (
            .O(N__6541),
            .I(N__6522));
    Odrv4 I__1185 (
            .O(N__6538),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1184 (
            .O(N__6535),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1183 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1182 (
            .O(N__6525),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1181 (
            .O(N__6522),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1180 (
            .O(N__6511),
            .I(N__6508));
    LocalMux I__1179 (
            .O(N__6508),
            .I(N__6505));
    Span4Mux_v I__1178 (
            .O(N__6505),
            .I(N__6501));
    InMux I__1177 (
            .O(N__6504),
            .I(N__6498));
    Odrv4 I__1176 (
            .O(N__6501),
            .I(LATCH_RAM));
    LocalMux I__1175 (
            .O(N__6498),
            .I(LATCH_RAM));
    InMux I__1174 (
            .O(N__6493),
            .I(N__6488));
    InMux I__1173 (
            .O(N__6492),
            .I(N__6484));
    InMux I__1172 (
            .O(N__6491),
            .I(N__6481));
    LocalMux I__1171 (
            .O(N__6488),
            .I(N__6478));
    CascadeMux I__1170 (
            .O(N__6487),
            .I(N__6475));
    LocalMux I__1169 (
            .O(N__6484),
            .I(N__6468));
    LocalMux I__1168 (
            .O(N__6481),
            .I(N__6468));
    Span4Mux_h I__1167 (
            .O(N__6478),
            .I(N__6468));
    InMux I__1166 (
            .O(N__6475),
            .I(N__6465));
    Odrv4 I__1165 (
            .O(N__6468),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1164 (
            .O(N__6465),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1163 (
            .O(N__6460),
            .I(N__6457));
    LocalMux I__1162 (
            .O(N__6457),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__1161 (
            .O(N__6454),
            .I(N__6450));
    InMux I__1160 (
            .O(N__6453),
            .I(N__6447));
    InMux I__1159 (
            .O(N__6450),
            .I(N__6444));
    LocalMux I__1158 (
            .O(N__6447),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1157 (
            .O(N__6444),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1156 (
            .O(N__6439),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1155 (
            .O(N__6436),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1154 (
            .O(N__6433),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1153 (
            .O(N__6430),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__1152 (
            .O(N__6427),
            .I(N__6409));
    ClkMux I__1151 (
            .O(N__6426),
            .I(N__6409));
    ClkMux I__1150 (
            .O(N__6425),
            .I(N__6409));
    ClkMux I__1149 (
            .O(N__6424),
            .I(N__6409));
    ClkMux I__1148 (
            .O(N__6423),
            .I(N__6409));
    ClkMux I__1147 (
            .O(N__6422),
            .I(N__6409));
    GlobalMux I__1146 (
            .O(N__6409),
            .I(N__6406));
    gio2CtrlBuf I__1145 (
            .O(N__6406),
            .I(C1_c_g));
    SRMux I__1144 (
            .O(N__6403),
            .I(N__6400));
    LocalMux I__1143 (
            .O(N__6400),
            .I(N__6397));
    Span4Mux_h I__1142 (
            .O(N__6397),
            .I(N__6394));
    Odrv4 I__1141 (
            .O(N__6394),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    IoInMux I__1140 (
            .O(N__6391),
            .I(N__6388));
    LocalMux I__1139 (
            .O(N__6388),
            .I(N__6385));
    Span4Mux_s2_v I__1138 (
            .O(N__6385),
            .I(N__6382));
    Sp12to4 I__1137 (
            .O(N__6382),
            .I(N__6379));
    Span12Mux_h I__1136 (
            .O(N__6379),
            .I(N__6376));
    Odrv12 I__1135 (
            .O(N__6376),
            .I(BANK0_c));
    InMux I__1134 (
            .O(N__6373),
            .I(N__6370));
    LocalMux I__1133 (
            .O(N__6370),
            .I(N__6367));
    Span12Mux_v I__1132 (
            .O(N__6367),
            .I(N__6364));
    Span12Mux_h I__1131 (
            .O(N__6364),
            .I(N__6361));
    Odrv12 I__1130 (
            .O(N__6361),
            .I(A_c_20));
    InMux I__1129 (
            .O(N__6358),
            .I(N__6355));
    LocalMux I__1128 (
            .O(N__6355),
            .I(\U712_CHIP_RAM.N_307 ));
    CascadeMux I__1127 (
            .O(N__6352),
            .I(N__6348));
    CascadeMux I__1126 (
            .O(N__6351),
            .I(N__6345));
    InMux I__1125 (
            .O(N__6348),
            .I(N__6342));
    InMux I__1124 (
            .O(N__6345),
            .I(N__6338));
    LocalMux I__1123 (
            .O(N__6342),
            .I(N__6334));
    InMux I__1122 (
            .O(N__6341),
            .I(N__6331));
    LocalMux I__1121 (
            .O(N__6338),
            .I(N__6328));
    InMux I__1120 (
            .O(N__6337),
            .I(N__6324));
    Sp12to4 I__1119 (
            .O(N__6334),
            .I(N__6321));
    LocalMux I__1118 (
            .O(N__6331),
            .I(N__6316));
    Span4Mux_h I__1117 (
            .O(N__6328),
            .I(N__6316));
    InMux I__1116 (
            .O(N__6327),
            .I(N__6313));
    LocalMux I__1115 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv12 I__1114 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__1113 (
            .O(N__6316),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1112 (
            .O(N__6313),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__1111 (
            .O(N__6304),
            .I(N__6301));
    LocalMux I__1110 (
            .O(N__6301),
            .I(\U712_CHIP_RAM.N_405 ));
    InMux I__1109 (
            .O(N__6298),
            .I(N__6287));
    InMux I__1108 (
            .O(N__6297),
            .I(N__6287));
    InMux I__1107 (
            .O(N__6296),
            .I(N__6287));
    InMux I__1106 (
            .O(N__6295),
            .I(N__6281));
    InMux I__1105 (
            .O(N__6294),
            .I(N__6278));
    LocalMux I__1104 (
            .O(N__6287),
            .I(N__6275));
    InMux I__1103 (
            .O(N__6286),
            .I(N__6271));
    InMux I__1102 (
            .O(N__6285),
            .I(N__6265));
    InMux I__1101 (
            .O(N__6284),
            .I(N__6265));
    LocalMux I__1100 (
            .O(N__6281),
            .I(N__6262));
    LocalMux I__1099 (
            .O(N__6278),
            .I(N__6259));
    Span4Mux_h I__1098 (
            .O(N__6275),
            .I(N__6256));
    InMux I__1097 (
            .O(N__6274),
            .I(N__6253));
    LocalMux I__1096 (
            .O(N__6271),
            .I(N__6250));
    InMux I__1095 (
            .O(N__6270),
            .I(N__6247));
    LocalMux I__1094 (
            .O(N__6265),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1093 (
            .O(N__6262),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1092 (
            .O(N__6259),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1091 (
            .O(N__6256),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1090 (
            .O(N__6253),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv12 I__1089 (
            .O(N__6250),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1088 (
            .O(N__6247),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1087 (
            .O(N__6232),
            .I(\U712_CHIP_RAM.N_405_cascade_ ));
    CascadeMux I__1086 (
            .O(N__6229),
            .I(N__6225));
    InMux I__1085 (
            .O(N__6228),
            .I(N__6221));
    InMux I__1084 (
            .O(N__6225),
            .I(N__6218));
    CascadeMux I__1083 (
            .O(N__6224),
            .I(N__6211));
    LocalMux I__1082 (
            .O(N__6221),
            .I(N__6207));
    LocalMux I__1081 (
            .O(N__6218),
            .I(N__6204));
    InMux I__1080 (
            .O(N__6217),
            .I(N__6201));
    InMux I__1079 (
            .O(N__6216),
            .I(N__6198));
    InMux I__1078 (
            .O(N__6215),
            .I(N__6194));
    InMux I__1077 (
            .O(N__6214),
            .I(N__6191));
    InMux I__1076 (
            .O(N__6211),
            .I(N__6188));
    CascadeMux I__1075 (
            .O(N__6210),
            .I(N__6185));
    Span4Mux_v I__1074 (
            .O(N__6207),
            .I(N__6178));
    Span4Mux_h I__1073 (
            .O(N__6204),
            .I(N__6173));
    LocalMux I__1072 (
            .O(N__6201),
            .I(N__6173));
    LocalMux I__1071 (
            .O(N__6198),
            .I(N__6170));
    InMux I__1070 (
            .O(N__6197),
            .I(N__6167));
    LocalMux I__1069 (
            .O(N__6194),
            .I(N__6160));
    LocalMux I__1068 (
            .O(N__6191),
            .I(N__6160));
    LocalMux I__1067 (
            .O(N__6188),
            .I(N__6160));
    InMux I__1066 (
            .O(N__6185),
            .I(N__6155));
    InMux I__1065 (
            .O(N__6184),
            .I(N__6155));
    InMux I__1064 (
            .O(N__6183),
            .I(N__6148));
    InMux I__1063 (
            .O(N__6182),
            .I(N__6148));
    InMux I__1062 (
            .O(N__6181),
            .I(N__6148));
    Odrv4 I__1061 (
            .O(N__6178),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1060 (
            .O(N__6173),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1059 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1058 (
            .O(N__6167),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1057 (
            .O(N__6160),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1056 (
            .O(N__6155),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1055 (
            .O(N__6148),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1054 (
            .O(N__6133),
            .I(\U712_CHIP_RAM.N_303_cascade_ ));
    CEMux I__1053 (
            .O(N__6130),
            .I(N__6127));
    LocalMux I__1052 (
            .O(N__6127),
            .I(N__6124));
    Span4Mux_v I__1051 (
            .O(N__6124),
            .I(N__6121));
    Span4Mux_h I__1050 (
            .O(N__6121),
            .I(N__6118));
    Odrv4 I__1049 (
            .O(N__6118),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ));
    CascadeMux I__1048 (
            .O(N__6115),
            .I(N__6112));
    InMux I__1047 (
            .O(N__6112),
            .I(N__6109));
    LocalMux I__1046 (
            .O(N__6109),
            .I(\U712_CHIP_RAM.N_136 ));
    InMux I__1045 (
            .O(N__6106),
            .I(N__6100));
    InMux I__1044 (
            .O(N__6105),
            .I(N__6100));
    LocalMux I__1043 (
            .O(N__6100),
            .I(N__6097));
    Span12Mux_v I__1042 (
            .O(N__6097),
            .I(N__6094));
    Span12Mux_h I__1041 (
            .O(N__6094),
            .I(N__6091));
    Odrv12 I__1040 (
            .O(N__6091),
            .I(A_c_10));
    InMux I__1039 (
            .O(N__6088),
            .I(N__6085));
    LocalMux I__1038 (
            .O(N__6085),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1037 (
            .O(N__6082),
            .I(bfn_10_8_0_));
    InMux I__1036 (
            .O(N__6079),
            .I(N__6075));
    InMux I__1035 (
            .O(N__6078),
            .I(N__6072));
    LocalMux I__1034 (
            .O(N__6075),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__1033 (
            .O(N__6072),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1032 (
            .O(N__6067),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1031 (
            .O(N__6064),
            .I(N__6060));
    InMux I__1030 (
            .O(N__6063),
            .I(N__6057));
    LocalMux I__1029 (
            .O(N__6060),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__1028 (
            .O(N__6057),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__1027 (
            .O(N__6052),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1026 (
            .O(N__6049),
            .I(N__6045));
    InMux I__1025 (
            .O(N__6048),
            .I(N__6042));
    LocalMux I__1024 (
            .O(N__6045),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1023 (
            .O(N__6042),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1022 (
            .O(N__6037),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1021 (
            .O(N__6034),
            .I(\U712_REG_SM.N_209_cascade_ ));
    InMux I__1020 (
            .O(N__6031),
            .I(N__6028));
    LocalMux I__1019 (
            .O(N__6028),
            .I(N__6025));
    Odrv4 I__1018 (
            .O(N__6025),
            .I(\U712_REG_SM.LDSn_7_iv_i_0 ));
    CascadeMux I__1017 (
            .O(N__6022),
            .I(\U712_REG_SM.N_297_cascade_ ));
    IoInMux I__1016 (
            .O(N__6019),
            .I(N__6016));
    LocalMux I__1015 (
            .O(N__6016),
            .I(N__6013));
    Span12Mux_s11_v I__1014 (
            .O(N__6013),
            .I(N__6010));
    Span12Mux_h I__1013 (
            .O(N__6010),
            .I(N__6005));
    InMux I__1012 (
            .O(N__6009),
            .I(N__6000));
    InMux I__1011 (
            .O(N__6008),
            .I(N__6000));
    Odrv12 I__1010 (
            .O(N__6005),
            .I(LDSn_c));
    LocalMux I__1009 (
            .O(N__6000),
            .I(LDSn_c));
    CascadeMux I__1008 (
            .O(N__5995),
            .I(\U712_REG_SM.N_295_cascade_ ));
    InMux I__1007 (
            .O(N__5992),
            .I(N__5986));
    InMux I__1006 (
            .O(N__5991),
            .I(N__5986));
    LocalMux I__1005 (
            .O(N__5986),
            .I(\U712_REG_SM.N_153 ));
    IoInMux I__1004 (
            .O(N__5983),
            .I(N__5980));
    LocalMux I__1003 (
            .O(N__5980),
            .I(N__5977));
    Span4Mux_s0_v I__1002 (
            .O(N__5977),
            .I(N__5974));
    Span4Mux_v I__1001 (
            .O(N__5974),
            .I(N__5971));
    Sp12to4 I__1000 (
            .O(N__5971),
            .I(N__5968));
    Span12Mux_h I__999 (
            .O(N__5968),
            .I(N__5963));
    InMux I__998 (
            .O(N__5967),
            .I(N__5958));
    InMux I__997 (
            .O(N__5966),
            .I(N__5958));
    Odrv12 I__996 (
            .O(N__5963),
            .I(UDSn_c));
    LocalMux I__995 (
            .O(N__5958),
            .I(UDSn_c));
    InMux I__994 (
            .O(N__5953),
            .I(N__5949));
    IoInMux I__993 (
            .O(N__5952),
            .I(N__5946));
    LocalMux I__992 (
            .O(N__5949),
            .I(N__5943));
    LocalMux I__991 (
            .O(N__5946),
            .I(N__5940));
    Span4Mux_v I__990 (
            .O(N__5943),
            .I(N__5937));
    IoSpan4Mux I__989 (
            .O(N__5940),
            .I(N__5934));
    Sp12to4 I__988 (
            .O(N__5937),
            .I(N__5931));
    IoSpan4Mux I__987 (
            .O(N__5934),
            .I(N__5928));
    Span12Mux_h I__986 (
            .O(N__5931),
            .I(N__5925));
    IoSpan4Mux I__985 (
            .O(N__5928),
            .I(N__5922));
    Odrv12 I__984 (
            .O(N__5925),
            .I(C1_c));
    Odrv4 I__983 (
            .O(N__5922),
            .I(C1_c));
    InMux I__982 (
            .O(N__5917),
            .I(N__5914));
    LocalMux I__981 (
            .O(N__5914),
            .I(N__5911));
    Odrv4 I__980 (
            .O(N__5911),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__979 (
            .O(N__5908),
            .I(N__5905));
    LocalMux I__978 (
            .O(N__5905),
            .I(N__5902));
    Span4Mux_v I__977 (
            .O(N__5902),
            .I(N__5899));
    Sp12to4 I__976 (
            .O(N__5899),
            .I(N__5896));
    Span12Mux_h I__975 (
            .O(N__5896),
            .I(N__5893));
    Span12Mux_v I__974 (
            .O(N__5893),
            .I(N__5890));
    Odrv12 I__973 (
            .O(N__5890),
            .I(REGSPACEn_c));
    InMux I__972 (
            .O(N__5887),
            .I(N__5884));
    LocalMux I__971 (
            .O(N__5884),
            .I(N__5880));
    InMux I__970 (
            .O(N__5883),
            .I(N__5877));
    Span4Mux_v I__969 (
            .O(N__5880),
            .I(N__5874));
    LocalMux I__968 (
            .O(N__5877),
            .I(\U712_REG_SM.CYCLE_RUNZ0 ));
    Odrv4 I__967 (
            .O(N__5874),
            .I(\U712_REG_SM.CYCLE_RUNZ0 ));
    CascadeMux I__966 (
            .O(N__5869),
            .I(N__5866));
    InMux I__965 (
            .O(N__5866),
            .I(N__5863));
    LocalMux I__964 (
            .O(N__5863),
            .I(N__5859));
    InMux I__963 (
            .O(N__5862),
            .I(N__5856));
    Span4Mux_v I__962 (
            .O(N__5859),
            .I(N__5853));
    LocalMux I__961 (
            .O(N__5856),
            .I(N__5850));
    Span4Mux_v I__960 (
            .O(N__5853),
            .I(N__5847));
    Span4Mux_v I__959 (
            .O(N__5850),
            .I(N__5844));
    Sp12to4 I__958 (
            .O(N__5847),
            .I(N__5839));
    Sp12to4 I__957 (
            .O(N__5844),
            .I(N__5839));
    Span12Mux_h I__956 (
            .O(N__5839),
            .I(N__5836));
    Odrv12 I__955 (
            .O(N__5836),
            .I(TSn_c));
    CascadeMux I__954 (
            .O(N__5833),
            .I(N__5829));
    InMux I__953 (
            .O(N__5832),
            .I(N__5825));
    InMux I__952 (
            .O(N__5829),
            .I(N__5822));
    InMux I__951 (
            .O(N__5828),
            .I(N__5819));
    LocalMux I__950 (
            .O(N__5825),
            .I(N__5816));
    LocalMux I__949 (
            .O(N__5822),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__948 (
            .O(N__5819),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv12 I__947 (
            .O(N__5816),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__946 (
            .O(N__5809),
            .I(N__5806));
    LocalMux I__945 (
            .O(N__5806),
            .I(N__5803));
    Odrv4 I__944 (
            .O(N__5803),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ));
    CascadeMux I__943 (
            .O(N__5800),
            .I(\U712_REG_SM.N_229_cascade_ ));
    InMux I__942 (
            .O(N__5797),
            .I(N__5788));
    InMux I__941 (
            .O(N__5796),
            .I(N__5788));
    InMux I__940 (
            .O(N__5795),
            .I(N__5783));
    InMux I__939 (
            .O(N__5794),
            .I(N__5783));
    InMux I__938 (
            .O(N__5793),
            .I(N__5780));
    LocalMux I__937 (
            .O(N__5788),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    LocalMux I__936 (
            .O(N__5783),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    LocalMux I__935 (
            .O(N__5780),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    InMux I__934 (
            .O(N__5773),
            .I(N__5768));
    InMux I__933 (
            .O(N__5772),
            .I(N__5765));
    InMux I__932 (
            .O(N__5771),
            .I(N__5762));
    LocalMux I__931 (
            .O(N__5768),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    LocalMux I__930 (
            .O(N__5765),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    LocalMux I__929 (
            .O(N__5762),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    CascadeMux I__928 (
            .O(N__5755),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_ ));
    InMux I__927 (
            .O(N__5752),
            .I(N__5749));
    LocalMux I__926 (
            .O(N__5749),
            .I(\U712_REG_SM.REG_CPU_CYCLE_e_1 ));
    InMux I__925 (
            .O(N__5746),
            .I(N__5743));
    LocalMux I__924 (
            .O(N__5743),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__923 (
            .O(N__5740),
            .I(N__5737));
    LocalMux I__922 (
            .O(N__5737),
            .I(\U712_REG_SM.N_224 ));
    CascadeMux I__921 (
            .O(N__5734),
            .I(\U712_REG_SM.N_224_cascade_ ));
    InMux I__920 (
            .O(N__5731),
            .I(N__5728));
    LocalMux I__919 (
            .O(N__5728),
            .I(\U712_CHIP_RAM.N_234 ));
    InMux I__918 (
            .O(N__5725),
            .I(N__5719));
    InMux I__917 (
            .O(N__5724),
            .I(N__5719));
    LocalMux I__916 (
            .O(N__5719),
            .I(N__5715));
    InMux I__915 (
            .O(N__5718),
            .I(N__5712));
    Odrv4 I__914 (
            .O(N__5715),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0 ));
    LocalMux I__913 (
            .O(N__5712),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0 ));
    InMux I__912 (
            .O(N__5707),
            .I(N__5702));
    InMux I__911 (
            .O(N__5706),
            .I(N__5698));
    InMux I__910 (
            .O(N__5705),
            .I(N__5695));
    LocalMux I__909 (
            .O(N__5702),
            .I(N__5692));
    InMux I__908 (
            .O(N__5701),
            .I(N__5688));
    LocalMux I__907 (
            .O(N__5698),
            .I(N__5684));
    LocalMux I__906 (
            .O(N__5695),
            .I(N__5681));
    Span4Mux_h I__905 (
            .O(N__5692),
            .I(N__5678));
    CascadeMux I__904 (
            .O(N__5691),
            .I(N__5675));
    LocalMux I__903 (
            .O(N__5688),
            .I(N__5671));
    InMux I__902 (
            .O(N__5687),
            .I(N__5668));
    Span4Mux_v I__901 (
            .O(N__5684),
            .I(N__5661));
    Span4Mux_v I__900 (
            .O(N__5681),
            .I(N__5661));
    Span4Mux_h I__899 (
            .O(N__5678),
            .I(N__5661));
    InMux I__898 (
            .O(N__5675),
            .I(N__5656));
    InMux I__897 (
            .O(N__5674),
            .I(N__5656));
    Odrv4 I__896 (
            .O(N__5671),
            .I(WRITE_CYCLE));
    LocalMux I__895 (
            .O(N__5668),
            .I(WRITE_CYCLE));
    Odrv4 I__894 (
            .O(N__5661),
            .I(WRITE_CYCLE));
    LocalMux I__893 (
            .O(N__5656),
            .I(WRITE_CYCLE));
    InMux I__892 (
            .O(N__5647),
            .I(N__5638));
    InMux I__891 (
            .O(N__5646),
            .I(N__5635));
    CascadeMux I__890 (
            .O(N__5645),
            .I(N__5632));
    CascadeMux I__889 (
            .O(N__5644),
            .I(N__5626));
    InMux I__888 (
            .O(N__5643),
            .I(N__5622));
    InMux I__887 (
            .O(N__5642),
            .I(N__5619));
    InMux I__886 (
            .O(N__5641),
            .I(N__5615));
    LocalMux I__885 (
            .O(N__5638),
            .I(N__5610));
    LocalMux I__884 (
            .O(N__5635),
            .I(N__5610));
    InMux I__883 (
            .O(N__5632),
            .I(N__5607));
    InMux I__882 (
            .O(N__5631),
            .I(N__5604));
    InMux I__881 (
            .O(N__5630),
            .I(N__5601));
    InMux I__880 (
            .O(N__5629),
            .I(N__5596));
    InMux I__879 (
            .O(N__5626),
            .I(N__5596));
    InMux I__878 (
            .O(N__5625),
            .I(N__5593));
    LocalMux I__877 (
            .O(N__5622),
            .I(N__5588));
    LocalMux I__876 (
            .O(N__5619),
            .I(N__5588));
    InMux I__875 (
            .O(N__5618),
            .I(N__5585));
    LocalMux I__874 (
            .O(N__5615),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__873 (
            .O(N__5610),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__872 (
            .O(N__5607),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__871 (
            .O(N__5604),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__870 (
            .O(N__5601),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__869 (
            .O(N__5596),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__868 (
            .O(N__5593),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__867 (
            .O(N__5588),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__866 (
            .O(N__5585),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__865 (
            .O(N__5566),
            .I(N__5563));
    LocalMux I__864 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ));
    CascadeMux I__863 (
            .O(N__5560),
            .I(N__5557));
    InMux I__862 (
            .O(N__5557),
            .I(N__5554));
    LocalMux I__861 (
            .O(N__5554),
            .I(\U712_CHIP_RAM.N_292 ));
    InMux I__860 (
            .O(N__5551),
            .I(N__5548));
    LocalMux I__859 (
            .O(N__5548),
            .I(N__5545));
    Odrv12 I__858 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.N_19 ));
    CascadeMux I__857 (
            .O(N__5542),
            .I(N__5539));
    InMux I__856 (
            .O(N__5539),
            .I(N__5536));
    LocalMux I__855 (
            .O(N__5536),
            .I(\U712_BYTE_ENABLE.N_185_i ));
    InMux I__854 (
            .O(N__5533),
            .I(N__5530));
    LocalMux I__853 (
            .O(N__5530),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_5 ));
    CascadeMux I__852 (
            .O(N__5527),
            .I(\U712_CHIP_RAM.N_391_cascade_ ));
    InMux I__851 (
            .O(N__5524),
            .I(N__5521));
    LocalMux I__850 (
            .O(N__5521),
            .I(\U712_CHIP_RAM.N_387 ));
    InMux I__849 (
            .O(N__5518),
            .I(N__5514));
    InMux I__848 (
            .O(N__5517),
            .I(N__5511));
    LocalMux I__847 (
            .O(N__5514),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ));
    LocalMux I__846 (
            .O(N__5511),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ));
    CascadeMux I__845 (
            .O(N__5506),
            .I(N__5502));
    InMux I__844 (
            .O(N__5505),
            .I(N__5496));
    InMux I__843 (
            .O(N__5502),
            .I(N__5493));
    InMux I__842 (
            .O(N__5501),
            .I(N__5488));
    InMux I__841 (
            .O(N__5500),
            .I(N__5488));
    InMux I__840 (
            .O(N__5499),
            .I(N__5484));
    LocalMux I__839 (
            .O(N__5496),
            .I(N__5480));
    LocalMux I__838 (
            .O(N__5493),
            .I(N__5475));
    LocalMux I__837 (
            .O(N__5488),
            .I(N__5475));
    InMux I__836 (
            .O(N__5487),
            .I(N__5472));
    LocalMux I__835 (
            .O(N__5484),
            .I(N__5469));
    InMux I__834 (
            .O(N__5483),
            .I(N__5466));
    Odrv4 I__833 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.N_352 ));
    Odrv4 I__832 (
            .O(N__5475),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__831 (
            .O(N__5472),
            .I(\U712_CHIP_RAM.N_352 ));
    Odrv4 I__830 (
            .O(N__5469),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__829 (
            .O(N__5466),
            .I(\U712_CHIP_RAM.N_352 ));
    InMux I__828 (
            .O(N__5455),
            .I(N__5449));
    InMux I__827 (
            .O(N__5454),
            .I(N__5446));
    InMux I__826 (
            .O(N__5453),
            .I(N__5435));
    InMux I__825 (
            .O(N__5452),
            .I(N__5435));
    LocalMux I__824 (
            .O(N__5449),
            .I(N__5430));
    LocalMux I__823 (
            .O(N__5446),
            .I(N__5430));
    InMux I__822 (
            .O(N__5445),
            .I(N__5423));
    InMux I__821 (
            .O(N__5444),
            .I(N__5423));
    InMux I__820 (
            .O(N__5443),
            .I(N__5423));
    InMux I__819 (
            .O(N__5442),
            .I(N__5418));
    InMux I__818 (
            .O(N__5441),
            .I(N__5418));
    InMux I__817 (
            .O(N__5440),
            .I(N__5415));
    LocalMux I__816 (
            .O(N__5435),
            .I(N__5412));
    Odrv4 I__815 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__814 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__813 (
            .O(N__5418),
            .I(\U712_CHIP_RAM.N_343 ));
    LocalMux I__812 (
            .O(N__5415),
            .I(\U712_CHIP_RAM.N_343 ));
    Odrv4 I__811 (
            .O(N__5412),
            .I(\U712_CHIP_RAM.N_343 ));
    CascadeMux I__810 (
            .O(N__5401),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_ ));
    InMux I__809 (
            .O(N__5398),
            .I(N__5386));
    InMux I__808 (
            .O(N__5397),
            .I(N__5386));
    InMux I__807 (
            .O(N__5396),
            .I(N__5378));
    InMux I__806 (
            .O(N__5395),
            .I(N__5371));
    InMux I__805 (
            .O(N__5394),
            .I(N__5371));
    InMux I__804 (
            .O(N__5393),
            .I(N__5371));
    InMux I__803 (
            .O(N__5392),
            .I(N__5368));
    InMux I__802 (
            .O(N__5391),
            .I(N__5365));
    LocalMux I__801 (
            .O(N__5386),
            .I(N__5362));
    InMux I__800 (
            .O(N__5385),
            .I(N__5355));
    InMux I__799 (
            .O(N__5384),
            .I(N__5355));
    InMux I__798 (
            .O(N__5383),
            .I(N__5355));
    InMux I__797 (
            .O(N__5382),
            .I(N__5350));
    InMux I__796 (
            .O(N__5381),
            .I(N__5350));
    LocalMux I__795 (
            .O(N__5378),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__794 (
            .O(N__5371),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__793 (
            .O(N__5368),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__792 (
            .O(N__5365),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__791 (
            .O(N__5362),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__790 (
            .O(N__5355),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__789 (
            .O(N__5350),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__788 (
            .O(N__5335),
            .I(N__5332));
    LocalMux I__787 (
            .O(N__5332),
            .I(N__5329));
    Span4Mux_v I__786 (
            .O(N__5329),
            .I(N__5325));
    InMux I__785 (
            .O(N__5328),
            .I(N__5322));
    Sp12to4 I__784 (
            .O(N__5325),
            .I(N__5317));
    LocalMux I__783 (
            .O(N__5322),
            .I(N__5317));
    Span12Mux_h I__782 (
            .O(N__5317),
            .I(N__5314));
    Span12Mux_v I__781 (
            .O(N__5314),
            .I(N__5311));
    Odrv12 I__780 (
            .O(N__5311),
            .I(AWEn_c));
    IoInMux I__779 (
            .O(N__5308),
            .I(N__5305));
    LocalMux I__778 (
            .O(N__5305),
            .I(N__5302));
    Span4Mux_s2_v I__777 (
            .O(N__5302),
            .I(N__5299));
    Span4Mux_v I__776 (
            .O(N__5299),
            .I(N__5296));
    Span4Mux_v I__775 (
            .O(N__5296),
            .I(N__5293));
    Span4Mux_v I__774 (
            .O(N__5293),
            .I(N__5289));
    InMux I__773 (
            .O(N__5292),
            .I(N__5286));
    Odrv4 I__772 (
            .O(N__5289),
            .I(DBDIR_c));
    LocalMux I__771 (
            .O(N__5286),
            .I(DBDIR_c));
    InMux I__770 (
            .O(N__5281),
            .I(N__5278));
    LocalMux I__769 (
            .O(N__5278),
            .I(\U712_CHIP_RAM.N_304 ));
    InMux I__768 (
            .O(N__5275),
            .I(N__5269));
    InMux I__767 (
            .O(N__5274),
            .I(N__5269));
    LocalMux I__766 (
            .O(N__5269),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0 ));
    InMux I__765 (
            .O(N__5266),
            .I(N__5263));
    LocalMux I__764 (
            .O(N__5263),
            .I(N__5260));
    Span4Mux_h I__763 (
            .O(N__5260),
            .I(N__5257));
    Odrv4 I__762 (
            .O(N__5257),
            .I(\U712_CHIP_RAM.N_399 ));
    CascadeMux I__761 (
            .O(N__5254),
            .I(\U712_CHIP_RAM.N_399_cascade_ ));
    InMux I__760 (
            .O(N__5251),
            .I(N__5248));
    LocalMux I__759 (
            .O(N__5248),
            .I(N__5245));
    Span4Mux_v I__758 (
            .O(N__5245),
            .I(N__5242));
    Odrv4 I__757 (
            .O(N__5242),
            .I(\U712_CHIP_RAM.N_277 ));
    CascadeMux I__756 (
            .O(N__5239),
            .I(\U712_CHIP_RAM.N_277_cascade_ ));
    CascadeMux I__755 (
            .O(N__5236),
            .I(\U712_CHIP_RAM.N_347_cascade_ ));
    InMux I__754 (
            .O(N__5233),
            .I(N__5229));
    CascadeMux I__753 (
            .O(N__5232),
            .I(N__5226));
    LocalMux I__752 (
            .O(N__5229),
            .I(N__5221));
    InMux I__751 (
            .O(N__5226),
            .I(N__5218));
    InMux I__750 (
            .O(N__5225),
            .I(N__5215));
    InMux I__749 (
            .O(N__5224),
            .I(N__5212));
    Span4Mux_h I__748 (
            .O(N__5221),
            .I(N__5209));
    LocalMux I__747 (
            .O(N__5218),
            .I(\U712_CHIP_RAM.N_353 ));
    LocalMux I__746 (
            .O(N__5215),
            .I(\U712_CHIP_RAM.N_353 ));
    LocalMux I__745 (
            .O(N__5212),
            .I(\U712_CHIP_RAM.N_353 ));
    Odrv4 I__744 (
            .O(N__5209),
            .I(\U712_CHIP_RAM.N_353 ));
    InMux I__743 (
            .O(N__5200),
            .I(N__5197));
    LocalMux I__742 (
            .O(N__5197),
            .I(N__5192));
    InMux I__741 (
            .O(N__5196),
            .I(N__5188));
    InMux I__740 (
            .O(N__5195),
            .I(N__5185));
    Span4Mux_h I__739 (
            .O(N__5192),
            .I(N__5182));
    InMux I__738 (
            .O(N__5191),
            .I(N__5179));
    LocalMux I__737 (
            .O(N__5188),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__736 (
            .O(N__5185),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv4 I__735 (
            .O(N__5182),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__734 (
            .O(N__5179),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__733 (
            .O(N__5170),
            .I(N__5164));
    InMux I__732 (
            .O(N__5169),
            .I(N__5161));
    InMux I__731 (
            .O(N__5168),
            .I(N__5158));
    InMux I__730 (
            .O(N__5167),
            .I(N__5155));
    InMux I__729 (
            .O(N__5164),
            .I(N__5152));
    LocalMux I__728 (
            .O(N__5161),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__727 (
            .O(N__5158),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__726 (
            .O(N__5155),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__725 (
            .O(N__5152),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__724 (
            .O(N__5143),
            .I(N__5138));
    InMux I__723 (
            .O(N__5142),
            .I(N__5134));
    InMux I__722 (
            .O(N__5141),
            .I(N__5131));
    InMux I__721 (
            .O(N__5138),
            .I(N__5128));
    InMux I__720 (
            .O(N__5137),
            .I(N__5125));
    LocalMux I__719 (
            .O(N__5134),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__718 (
            .O(N__5131),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__717 (
            .O(N__5128),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__716 (
            .O(N__5125),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__715 (
            .O(N__5116),
            .I(N__5110));
    InMux I__714 (
            .O(N__5115),
            .I(N__5110));
    LocalMux I__713 (
            .O(N__5110),
            .I(N__5106));
    InMux I__712 (
            .O(N__5109),
            .I(N__5103));
    Odrv4 I__711 (
            .O(N__5106),
            .I(\U712_CHIP_RAM.N_347 ));
    LocalMux I__710 (
            .O(N__5103),
            .I(\U712_CHIP_RAM.N_347 ));
    CascadeMux I__709 (
            .O(N__5098),
            .I(\U712_CHIP_RAM.N_343_cascade_ ));
    InMux I__708 (
            .O(N__5095),
            .I(N__5083));
    InMux I__707 (
            .O(N__5094),
            .I(N__5083));
    InMux I__706 (
            .O(N__5093),
            .I(N__5083));
    CascadeMux I__705 (
            .O(N__5092),
            .I(N__5080));
    CascadeMux I__704 (
            .O(N__5091),
            .I(N__5077));
    InMux I__703 (
            .O(N__5090),
            .I(N__5071));
    LocalMux I__702 (
            .O(N__5083),
            .I(N__5068));
    InMux I__701 (
            .O(N__5080),
            .I(N__5065));
    InMux I__700 (
            .O(N__5077),
            .I(N__5062));
    InMux I__699 (
            .O(N__5076),
            .I(N__5059));
    InMux I__698 (
            .O(N__5075),
            .I(N__5054));
    InMux I__697 (
            .O(N__5074),
            .I(N__5054));
    LocalMux I__696 (
            .O(N__5071),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__695 (
            .O(N__5068),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__694 (
            .O(N__5065),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__693 (
            .O(N__5062),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__692 (
            .O(N__5059),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__691 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__690 (
            .O(N__5041),
            .I(N__5031));
    InMux I__689 (
            .O(N__5040),
            .I(N__5028));
    InMux I__688 (
            .O(N__5039),
            .I(N__5025));
    InMux I__687 (
            .O(N__5038),
            .I(N__5022));
    InMux I__686 (
            .O(N__5037),
            .I(N__5019));
    InMux I__685 (
            .O(N__5036),
            .I(N__5014));
    InMux I__684 (
            .O(N__5035),
            .I(N__5014));
    InMux I__683 (
            .O(N__5034),
            .I(N__5011));
    LocalMux I__682 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__681 (
            .O(N__5028),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__680 (
            .O(N__5025),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__679 (
            .O(N__5022),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__678 (
            .O(N__5019),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__677 (
            .O(N__5014),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__676 (
            .O(N__5011),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__675 (
            .O(N__4996),
            .I(N__4991));
    InMux I__674 (
            .O(N__4995),
            .I(N__4988));
    InMux I__673 (
            .O(N__4994),
            .I(N__4985));
    LocalMux I__672 (
            .O(N__4991),
            .I(N__4981));
    LocalMux I__671 (
            .O(N__4988),
            .I(N__4978));
    LocalMux I__670 (
            .O(N__4985),
            .I(N__4975));
    InMux I__669 (
            .O(N__4984),
            .I(N__4972));
    Span4Mux_h I__668 (
            .O(N__4981),
            .I(N__4969));
    Odrv12 I__667 (
            .O(N__4978),
            .I(\U712_CHIP_RAM.N_391 ));
    Odrv4 I__666 (
            .O(N__4975),
            .I(\U712_CHIP_RAM.N_391 ));
    LocalMux I__665 (
            .O(N__4972),
            .I(\U712_CHIP_RAM.N_391 ));
    Odrv4 I__664 (
            .O(N__4969),
            .I(\U712_CHIP_RAM.N_391 ));
    IoInMux I__663 (
            .O(N__4960),
            .I(N__4957));
    LocalMux I__662 (
            .O(N__4957),
            .I(N__4954));
    IoSpan4Mux I__661 (
            .O(N__4954),
            .I(N__4951));
    Span4Mux_s0_h I__660 (
            .O(N__4951),
            .I(N__4948));
    Span4Mux_h I__659 (
            .O(N__4948),
            .I(N__4945));
    Sp12to4 I__658 (
            .O(N__4945),
            .I(N__4942));
    Span12Mux_v I__657 (
            .O(N__4942),
            .I(N__4938));
    InMux I__656 (
            .O(N__4941),
            .I(N__4935));
    Span12Mux_h I__655 (
            .O(N__4938),
            .I(N__4932));
    LocalMux I__654 (
            .O(N__4935),
            .I(N__4929));
    Span12Mux_h I__653 (
            .O(N__4932),
            .I(N__4926));
    Span12Mux_h I__652 (
            .O(N__4929),
            .I(N__4923));
    Odrv12 I__651 (
            .O(N__4926),
            .I(C3_c));
    Odrv12 I__650 (
            .O(N__4923),
            .I(C3_c));
    InMux I__649 (
            .O(N__4918),
            .I(N__4915));
    LocalMux I__648 (
            .O(N__4915),
            .I(N__4912));
    Span4Mux_v I__647 (
            .O(N__4912),
            .I(N__4909));
    Sp12to4 I__646 (
            .O(N__4909),
            .I(N__4906));
    Odrv12 I__645 (
            .O(N__4906),
            .I(A_c_9));
    InMux I__644 (
            .O(N__4903),
            .I(N__4900));
    LocalMux I__643 (
            .O(N__4900),
            .I(N__4897));
    Span4Mux_v I__642 (
            .O(N__4897),
            .I(N__4894));
    Sp12to4 I__641 (
            .O(N__4894),
            .I(N__4891));
    Span12Mux_h I__640 (
            .O(N__4891),
            .I(N__4888));
    Span12Mux_v I__639 (
            .O(N__4888),
            .I(N__4885));
    Odrv12 I__638 (
            .O(N__4885),
            .I(A_c_2));
    InMux I__637 (
            .O(N__4882),
            .I(N__4879));
    LocalMux I__636 (
            .O(N__4879),
            .I(N__4876));
    Span4Mux_v I__635 (
            .O(N__4876),
            .I(N__4873));
    Sp12to4 I__634 (
            .O(N__4873),
            .I(N__4870));
    Span12Mux_h I__633 (
            .O(N__4870),
            .I(N__4867));
    Odrv12 I__632 (
            .O(N__4867),
            .I(A_c_12));
    InMux I__631 (
            .O(N__4864),
            .I(N__4861));
    LocalMux I__630 (
            .O(N__4861),
            .I(N__4858));
    Span4Mux_v I__629 (
            .O(N__4858),
            .I(N__4855));
    Span4Mux_v I__628 (
            .O(N__4855),
            .I(N__4852));
    Sp12to4 I__627 (
            .O(N__4852),
            .I(N__4849));
    Odrv12 I__626 (
            .O(N__4849),
            .I(A_c_5));
    CascadeMux I__625 (
            .O(N__4846),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__624 (
            .O(N__4843),
            .I(N__4840));
    LocalMux I__623 (
            .O(N__4840),
            .I(N__4837));
    Span12Mux_h I__622 (
            .O(N__4837),
            .I(N__4834));
    Span12Mux_v I__621 (
            .O(N__4834),
            .I(N__4831));
    Odrv12 I__620 (
            .O(N__4831),
            .I(A_c_3));
    InMux I__619 (
            .O(N__4828),
            .I(N__4825));
    LocalMux I__618 (
            .O(N__4825),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ));
    InMux I__617 (
            .O(N__4822),
            .I(N__4819));
    LocalMux I__616 (
            .O(N__4819),
            .I(N__4816));
    Span4Mux_h I__615 (
            .O(N__4816),
            .I(N__4813));
    Span4Mux_v I__614 (
            .O(N__4813),
            .I(N__4810));
    Span4Mux_v I__613 (
            .O(N__4810),
            .I(N__4807));
    Span4Mux_v I__612 (
            .O(N__4807),
            .I(N__4804));
    Odrv4 I__611 (
            .O(N__4804),
            .I(RAMSPACEn_c));
    IoInMux I__610 (
            .O(N__4801),
            .I(N__4797));
    IoInMux I__609 (
            .O(N__4800),
            .I(N__4794));
    LocalMux I__608 (
            .O(N__4797),
            .I(N__4791));
    LocalMux I__607 (
            .O(N__4794),
            .I(N__4788));
    Span12Mux_s3_h I__606 (
            .O(N__4791),
            .I(N__4785));
    Span4Mux_s3_v I__605 (
            .O(N__4788),
            .I(N__4782));
    Span12Mux_v I__604 (
            .O(N__4785),
            .I(N__4779));
    Span4Mux_h I__603 (
            .O(N__4782),
            .I(N__4776));
    Span12Mux_h I__602 (
            .O(N__4779),
            .I(N__4773));
    Sp12to4 I__601 (
            .O(N__4776),
            .I(N__4770));
    Odrv12 I__600 (
            .O(N__4773),
            .I(N_246));
    Odrv12 I__599 (
            .O(N__4770),
            .I(N_246));
    IoInMux I__598 (
            .O(N__4765),
            .I(N__4762));
    LocalMux I__597 (
            .O(N__4762),
            .I(N__4759));
    IoSpan4Mux I__596 (
            .O(N__4759),
            .I(N__4756));
    Sp12to4 I__595 (
            .O(N__4756),
            .I(N__4753));
    Span12Mux_v I__594 (
            .O(N__4753),
            .I(N__4749));
    InMux I__593 (
            .O(N__4752),
            .I(N__4746));
    Odrv12 I__592 (
            .O(N__4749),
            .I(REGENn_c));
    LocalMux I__591 (
            .O(N__4746),
            .I(REGENn_c));
    InMux I__590 (
            .O(N__4741),
            .I(N__4737));
    InMux I__589 (
            .O(N__4740),
            .I(N__4734));
    LocalMux I__588 (
            .O(N__4737),
            .I(LATCH_REG));
    LocalMux I__587 (
            .O(N__4734),
            .I(LATCH_REG));
    InMux I__586 (
            .O(N__4729),
            .I(N__4726));
    LocalMux I__585 (
            .O(N__4726),
            .I(N__4723));
    Span12Mux_v I__584 (
            .O(N__4723),
            .I(N__4719));
    InMux I__583 (
            .O(N__4722),
            .I(N__4716));
    Odrv12 I__582 (
            .O(N__4719),
            .I(REG_CPU_CYCLE));
    LocalMux I__581 (
            .O(N__4716),
            .I(REG_CPU_CYCLE));
    IoInMux I__580 (
            .O(N__4711),
            .I(N__4708));
    LocalMux I__579 (
            .O(N__4708),
            .I(N__4705));
    Span4Mux_s3_v I__578 (
            .O(N__4705),
            .I(N__4702));
    Span4Mux_h I__577 (
            .O(N__4702),
            .I(N__4699));
    Sp12to4 I__576 (
            .O(N__4699),
            .I(N__4696));
    Span12Mux_h I__575 (
            .O(N__4696),
            .I(N__4692));
    InMux I__574 (
            .O(N__4695),
            .I(N__4689));
    Odrv12 I__573 (
            .O(N__4692),
            .I(ASn_c));
    LocalMux I__572 (
            .O(N__4689),
            .I(ASn_c));
    CascadeMux I__571 (
            .O(N__4684),
            .I(\U712_CHIP_RAM.N_400_cascade_ ));
    CascadeMux I__570 (
            .O(N__4681),
            .I(N__4678));
    InMux I__569 (
            .O(N__4678),
            .I(N__4674));
    InMux I__568 (
            .O(N__4677),
            .I(N__4671));
    LocalMux I__567 (
            .O(N__4674),
            .I(N__4666));
    LocalMux I__566 (
            .O(N__4671),
            .I(N__4666));
    Span4Mux_v I__565 (
            .O(N__4666),
            .I(N__4663));
    Odrv4 I__564 (
            .O(N__4663),
            .I(\U712_CHIP_RAM.N_266 ));
    CascadeMux I__563 (
            .O(N__4660),
            .I(\U712_CHIP_RAM.N_304_cascade_ ));
    InMux I__562 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__561 (
            .O(N__4654),
            .I(\U712_CHIP_RAM.N_249 ));
    InMux I__560 (
            .O(N__4651),
            .I(N__4646));
    InMux I__559 (
            .O(N__4650),
            .I(N__4643));
    InMux I__558 (
            .O(N__4649),
            .I(N__4639));
    LocalMux I__557 (
            .O(N__4646),
            .I(N__4636));
    LocalMux I__556 (
            .O(N__4643),
            .I(N__4633));
    InMux I__555 (
            .O(N__4642),
            .I(N__4630));
    LocalMux I__554 (
            .O(N__4639),
            .I(\U712_CHIP_RAM.N_355 ));
    Odrv4 I__553 (
            .O(N__4636),
            .I(\U712_CHIP_RAM.N_355 ));
    Odrv4 I__552 (
            .O(N__4633),
            .I(\U712_CHIP_RAM.N_355 ));
    LocalMux I__551 (
            .O(N__4630),
            .I(\U712_CHIP_RAM.N_355 ));
    InMux I__550 (
            .O(N__4621),
            .I(N__4617));
    InMux I__549 (
            .O(N__4620),
            .I(N__4614));
    LocalMux I__548 (
            .O(N__4617),
            .I(N__4610));
    LocalMux I__547 (
            .O(N__4614),
            .I(N__4607));
    InMux I__546 (
            .O(N__4613),
            .I(N__4604));
    Odrv4 I__545 (
            .O(N__4610),
            .I(\U712_CHIP_RAM.N_350_0 ));
    Odrv4 I__544 (
            .O(N__4607),
            .I(\U712_CHIP_RAM.N_350_0 ));
    LocalMux I__543 (
            .O(N__4604),
            .I(\U712_CHIP_RAM.N_350_0 ));
    CascadeMux I__542 (
            .O(N__4597),
            .I(\U712_CHIP_RAM.N_291_cascade_ ));
    InMux I__541 (
            .O(N__4594),
            .I(N__4591));
    LocalMux I__540 (
            .O(N__4591),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0 ));
    InMux I__539 (
            .O(N__4588),
            .I(N__4585));
    LocalMux I__538 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ));
    InMux I__537 (
            .O(N__4582),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__536 (
            .O(N__4579),
            .I(N__4576));
    LocalMux I__535 (
            .O(N__4576),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__534 (
            .O(N__4573),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__533 (
            .O(N__4570),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__532 (
            .O(N__4567),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__531 (
            .O(N__4564),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__530 (
            .O(N__4561),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__529 (
            .O(N__4558),
            .I(N__4551));
    InMux I__528 (
            .O(N__4557),
            .I(N__4551));
    CascadeMux I__527 (
            .O(N__4556),
            .I(N__4543));
    LocalMux I__526 (
            .O(N__4551),
            .I(N__4540));
    InMux I__525 (
            .O(N__4550),
            .I(N__4533));
    InMux I__524 (
            .O(N__4549),
            .I(N__4533));
    InMux I__523 (
            .O(N__4548),
            .I(N__4533));
    InMux I__522 (
            .O(N__4547),
            .I(N__4526));
    InMux I__521 (
            .O(N__4546),
            .I(N__4526));
    InMux I__520 (
            .O(N__4543),
            .I(N__4526));
    Odrv4 I__519 (
            .O(N__4540),
            .I(\U712_CHIP_RAM.N_100 ));
    LocalMux I__518 (
            .O(N__4533),
            .I(\U712_CHIP_RAM.N_100 ));
    LocalMux I__517 (
            .O(N__4526),
            .I(\U712_CHIP_RAM.N_100 ));
    InMux I__516 (
            .O(N__4519),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__515 (
            .O(N__4516),
            .I(N__4512));
    CEMux I__514 (
            .O(N__4515),
            .I(N__4509));
    LocalMux I__513 (
            .O(N__4512),
            .I(N__4506));
    LocalMux I__512 (
            .O(N__4509),
            .I(N__4503));
    Span4Mux_v I__511 (
            .O(N__4506),
            .I(N__4500));
    Span4Mux_v I__510 (
            .O(N__4503),
            .I(N__4497));
    Span4Mux_h I__509 (
            .O(N__4500),
            .I(N__4494));
    Odrv4 I__508 (
            .O(N__4497),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__507 (
            .O(N__4494),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__506 (
            .O(N__4489),
            .I(N__4481));
    InMux I__505 (
            .O(N__4488),
            .I(N__4481));
    InMux I__504 (
            .O(N__4487),
            .I(N__4476));
    InMux I__503 (
            .O(N__4486),
            .I(N__4476));
    LocalMux I__502 (
            .O(N__4481),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ));
    LocalMux I__501 (
            .O(N__4476),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ));
    CascadeMux I__500 (
            .O(N__4471),
            .I(N__4467));
    InMux I__499 (
            .O(N__4470),
            .I(N__4460));
    InMux I__498 (
            .O(N__4467),
            .I(N__4460));
    InMux I__497 (
            .O(N__4466),
            .I(N__4455));
    InMux I__496 (
            .O(N__4465),
            .I(N__4455));
    LocalMux I__495 (
            .O(N__4460),
            .I(\U712_CHIP_RAM.N_280 ));
    LocalMux I__494 (
            .O(N__4455),
            .I(\U712_CHIP_RAM.N_280 ));
    CascadeMux I__493 (
            .O(N__4450),
            .I(\U712_CHIP_RAM.N_301_cascade_ ));
    InMux I__492 (
            .O(N__4447),
            .I(N__4443));
    InMux I__491 (
            .O(N__4446),
            .I(N__4440));
    LocalMux I__490 (
            .O(N__4443),
            .I(\U712_CHIP_RAM.N_280_2 ));
    LocalMux I__489 (
            .O(N__4440),
            .I(\U712_CHIP_RAM.N_280_2 ));
    CascadeMux I__488 (
            .O(N__4435),
            .I(N__4432));
    InMux I__487 (
            .O(N__4432),
            .I(N__4429));
    LocalMux I__486 (
            .O(N__4429),
            .I(\U712_CHIP_RAM.N_192 ));
    CascadeMux I__485 (
            .O(N__4426),
            .I(\U712_CHIP_RAM.N_192_cascade_ ));
    InMux I__484 (
            .O(N__4423),
            .I(N__4420));
    LocalMux I__483 (
            .O(N__4420),
            .I(\U712_CHIP_RAM.N_215 ));
    CascadeMux I__482 (
            .O(N__4417),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_ ));
    InMux I__481 (
            .O(N__4414),
            .I(N__4411));
    LocalMux I__480 (
            .O(N__4411),
            .I(\U712_CHIP_RAM.N_345 ));
    IoInMux I__479 (
            .O(N__4408),
            .I(N__4405));
    LocalMux I__478 (
            .O(N__4405),
            .I(N__4402));
    IoSpan4Mux I__477 (
            .O(N__4402),
            .I(N__4399));
    Span4Mux_s2_v I__476 (
            .O(N__4399),
            .I(N__4396));
    Sp12to4 I__475 (
            .O(N__4396),
            .I(N__4393));
    Odrv12 I__474 (
            .O(N__4393),
            .I(LATCH_CLK_0_i));
    IoInMux I__473 (
            .O(N__4390),
            .I(N__4386));
    IoInMux I__472 (
            .O(N__4389),
            .I(N__4383));
    LocalMux I__471 (
            .O(N__4386),
            .I(N__4377));
    LocalMux I__470 (
            .O(N__4383),
            .I(N__4377));
    IoInMux I__469 (
            .O(N__4382),
            .I(N__4374));
    IoSpan4Mux I__468 (
            .O(N__4377),
            .I(N__4371));
    LocalMux I__467 (
            .O(N__4374),
            .I(N__4368));
    Sp12to4 I__466 (
            .O(N__4371),
            .I(N__4365));
    Span4Mux_s3_h I__465 (
            .O(N__4368),
            .I(N__4362));
    Span12Mux_v I__464 (
            .O(N__4365),
            .I(N__4359));
    Span4Mux_v I__463 (
            .O(N__4362),
            .I(N__4356));
    Span12Mux_h I__462 (
            .O(N__4359),
            .I(N__4353));
    Span4Mux_h I__461 (
            .O(N__4356),
            .I(N__4350));
    Odrv12 I__460 (
            .O(N__4353),
            .I(CLK40_PLL_iso_i));
    Odrv4 I__459 (
            .O(N__4350),
            .I(CLK40_PLL_iso_i));
    IoInMux I__458 (
            .O(N__4345),
            .I(N__4342));
    LocalMux I__457 (
            .O(N__4342),
            .I(N__4339));
    Span12Mux_s5_v I__456 (
            .O(N__4339),
            .I(N__4336));
    Odrv12 I__455 (
            .O(N__4336),
            .I(VBENn_c));
    InMux I__454 (
            .O(N__4333),
            .I(N__4330));
    LocalMux I__453 (
            .O(N__4330),
            .I(N__4327));
    Span12Mux_h I__452 (
            .O(N__4327),
            .I(N__4324));
    Odrv12 I__451 (
            .O(N__4324),
            .I(A_c_11));
    InMux I__450 (
            .O(N__4321),
            .I(N__4318));
    LocalMux I__449 (
            .O(N__4318),
            .I(N__4315));
    Span4Mux_h I__448 (
            .O(N__4315),
            .I(N__4312));
    Sp12to4 I__447 (
            .O(N__4312),
            .I(N__4309));
    Span12Mux_v I__446 (
            .O(N__4309),
            .I(N__4306));
    Odrv12 I__445 (
            .O(N__4306),
            .I(A_c_4));
    CascadeMux I__444 (
            .O(N__4303),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ));
    InMux I__443 (
            .O(N__4300),
            .I(N__4297));
    LocalMux I__442 (
            .O(N__4297),
            .I(\U712_CHIP_RAM.N_350 ));
    InMux I__441 (
            .O(N__4294),
            .I(N__4291));
    LocalMux I__440 (
            .O(N__4291),
            .I(\U712_CHIP_RAM.N_283 ));
    InMux I__439 (
            .O(N__4288),
            .I(N__4284));
    InMux I__438 (
            .O(N__4287),
            .I(N__4281));
    LocalMux I__437 (
            .O(N__4284),
            .I(N__4276));
    LocalMux I__436 (
            .O(N__4281),
            .I(N__4276));
    Odrv4 I__435 (
            .O(N__4276),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0 ));
    InMux I__434 (
            .O(N__4273),
            .I(N__4268));
    InMux I__433 (
            .O(N__4272),
            .I(N__4263));
    InMux I__432 (
            .O(N__4271),
            .I(N__4263));
    LocalMux I__431 (
            .O(N__4268),
            .I(\U712_CHIP_RAM.N_403 ));
    LocalMux I__430 (
            .O(N__4263),
            .I(\U712_CHIP_RAM.N_403 ));
    CascadeMux I__429 (
            .O(N__4258),
            .I(\U712_CHIP_RAM.N_389_cascade_ ));
    InMux I__428 (
            .O(N__4255),
            .I(N__4252));
    LocalMux I__427 (
            .O(N__4252),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ));
    CascadeMux I__426 (
            .O(N__4249),
            .I(\U712_CHIP_RAM.N_348_cascade_ ));
    InMux I__425 (
            .O(N__4246),
            .I(N__4243));
    LocalMux I__424 (
            .O(N__4243),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0 ));
    IoInMux I__423 (
            .O(N__4240),
            .I(N__4237));
    LocalMux I__422 (
            .O(N__4237),
            .I(N__4234));
    IoSpan4Mux I__421 (
            .O(N__4234),
            .I(N__4231));
    Sp12to4 I__420 (
            .O(N__4231),
            .I(N__4228));
    Span12Mux_s9_h I__419 (
            .O(N__4228),
            .I(N__4225));
    Span12Mux_h I__418 (
            .O(N__4225),
            .I(N__4221));
    InMux I__417 (
            .O(N__4224),
            .I(N__4218));
    Odrv12 I__416 (
            .O(N__4221),
            .I(CLK_EN_c));
    LocalMux I__415 (
            .O(N__4218),
            .I(CLK_EN_c));
    CascadeMux I__414 (
            .O(N__4213),
            .I(DBRn_c_i_cascade_));
    IoInMux I__413 (
            .O(N__4210),
            .I(N__4207));
    LocalMux I__412 (
            .O(N__4207),
            .I(N__4204));
    Span12Mux_s5_h I__411 (
            .O(N__4204),
            .I(N__4201));
    Odrv12 I__410 (
            .O(N__4201),
            .I(DBRn_c_i_0));
    CascadeMux I__409 (
            .O(N__4198),
            .I(\U712_CHIP_RAM.N_288_cascade_ ));
    CascadeMux I__408 (
            .O(N__4195),
            .I(\U712_CHIP_RAM.N_325_cascade_ ));
    CascadeMux I__407 (
            .O(N__4192),
            .I(\U712_CHIP_RAM.N_308_cascade_ ));
    CascadeMux I__406 (
            .O(N__4189),
            .I(\U712_CHIP_RAM.N_350_0_cascade_ ));
    CascadeMux I__405 (
            .O(N__4186),
            .I(\U712_CHIP_RAM.N_355_cascade_ ));
    IoInMux I__404 (
            .O(N__4183),
            .I(N__4180));
    LocalMux I__403 (
            .O(N__4180),
            .I(N__4177));
    Span4Mux_s2_v I__402 (
            .O(N__4177),
            .I(N__4174));
    Span4Mux_v I__401 (
            .O(N__4174),
            .I(N__4171));
    Span4Mux_h I__400 (
            .O(N__4171),
            .I(N__4168));
    Odrv4 I__399 (
            .O(N__4168),
            .I(CLK80_PLL_i_i));
    InMux I__398 (
            .O(N__4165),
            .I(N__4162));
    LocalMux I__397 (
            .O(N__4162),
            .I(N__4159));
    Span4Mux_v I__396 (
            .O(N__4159),
            .I(N__4156));
    Span4Mux_v I__395 (
            .O(N__4156),
            .I(N__4153));
    Sp12to4 I__394 (
            .O(N__4153),
            .I(N__4150));
    Odrv12 I__393 (
            .O(N__4150),
            .I(A_c_14));
    InMux I__392 (
            .O(N__4147),
            .I(N__4144));
    LocalMux I__391 (
            .O(N__4144),
            .I(N__4141));
    Span4Mux_v I__390 (
            .O(N__4141),
            .I(N__4138));
    Span4Mux_v I__389 (
            .O(N__4138),
            .I(N__4135));
    Sp12to4 I__388 (
            .O(N__4135),
            .I(N__4132));
    Odrv12 I__387 (
            .O(N__4132),
            .I(A_c_7));
    InMux I__386 (
            .O(N__4129),
            .I(N__4126));
    LocalMux I__385 (
            .O(N__4126),
            .I(N__4123));
    Span4Mux_v I__384 (
            .O(N__4123),
            .I(N__4120));
    Span4Mux_v I__383 (
            .O(N__4120),
            .I(N__4117));
    Sp12to4 I__382 (
            .O(N__4117),
            .I(N__4114));
    Odrv12 I__381 (
            .O(N__4114),
            .I(A_c_16));
    InMux I__380 (
            .O(N__4111),
            .I(N__4108));
    LocalMux I__379 (
            .O(N__4108),
            .I(N__4105));
    Span4Mux_v I__378 (
            .O(N__4105),
            .I(N__4102));
    Span4Mux_v I__377 (
            .O(N__4102),
            .I(N__4099));
    Sp12to4 I__376 (
            .O(N__4099),
            .I(N__4096));
    Odrv12 I__375 (
            .O(N__4096),
            .I(A_c_18));
    InMux I__374 (
            .O(N__4093),
            .I(N__4090));
    LocalMux I__373 (
            .O(N__4090),
            .I(N__4087));
    Sp12to4 I__372 (
            .O(N__4087),
            .I(N__4084));
    Span12Mux_v I__371 (
            .O(N__4084),
            .I(N__4081));
    Odrv12 I__370 (
            .O(N__4081),
            .I(A_c_15));
    InMux I__369 (
            .O(N__4078),
            .I(N__4075));
    LocalMux I__368 (
            .O(N__4075),
            .I(N__4072));
    Span4Mux_v I__367 (
            .O(N__4072),
            .I(N__4069));
    Span4Mux_v I__366 (
            .O(N__4069),
            .I(N__4066));
    Sp12to4 I__365 (
            .O(N__4066),
            .I(N__4063));
    Odrv12 I__364 (
            .O(N__4063),
            .I(A_c_8));
    CascadeMux I__363 (
            .O(N__4060),
            .I(\U712_CHIP_RAM.N_350_cascade_ ));
    CascadeMux I__362 (
            .O(N__4057),
            .I(\U712_CHIP_RAM.N_376_cascade_ ));
    CascadeMux I__361 (
            .O(N__4054),
            .I(\U712_CHIP_RAM.N_280_cascade_ ));
    IoInMux I__360 (
            .O(N__4051),
            .I(N__4048));
    LocalMux I__359 (
            .O(N__4048),
            .I(N__4045));
    Span4Mux_s0_v I__358 (
            .O(N__4045),
            .I(N__4042));
    Span4Mux_v I__357 (
            .O(N__4042),
            .I(N__4039));
    Sp12to4 I__356 (
            .O(N__4039),
            .I(N__4036));
    Span12Mux_h I__355 (
            .O(N__4036),
            .I(N__4033));
    Span12Mux_v I__354 (
            .O(N__4033),
            .I(N__4030));
    Odrv12 I__353 (
            .O(N__4030),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__6422));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__6423));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__6424));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__6426));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__6425));
    INV \INVU712_REG_SM.DBR_SYNC_0C  (
            .O(\INVU712_REG_SM.DBR_SYNC_0C_net ),
            .I(N__9081));
    INV \INVU712_REG_SM.REG_TACKC  (
            .O(\INVU712_REG_SM.REG_TACKC_net ),
            .I(N__9077));
    INV \INVU712_REG_SM.C1_SYNC_0C  (
            .O(\INVU712_REG_SM.C1_SYNC_0C_net ),
            .I(N__9086));
    INV \INVU712_REG_SM.C3_SYNC_1C  (
            .O(\INVU712_REG_SM.C3_SYNC_1C_net ),
            .I(N__9080));
    INV \INVU712_REG_SM.STATE_COUNTER_0C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_0C_net ),
            .I(N__9078));
    INV \INVU712_REG_SM.CYCLE_RUNC  (
            .O(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .I(N__9076));
    INV \INVU712_REG_SM.ASnC  (
            .O(\INVU712_REG_SM.ASnC_net ),
            .I(N__9085));
    INV \INVU712_REG_SM.REGENnC  (
            .O(\INVU712_REG_SM.REGENnC_net ),
            .I(N__9079));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    ICE_GB CLK40_PLL_derived_clock_RNIIOT (
            .USERSIGNALTOGLOBALBUFFER(N__8454),
            .GLOBALBUFFEROUTPUT(CLK40_PLL_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8770),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5952),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4210),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4960),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_6_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_6_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_6_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_6_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10393),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_6_1  (
            .in0(N__4165),
            .in1(N__4147),
            .in2(_gnd_net_),
            .in3(N__9237),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_2  (
            .in0(N__9238),
            .in1(N__4129),
            .in2(_gnd_net_),
            .in3(N__4111),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_6_4  (
            .in0(N__9239),
            .in1(N__4093),
            .in2(_gnd_net_),
            .in3(N__4078),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILSBFD_4_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILSBFD_4_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILSBFD_4_LC_7_7_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILSBFD_4_LC_7_7_0  (
            .in0(N__5094),
            .in1(N__5233),
            .in2(N__9003),
            .in3(N__4423),
            .lcout(\U712_CHIP_RAM.N_350 ),
            .ltout(\U712_CHIP_RAM.N_350_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_7_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4060),
            .in3(N__4271),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_7_2 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_7_2  (
            .in0(N__4465),
            .in1(N__4489),
            .in2(N__4057),
            .in3(N__8541),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10374),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_7_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_7_7_3 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_7_7_3  (
            .in0(N__6493),
            .in1(N__6613),
            .in2(N__6352),
            .in3(N__4446),
            .lcout(\U712_CHIP_RAM.N_280 ),
            .ltout(\U712_CHIP_RAM.N_280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1RLTB_4_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1RLTB_4_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1RLTB_4_LC_7_7_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1RLTB_4_LC_7_7_4  (
            .in0(N__5093),
            .in1(N__4677),
            .in2(N__4054),
            .in3(N__4287),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_5  (
            .in0(N__6215),
            .in1(N__8995),
            .in2(N__4435),
            .in3(N__5095),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_7_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_7_6  (
            .in0(N__4272),
            .in1(N__6614),
            .in2(N__4198),
            .in3(N__4447),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_7_7 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_7_7  (
            .in0(N__4488),
            .in1(N__4466),
            .in2(N__4195),
            .in3(N__9245),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10374),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISJJB2_7_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISJJB2_7_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISJJB2_7_LC_7_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISJJB2_7_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__5452),
            .in2(_gnd_net_),
            .in3(N__8992),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVENA4_1_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVENA4_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVENA4_1_LC_7_8_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVENA4_1_LC_7_8_1  (
            .in0(N__5453),
            .in1(N__5382),
            .in2(_gnd_net_),
            .in3(N__4246),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILAVHF_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILAVHF_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILAVHF_LC_7_8_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILAVHF_LC_7_8_2  (
            .in0(N__4255),
            .in1(N__8993),
            .in2(N__4192),
            .in3(N__6837),
            .lcout(\U712_CHIP_RAM.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7BNR1_7_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7BNR1_7_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7BNR1_7_LC_7_8_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7BNR1_7_LC_7_8_3  (
            .in0(N__5191),
            .in1(N__5137),
            .in2(N__5170),
            .in3(N__5381),
            .lcout(\U712_CHIP_RAM.N_350_0 ),
            .ltout(\U712_CHIP_RAM.N_350_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_7_8_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__5631),
            .in2(N__4189),
            .in3(N__6543),
            .lcout(\U712_CHIP_RAM.N_355 ),
            .ltout(\U712_CHIP_RAM.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_7_8_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_7_8_5  (
            .in0(N__8991),
            .in1(_gnd_net_),
            .in2(N__4186),
            .in3(N__6881),
            .lcout(\U712_CHIP_RAM.N_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_7_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_7_8_6  (
            .in0(N__4613),
            .in1(N__5483),
            .in2(_gnd_net_),
            .in3(N__6542),
            .lcout(\U712_CHIP_RAM.N_389 ),
            .ltout(\U712_CHIP_RAM.N_389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_7_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_7_8_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_7_8_7  (
            .in0(N__5707),
            .in1(N__4996),
            .in2(N__4258),
            .in3(N__4642),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_7_9_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_7_9_0  (
            .in0(N__6181),
            .in1(N__5074),
            .in2(_gnd_net_),
            .in3(N__5035),
            .lcout(\U712_CHIP_RAM.N_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_9_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_9_4  (
            .in0(N__6183),
            .in1(N__4995),
            .in2(_gnd_net_),
            .in3(N__4649),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10382),
            .ce(),
            .sr(N__10645));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_5  (
            .in0(N__5075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6182),
            .lcout(\U712_CHIP_RAM.N_348 ),
            .ltout(\U712_CHIP_RAM.N_348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRD202_3_LC_7_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRD202_3_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRD202_3_LC_7_9_6 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRD202_3_LC_7_9_6  (
            .in0(N__6988),
            .in1(N__5036),
            .in2(N__4249),
            .in3(N__5646),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_7_10_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_7_10_4 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_7_10_4  (
            .in0(N__7022),
            .in1(N__5517),
            .in2(N__6847),
            .in3(N__9628),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10386),
            .ce(),
            .sr(N__10640));
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_10_5 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_7_10_5  (
            .in0(N__5266),
            .in1(N__4224),
            .in2(N__5506),
            .in3(N__5251),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10386),
            .ce(),
            .sr(N__10640));
    defparam DBRn_ibuf_RNIBAB_LC_7_11_0.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_7_11_0 (
            .in0(N__8128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(DBRn_c_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4213),
            .in3(N__10663),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_14_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_14_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BUFFERS.LATCH_CLK_0_i_LC_7_14_2  (
            .in0(N__4741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6511),
            .lcout(LATCH_CLK_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_14_7.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_14_7.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_14_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_0_LC_7_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9094),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_8_5_7  (
            .in0(N__4729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9450),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_6_2  (
            .in0(N__4333),
            .in1(N__4321),
            .in2(_gnd_net_),
            .in3(N__9236),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_8_6_5 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_8_6_5  (
            .in0(N__4294),
            .in1(N__4621),
            .in2(N__9004),
            .in3(N__5505),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_0_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_0_LC_8_6_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_0_LC_8_6_6  (
            .in0(N__4994),
            .in1(N__8999),
            .in2(N__4303),
            .in3(N__4651),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_7_0 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_7_0  (
            .in0(N__4300),
            .in1(N__4487),
            .in2(N__4471),
            .in3(N__8606),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10372),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_1_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_1_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_1_LC_8_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_1_LC_8_7_1  (
            .in0(N__5393),
            .in1(N__4594),
            .in2(_gnd_net_),
            .in3(N__5443),
            .lcout(\U712_CHIP_RAM.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_7_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_7_2  (
            .in0(N__4288),
            .in1(N__4273),
            .in2(N__4681),
            .in3(N__5706),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_7_3 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_7_3  (
            .in0(N__4486),
            .in1(N__4470),
            .in2(N__4450),
            .in3(N__8497),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10372),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_8_7_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_8_7_4  (
            .in0(N__6286),
            .in1(N__8994),
            .in2(N__6224),
            .in3(N__6814),
            .lcout(\U712_CHIP_RAM.N_280_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_8_7_5 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_8_7_5  (
            .in0(N__5394),
            .in1(N__5444),
            .in2(N__5645),
            .in3(N__4414),
            .lcout(\U712_CHIP_RAM.N_192 ),
            .ltout(\U712_CHIP_RAM.N_192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_8_7_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_8_7_6  (
            .in0(N__5445),
            .in1(N__6214),
            .in2(N__4426),
            .in3(N__5395),
            .lcout(\U712_CHIP_RAM.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_0 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_0  (
            .in0(N__4546),
            .in1(N__8703),
            .in2(N__6552),
            .in3(N__4828),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10375),
            .ce(N__4516),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_8_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_8_1  (
            .in0(N__5038),
            .in1(N__5391),
            .in2(N__5644),
            .in3(N__6544),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_8_8_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_8_8_2  (
            .in0(N__5141),
            .in1(N__5195),
            .in2(N__4417),
            .in3(N__5168),
            .lcout(\U712_CHIP_RAM.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_3  (
            .in0(N__5724),
            .in1(N__4588),
            .in2(N__5232),
            .in3(N__4547),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10375),
            .ce(N__4516),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_8_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_8_4  (
            .in0(N__5225),
            .in1(N__4579),
            .in2(N__4556),
            .in3(N__5725),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10375),
            .ce(N__4516),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_4_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_4_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_4_LC_8_8_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_4_LC_8_8_5  (
            .in0(N__5629),
            .in1(N__8977),
            .in2(N__5092),
            .in3(N__6197),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_8_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__6548),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__5396),
            .in2(_gnd_net_),
            .in3(N__4582),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__5641),
            .in2(_gnd_net_),
            .in3(N__4573),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_9_3  (
            .in0(N__4548),
            .in1(N__5041),
            .in2(_gnd_net_),
            .in3(N__4570),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10379),
            .ce(N__4515),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_9_4  (
            .in0(N__4557),
            .in1(N__5090),
            .in2(_gnd_net_),
            .in3(N__4567),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10379),
            .ce(N__4515),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_9_5  (
            .in0(N__4549),
            .in1(N__5169),
            .in2(_gnd_net_),
            .in3(N__4564),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10379),
            .ce(N__4515),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_9_6  (
            .in0(N__4558),
            .in1(N__5196),
            .in2(_gnd_net_),
            .in3(N__4561),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10379),
            .ce(N__4515),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_9_7  (
            .in0(N__4550),
            .in1(N__5142),
            .in2(_gnd_net_),
            .in3(N__4519),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10379),
            .ce(N__4515),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPI372_4_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPI372_4_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPI372_4_LC_8_10_2 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPI372_4_LC_8_10_2  (
            .in0(N__6184),
            .in1(N__5115),
            .in2(N__5091),
            .in3(N__5397),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILMBG3_4_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILMBG3_4_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILMBG3_4_LC_8_10_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILMBG3_4_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4684),
            .in3(N__5487),
            .lcout(\U712_CHIP_RAM.N_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBO8O5_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBO8O5_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBO8O5_LC_8_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBO8O5_LC_8_10_4  (
            .in0(N__4657),
            .in1(N__5454),
            .in2(N__6210),
            .in3(N__5398),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(\U712_CHIP_RAM.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI34JU9_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI34JU9_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI34JU9_LC_8_10_5 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI34JU9_LC_8_10_5  (
            .in0(N__5687),
            .in1(N__6730),
            .in2(N__4660),
            .in3(N__5643),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC6723_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC6723_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC6723_LC_8_10_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIC6723_LC_8_10_6  (
            .in0(N__6274),
            .in1(N__5116),
            .in2(_gnd_net_),
            .in3(N__5524),
            .lcout(\U712_CHIP_RAM.N_249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_7  (
            .in0(N__6882),
            .in1(N__4650),
            .in2(_gnd_net_),
            .in3(N__5040),
            .lcout(\U712_CHIP_RAM.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_11_0 .LUT_INIT=16'b1110010011101100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_11_0  (
            .in0(N__8936),
            .in1(N__6285),
            .in2(N__6916),
            .in3(N__7002),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10387),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_1  (
            .in0(N__6765),
            .in1(N__4620),
            .in2(_gnd_net_),
            .in3(N__5500),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_2  (
            .in0(N__5501),
            .in1(N__5455),
            .in2(N__4597),
            .in3(N__5647),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMQBQ1_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMQBQ1_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMQBQ1_LC_8_11_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMQBQ1_LC_8_11_3  (
            .in0(N__6217),
            .in1(N__6861),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a3_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_11_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_11_6  (
            .in0(N__7567),
            .in1(N__5328),
            .in2(_gnd_net_),
            .in3(N__6284),
            .lcout(\U712_CHIP_RAM.N_234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_12_1 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_12_1  (
            .in0(N__4822),
            .in1(N__9411),
            .in2(N__5869),
            .in3(N__6337),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10389),
            .ce(),
            .sr(N__10618));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_8_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_x2_LC_8_13_2  (
            .in0(N__7831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7726),
            .lcout(\U712_BYTE_ENABLE.N_185_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_8_13_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_8_13_3  (
            .in0(N__7599),
            .in1(N__8052),
            .in2(_gnd_net_),
            .in3(N__5701),
            .lcout(N_246),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_LC_8_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_8_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_8_14_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.REGENn_LC_8_14_1  (
            .in0(N__4752),
            .in1(N__7339),
            .in2(_gnd_net_),
            .in3(N__5794),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REGENnC_net ),
            .ce(),
            .sr(N__10610));
    defparam \U712_REG_SM.LATCH_REG_LC_8_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LATCH_REG_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LATCH_REG_LC_8_14_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \U712_REG_SM.LATCH_REG_LC_8_14_3  (
            .in0(N__6900),
            .in1(N__5795),
            .in2(N__7600),
            .in3(N__4740),
            .lcout(LATCH_REG),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REGENnC_net ),
            .ce(),
            .sr(N__10610));
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_8_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_8_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_4_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6901),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REGENnC_net ),
            .ce(),
            .sr(N__10610));
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_14_5 .LUT_INIT=16'b0100111000000101;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_LC_8_14_5  (
            .in0(N__5772),
            .in1(N__4722),
            .in2(N__7477),
            .in3(N__5752),
            .lcout(REG_CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REGENnC_net ),
            .ce(),
            .sr(N__10610));
    defparam \U712_REG_SM.ASn_LC_8_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_8_15_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_8_15_0 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \U712_REG_SM.ASn_LC_8_15_0  (
            .in0(N__5797),
            .in1(N__5740),
            .in2(N__7297),
            .in3(N__4695),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.ASnC_net ),
            .ce(),
            .sr(N__10608));
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_15_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__4941),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.ASnC_net ),
            .ce(),
            .sr(N__10608));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_4 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_15_4  (
            .in0(N__5796),
            .in1(N__8045),
            .in2(_gnd_net_),
            .in3(N__7180),
            .lcout(REG_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.ASnC_net ),
            .ce(),
            .sr(N__10608));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_7_0  (
            .in0(N__4918),
            .in1(N__4903),
            .in2(_gnd_net_),
            .in3(N__9248),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_7_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__8600),
            .in2(_gnd_net_),
            .in3(N__8492),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_9_7_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_9_7_2  (
            .in0(N__8493),
            .in1(N__8611),
            .in2(_gnd_net_),
            .in3(N__9249),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_3  (
            .in0(N__9250),
            .in1(N__4882),
            .in2(_gnd_net_),
            .in3(N__4864),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_7_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_7_4  (
            .in0(N__9378),
            .in1(N__9251),
            .in2(N__4846),
            .in3(N__9658),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_7_5  (
            .in0(N__4843),
            .in1(N__9377),
            .in2(_gnd_net_),
            .in3(N__9682),
            .lcout(\U712_CHIP_RAM.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_8_0 .LUT_INIT=16'b0010101000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_8_0  (
            .in0(N__5224),
            .in1(N__6294),
            .in2(N__6229),
            .in3(N__6615),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_9_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__5442),
            .in2(_gnd_net_),
            .in3(N__5385),
            .lcout(\U712_CHIP_RAM.N_399 ),
            .ltout(\U712_CHIP_RAM.N_399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_9_8_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_9_8_2  (
            .in0(N__6773),
            .in1(N__9379),
            .in2(N__5254),
            .in3(N__4984),
            .lcout(\U712_CHIP_RAM.N_277 ),
            .ltout(\U712_CHIP_RAM.N_277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_8_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_8_3  (
            .in0(N__9380),
            .in1(N__5039),
            .in2(N__5239),
            .in3(N__5705),
            .lcout(\U712_CHIP_RAM.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__5034),
            .in2(_gnd_net_),
            .in3(N__5618),
            .lcout(\U712_CHIP_RAM.N_347 ),
            .ltout(\U712_CHIP_RAM.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_9_8_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_9_8_5  (
            .in0(N__8976),
            .in1(N__5441),
            .in2(N__5236),
            .in3(N__5384),
            .lcout(\U712_CHIP_RAM.N_353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ANR1_7_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ANR1_7_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ANR1_7_LC_9_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ANR1_7_LC_9_8_6  (
            .in0(N__5200),
            .in1(N__5167),
            .in2(N__5143),
            .in3(N__6541),
            .lcout(\U712_CHIP_RAM.N_343 ),
            .ltout(\U712_CHIP_RAM.N_343_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_1_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_1_LC_9_8_7 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_1_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__5109),
            .in2(N__5098),
            .in3(N__5383),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_9_9_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__5076),
            .in2(_gnd_net_),
            .in3(N__5037),
            .lcout(\U712_CHIP_RAM.N_391 ),
            .ltout(\U712_CHIP_RAM.N_391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNI0TLK1_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNI0TLK1_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNI0TLK1_LC_9_9_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNI0TLK1_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__6970),
            .in2(N__5527),
            .in3(N__5625),
            .lcout(\U712_CHIP_RAM.N_387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_9_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_9_9_4  (
            .in0(N__5274),
            .in1(N__6835),
            .in2(N__6987),
            .in3(N__5518),
            .lcout(DMA_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10376),
            .ce(),
            .sr(N__10632));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_9_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_9_9_5  (
            .in0(N__5630),
            .in1(N__5499),
            .in2(_gnd_net_),
            .in3(N__6971),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_9_9_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__5440),
            .in2(N__5401),
            .in3(N__5392),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_9_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_9_7 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_9_7  (
            .in0(N__5335),
            .in1(N__5292),
            .in2(N__6843),
            .in3(N__5275),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10376),
            .ce(),
            .sr(N__10632));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0  (
            .in0(N__6341),
            .in1(N__6492),
            .in2(N__6616),
            .in3(N__6842),
            .lcout(CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10380),
            .ce(N__6130),
            .sr(N__10625));
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_10_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_10_5  (
            .in0(N__6766),
            .in1(N__6736),
            .in2(_gnd_net_),
            .in3(N__5281),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_9_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_9_10_7  (
            .in0(N__6295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6228),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_11_0 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_11_0  (
            .in0(N__6270),
            .in1(N__6588),
            .in2(N__6487),
            .in3(N__6327),
            .lcout(\U712_CHIP_RAM.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_11_3  (
            .in0(N__5731),
            .in1(N__5718),
            .in2(N__5691),
            .in3(N__6841),
            .lcout(WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10383),
            .ce(),
            .sr(N__10619));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__5674),
            .in2(_gnd_net_),
            .in3(N__5642),
            .lcout(\U712_CHIP_RAM.N_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_9_11_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_9_11_7  (
            .in0(N__5566),
            .in1(N__8841),
            .in2(N__5560),
            .in3(N__5551),
            .lcout(CPU_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10383),
            .ce(),
            .sr(N__10619));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_9_12_1 .LUT_INIT=16'b0010101000001010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_9_12_1  (
            .in0(N__9412),
            .in1(N__7981),
            .in2(N__5542),
            .in3(N__7795),
            .lcout(\U712_BYTE_ENABLE.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_9_12_4 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_LC_9_12_4  (
            .in0(N__7845),
            .in1(N__7715),
            .in2(_gnd_net_),
            .in3(N__9413),
            .lcout(\U712_BYTE_ENABLE.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.CYCLE_RUN_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.CYCLE_RUN_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.CYCLE_RUN_LC_9_13_1 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \U712_REG_SM.CYCLE_RUN_LC_9_13_1  (
            .in0(N__7334),
            .in1(N__7401),
            .in2(N__7384),
            .in3(N__5883),
            .lcout(\U712_REG_SM.CYCLE_RUNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .ce(),
            .sr(N__10611));
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_5_LC_9_13_3  (
            .in0(N__5773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .ce(),
            .sr(N__10611));
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_6_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5533),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .ce(),
            .sr(N__10611));
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_13_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_3_LC_9_13_6  (
            .in0(N__8083),
            .in1(N__7428),
            .in2(_gnd_net_),
            .in3(N__7219),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .ce(),
            .sr(N__10611));
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_9_13_7 .LUT_INIT=16'b1100010111001100;
    LogicCell40 \U712_REG_SM.REG_WRITE_CYCLE_LC_9_13_7  (
            .in0(N__7555),
            .in1(N__7595),
            .in2(N__7405),
            .in3(N__7382),
            .lcout(REG_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.CYCLE_RUNC_net ),
            .ce(),
            .sr(N__10611));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_9_14_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_9_14_0  (
            .in0(N__5832),
            .in1(N__7292),
            .in2(_gnd_net_),
            .in3(N__7254),
            .lcout(\U712_REG_SM.N_229 ),
            .ltout(\U712_REG_SM.N_229_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_9_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_9_14_1 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_0_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__7376),
            .in2(N__5800),
            .in3(N__5793),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_0C_net ),
            .ce(),
            .sr(N__10609));
    defparam \U712_REG_SM.LDSn_RNO_1_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_9_14_2 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \U712_REG_SM.LDSn_RNO_1_LC_9_14_2  (
            .in0(N__7467),
            .in1(N__7885),
            .in2(N__7383),
            .in3(N__7562),
            .lcout(\U712_REG_SM.LDSn_7_iv_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5917),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_0C_net ),
            .ce(),
            .sr(N__10609));
    defparam \U712_REG_SM.C3_SYNC_RNIELLV_1_LC_9_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIELLV_1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIELLV_1_LC_9_14_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIELLV_1_LC_9_14_6  (
            .in0(N__7466),
            .in1(N__7291),
            .in2(_gnd_net_),
            .in3(N__7253),
            .lcout(\U712_REG_SM.LATCH_REG_0_sqmuxa ),
            .ltout(\U712_REG_SM.LATCH_REG_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_14_7 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_14_7  (
            .in0(N__7594),
            .in1(N__5771),
            .in2(N__5755),
            .in3(N__7175),
            .lcout(\U712_REG_SM.REG_CPU_CYCLE_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_15_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_15_0  (
            .in0(N__5746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_1C_net ),
            .ce(),
            .sr(N__10604));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_9_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_9_15_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_9_15_1  (
            .in0(N__7377),
            .in1(N__5828),
            .in2(N__7473),
            .in3(N__7252),
            .lcout(\U712_REG_SM.N_224 ),
            .ltout(\U712_REG_SM.N_224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNI5ITS1_2_LC_9_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNI5ITS1_2_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNI5ITS1_2_LC_9_15_2 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNI5ITS1_2_LC_9_15_2  (
            .in0(N__7290),
            .in1(_gnd_net_),
            .in2(N__5734),
            .in3(N__7216),
            .lcout(\U712_REG_SM.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_15_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__7289),
            .in2(_gnd_net_),
            .in3(N__7251),
            .lcout(\U712_REG_SM.N_209 ),
            .ltout(\U712_REG_SM.N_209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_9_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_9_15_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_9_15_4  (
            .in0(N__7884),
            .in1(N__6008),
            .in2(N__6034),
            .in3(N__7218),
            .lcout(),
            .ltout(\U712_REG_SM.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_LC_9_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_9_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_9_15_5 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \U712_REG_SM.LDSn_LC_9_15_5  (
            .in0(N__6009),
            .in1(N__6031),
            .in2(N__6022),
            .in3(N__5992),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_1C_net ),
            .ce(),
            .sr(N__10604));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_9_15_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_9_15_6  (
            .in0(N__5966),
            .in1(N__7217),
            .in2(N__7429),
            .in3(N__7960),
            .lcout(),
            .ltout(\U712_REG_SM.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_LC_9_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_9_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_9_15_7 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U712_REG_SM.UDSn_LC_9_15_7  (
            .in0(N__7513),
            .in1(N__5967),
            .in2(N__5995),
            .in3(N__5991),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_1C_net ),
            .ce(),
            .sr(N__10604));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_16_1  (
            .in0(N__5953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C1_SYNC_0C_net ),
            .ce(),
            .sr(N__10602));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_16_6 .LUT_INIT=16'b0011000001110101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_16_6  (
            .in0(N__5908),
            .in1(N__5887),
            .in2(N__5833),
            .in3(N__5862),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C1_SYNC_0C_net ),
            .ce(),
            .sr(N__10602));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_6_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_6_1  (
            .in0(N__9423),
            .in1(N__5809),
            .in2(N__9298),
            .in3(N__9616),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_7_0 .LUT_INIT=16'b0111001001110010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_7_0  (
            .in0(N__9808),
            .in1(N__9247),
            .in2(N__6115),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_7_3 .LUT_INIT=16'b1010110011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_7_3  (
            .in0(N__6106),
            .in1(N__9109),
            .in2(N__9453),
            .in3(N__8285),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_7_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_7_4  (
            .in0(N__6048),
            .in1(N__6078),
            .in2(N__6454),
            .in3(N__6063),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_7_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_7_5  (
            .in0(N__6105),
            .in1(N__9108),
            .in2(N__9454),
            .in3(N__8286),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_7_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_7_6  (
            .in0(N__8491),
            .in1(N__8607),
            .in2(N__8554),
            .in3(N__9246),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__6088),
            .in2(_gnd_net_),
            .in3(N__6082),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__6079),
            .in2(_gnd_net_),
            .in3(N__6067),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__6064),
            .in2(_gnd_net_),
            .in3(N__6052),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__6049),
            .in2(_gnd_net_),
            .in3(N__6037),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__6453),
            .in2(_gnd_net_),
            .in3(N__6439),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_8_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__6657),
            .in2(_gnd_net_),
            .in3(N__6436),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__6672),
            .in2(_gnd_net_),
            .in3(N__6433),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__6636),
            .in2(_gnd_net_),
            .in3(N__6430),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6427),
            .ce(),
            .sr(N__6403));
    defparam \U712_CHIP_RAM.BANK0_esr_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_10_9_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_LC_10_9_0  (
            .in0(N__6298),
            .in1(N__6358),
            .in2(N__6836),
            .in3(N__8139),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10373),
            .ce(N__6688),
            .sr(N__10626));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_10_9_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_10_9_1  (
            .in0(N__6373),
            .in1(N__6297),
            .in2(N__10993),
            .in3(N__6304),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_10_9_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_10_9_2  (
            .in0(N__6815),
            .in1(N__6594),
            .in2(N__6351),
            .in3(N__6491),
            .lcout(\U712_CHIP_RAM.N_405 ),
            .ltout(\U712_CHIP_RAM.N_405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_9_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__6296),
            .in2(N__6232),
            .in3(N__6216),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_9_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_9_4  (
            .in0(N__10662),
            .in1(N__6775),
            .in2(N__6133),
            .in3(N__6735),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_10_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_10_9_5  (
            .in0(N__6886),
            .in1(N__6862),
            .in2(_gnd_net_),
            .in3(N__6816),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_9_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_9_6  (
            .in0(N__6774),
            .in1(N__6734),
            .in2(N__6700),
            .in3(N__6697),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_9_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6691),
            .in3(N__10661),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_10_1  (
            .in0(N__6673),
            .in1(N__6658),
            .in2(N__6643),
            .in3(N__6625),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10377),
            .ce(),
            .sr(N__10620));
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_10_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_LC_10_10_6  (
            .in0(N__6981),
            .in1(N__6565),
            .in2(N__6559),
            .in3(N__6504),
            .lcout(LATCH_RAM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10377),
            .ce(),
            .sr(N__10620));
    defparam DBR_SYNC_1_LC_10_11_0.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_10_11_0.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_10_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_10_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6460),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10381),
            .ce(),
            .sr(N__10614));
    defparam DBR_SYNC_0_LC_10_11_6.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_10_11_6.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_10_11_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_10_11_6 (
            .in0(N__8127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10381),
            .ce(),
            .sr(N__10614));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_1_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_1_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_1_LC_10_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_1_LC_10_12_0  (
            .in0(N__10459),
            .in1(N__7006),
            .in2(_gnd_net_),
            .in3(N__7046),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_12_1 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \U712_BYTE_ENABLE.N_58_i_LC_10_12_1  (
            .in0(N__7793),
            .in1(N__7099),
            .in2(N__7159),
            .in3(N__7087),
            .lcout(N_58_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_10_12_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_10_12_2  (
            .in0(N__7722),
            .in1(N__9448),
            .in2(_gnd_net_),
            .in3(N__7982),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_56_i_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_10_12_3 .LUT_INIT=16'b0101010001010101;
    LogicCell40 \U712_BYTE_ENABLE.N_56_i_LC_10_12_3  (
            .in0(N__7129),
            .in1(N__10509),
            .in2(N__7050),
            .in3(N__7003),
            .lcout(N_56_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_10_12_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_10_12_4  (
            .in0(N__10458),
            .in1(N__7005),
            .in2(_gnd_net_),
            .in3(N__7045),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_54_i_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_54_i_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_54_i_LC_10_12_5 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_BYTE_ENABLE.N_54_i_LC_10_12_5  (
            .in0(N__7792),
            .in1(N__7098),
            .in2(N__7090),
            .in3(N__7086),
            .lcout(N_54_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_10_12_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_10_12_6  (
            .in0(N__9449),
            .in1(N__7794),
            .in2(_gnd_net_),
            .in3(N__7983),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_60_i_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_60_i_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_60_i_LC_10_12_7 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \U712_BYTE_ENABLE.N_60_i_LC_10_12_7  (
            .in0(N__7044),
            .in1(N__7004),
            .in2(N__6940),
            .in3(N__10510),
            .lcout(N_60_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__8353),
            .in2(_gnd_net_),
            .in3(N__10407),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_3  (
            .in0(N__7491),
            .in1(N__7462),
            .in2(_gnd_net_),
            .in3(N__6899),
            .lcout(\U712_REG_SM.un15_0_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_5  (
            .in0(N__7490),
            .in1(_gnd_net_),
            .in2(N__7224),
            .in3(N__7593),
            .lcout(\U712_REG_SM.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_1_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_10_13_6 .LUT_INIT=16'b1111110111110000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_1_LC_10_13_6  (
            .in0(N__7566),
            .in1(N__7987),
            .in2(N__7472),
            .in3(N__7372),
            .lcout(\U712_REG_SM.UDSn_7_iv_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_14_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_14_2  (
            .in0(N__7504),
            .in1(N__7176),
            .in2(N__8806),
            .in3(N__7498),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_TACKC_net ),
            .ce(),
            .sr(N__10605));
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_14_4 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_7_LC_10_14_4  (
            .in0(N__7471),
            .in1(N__7293),
            .in2(N__7258),
            .in3(N__7492),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_TACKC_net ),
            .ce(),
            .sr(N__10605));
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_6 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_2_LC_10_14_6  (
            .in0(N__8082),
            .in1(N__7427),
            .in2(N__7225),
            .in3(N__7335),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_TACKC_net ),
            .ce(),
            .sr(N__10605));
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_10_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_1_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__7400),
            .in2(_gnd_net_),
            .in3(N__7381),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_TACKC_net ),
            .ce(),
            .sr(N__10605));
    defparam TACKn_obuft_RNO_LC_10_15_2.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_10_15_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_10_15_2 (
            .in0(N__8338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_858_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_10_15_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_10_15_7  (
            .in0(N__7288),
            .in1(N__7250),
            .in2(N__8078),
            .in3(N__7223),
            .lcout(\U712_REG_SM.REG_TACK_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_0_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8120),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.DBR_SYNC_0C_net ),
            .ce(),
            .sr(N__10601));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8089),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.DBR_SYNC_0C_net ),
            .ce(),
            .sr(N__10601));
    defparam \U712_BYTE_ENABLE.LLBE_0_0_a2_LC_10_18_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_a2_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_a2_LC_10_18_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_0_a2_LC_10_18_0  (
            .in0(N__7857),
            .in1(N__7984),
            .in2(_gnd_net_),
            .in3(N__7711),
            .lcout(N_386),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_10_18_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_10_18_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_10_18_1  (
            .in0(N__10456),
            .in1(N__10502),
            .in2(_gnd_net_),
            .in3(N__8056),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_118_i_LC_10_19_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_118_i_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_118_i_LC_10_19_6 .LUT_INIT=16'b0100100001011010;
    LogicCell40 \U712_BYTE_ENABLE.N_118_i_LC_10_19_6  (
            .in0(N__7710),
            .in1(N__7985),
            .in2(N__7858),
            .in3(N__7750),
            .lcout(N_118_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_10_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_10_20_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_LC_10_20_4  (
            .in0(N__7986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7779),
            .lcout(U712_BYTE_ENABLE_UUBE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_10_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_0_LC_10_20_5 .LUT_INIT=16'b1010101110101110;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_0_LC_10_20_5  (
            .in0(N__7876),
            .in1(N__7846),
            .in2(N__7790),
            .in3(N__7708),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_0_0_LC_10_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_0_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_0_LC_10_20_7 .LUT_INIT=16'b1011101011101010;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_0_LC_10_20_7  (
            .in0(N__7877),
            .in1(N__7847),
            .in2(N__7791),
            .in3(N__7709),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_5_5 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_11_5_5  (
            .in0(N__7639),
            .in1(N__9456),
            .in2(N__8299),
            .in3(N__8161),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10363),
            .ce(N__9728),
            .sr(N__10646));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_11_5_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_11_5_7  (
            .in0(N__8298),
            .in1(N__8272),
            .in2(N__10063),
            .in3(N__9457),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10363),
            .ce(N__9728),
            .sr(N__10646));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_11_6_3  (
            .in0(N__8212),
            .in1(N__8206),
            .in2(_gnd_net_),
            .in3(N__8239),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10368),
            .ce(N__9735),
            .sr(N__10641));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_1 .LUT_INIT=16'b0000101001001010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_1  (
            .in0(N__9816),
            .in1(N__10302),
            .in2(N__9281),
            .in3(N__9437),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_4 .LUT_INIT=16'b0011001111111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_4  (
            .in0(N__10303),
            .in1(N__9262),
            .in2(N__9455),
            .in3(N__9817),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_7_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_11_7_7  (
            .in0(N__8200),
            .in1(_gnd_net_),
            .in2(N__8194),
            .in3(N__8185),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10370),
            .ce(N__9725),
            .sr(N__10633));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_11_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_11_8_0  (
            .in0(N__10137),
            .in1(N__10195),
            .in2(_gnd_net_),
            .in3(N__10992),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10717),
            .ce(N__10688),
            .sr(N__10627));
    defparam \U712_CHIP_RAM.DMA_A20_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_11_10_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_11_10_6  (
            .in0(N__8152),
            .in1(N__10988),
            .in2(N__10138),
            .in3(N__8140),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10615));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_11_1  (
            .in0(N__8453),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9045),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10378),
            .ce(),
            .sr(N__10612));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8386),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10378),
            .ce(),
            .sr(N__10612));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_11_7 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_11_11_7  (
            .in0(N__8397),
            .in1(N__8370),
            .in2(N__8455),
            .in3(N__9046),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10378),
            .ce(),
            .sr(N__10612));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_4  (
            .in0(N__8385),
            .in1(N__9037),
            .in2(N__8863),
            .in3(N__8369),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_13_1 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_11_13_1  (
            .in0(N__9039),
            .in1(N__8861),
            .in2(N__9013),
            .in3(N__8800),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10384),
            .ce(),
            .sr(N__10606));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8374),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10384),
            .ce(),
            .sr(N__10606));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10408),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10384),
            .ce(),
            .sr(N__10606));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_13_5 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_11_13_5  (
            .in0(N__9038),
            .in1(N__8875),
            .in2(N__8347),
            .in3(N__8799),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10384),
            .ce(),
            .sr(N__10606));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_14_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_14_6 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_14_6  (
            .in0(N__8975),
            .in1(N__8805),
            .in2(N__8862),
            .in3(N__8893),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10388),
            .ce(N__8752),
            .sr(N__10603));
    defparam \U712_CHIP_RAM.RASn_LC_12_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_12_4_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_12_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8619),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10361),
            .ce(),
            .sr(N__10644));
    defparam \U712_CHIP_RAM.WEn_LC_12_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8506),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10361),
            .ce(),
            .sr(N__10644));
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8565),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10361),
            .ce(),
            .sr(N__10644));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_5_1  (
            .in0(N__8620),
            .in1(N__9296),
            .in2(N__8566),
            .in3(N__8505),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10362),
            .ce(N__9727),
            .sr(N__10639));
    defparam CONSTANT_ONE_LUT4_LC_12_6_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_6_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_6_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_6_7  (
            .in0(N__9424),
            .in1(N__8680),
            .in2(N__9301),
            .in3(N__9118),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_7_0  (
            .in0(N__8671),
            .in1(N__9253),
            .in2(_gnd_net_),
            .in3(N__8650),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1  (
            .in0(N__9255),
            .in1(N__9442),
            .in2(N__8635),
            .in3(N__9637),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3  (
            .in0(N__9254),
            .in1(N__9441),
            .in2(N__8632),
            .in3(N__9124),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_7_4 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_7_4  (
            .in0(N__8618),
            .in1(N__9252),
            .in2(N__8564),
            .in3(N__8504),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_7_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_7_5  (
            .in0(N__10660),
            .in1(_gnd_net_),
            .in2(N__9127),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_8_3  (
            .in0(N__9901),
            .in1(N__10291),
            .in2(_gnd_net_),
            .in3(N__10980),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10691),
            .sr(N__10617));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_7  (
            .in0(N__10048),
            .in1(N__10002),
            .in2(_gnd_net_),
            .in3(N__10981),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10691),
            .sr(N__10617));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_9_3  (
            .in0(N__10983),
            .in1(N__9889),
            .in2(_gnd_net_),
            .in3(N__10290),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10715),
            .ce(N__10689),
            .sr(N__10613));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6  (
            .in0(N__9093),
            .in1(N__9036),
            .in2(_gnd_net_),
            .in3(N__8892),
            .lcout(\U712_CYCLE_TERM.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8949),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__8950),
            .in2(_gnd_net_),
            .in3(N__8891),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_227_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_6 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_6  (
            .in0(N__8874),
            .in1(N__8854),
            .in2(N__8809),
            .in3(N__8804),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_227_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_14_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_14_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8773),
            .in3(N__8763),
            .lcout(\U712_CYCLE_TERM.N_227_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_13_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_13_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9297),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10364),
            .ce(),
            .sr(N__10647));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_6_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_6_2  (
            .in0(N__9451),
            .in1(N__9300),
            .in2(N__9583),
            .in3(N__9646),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_13_6_3  (
            .in0(N__9839),
            .in1(N__9777),
            .in2(N__9568),
            .in3(N__10729),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10369),
            .ce(N__9736),
            .sr(N__10642));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_6_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_6_4  (
            .in0(N__9776),
            .in1(N__10201),
            .in2(N__9841),
            .in3(N__9544),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10369),
            .ce(N__9736),
            .sr(N__10642));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_5  (
            .in0(N__9299),
            .in1(N__9517),
            .in2(N__9670),
            .in3(N__9452),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_6_6  (
            .in0(N__9778),
            .in1(N__10147),
            .in2(N__9505),
            .in3(N__9840),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10369),
            .ce(N__9736),
            .sr(N__10642));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_7_4 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_13_7_4  (
            .in0(N__9774),
            .in1(N__9838),
            .in2(N__10246),
            .in3(N__9481),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10371),
            .ce(N__9726),
            .sr(N__10634));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__9430),
            .in2(_gnd_net_),
            .in3(N__9261),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6  (
            .in0(N__9847),
            .in1(N__9837),
            .in2(N__9157),
            .in3(N__9154),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10371),
            .ce(N__9726),
            .sr(N__10634));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_7_7 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_7_7  (
            .in0(N__9836),
            .in1(N__9787),
            .in2(N__9946),
            .in3(N__9775),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10371),
            .ce(N__9726),
            .sr(N__10634));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2  (
            .in0(N__10984),
            .in1(N__10289),
            .in2(_gnd_net_),
            .in3(N__10047),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10693),
            .sr(N__10628));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_4  (
            .in0(N__10987),
            .in1(N__10136),
            .in2(_gnd_net_),
            .in3(N__10194),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10693),
            .sr(N__10628));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5  (
            .in0(N__10237),
            .in1(N__10001),
            .in2(_gnd_net_),
            .in3(N__10985),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10693),
            .sr(N__10628));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7  (
            .in0(N__10193),
            .in1(N__10777),
            .in2(_gnd_net_),
            .in3(N__10986),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10693),
            .sr(N__10628));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_4  (
            .in0(N__10828),
            .in1(N__10233),
            .in2(_gnd_net_),
            .in3(N__10982),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10692),
            .sr(N__10621));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0  (
            .in0(N__9893),
            .in1(N__10954),
            .in2(_gnd_net_),
            .in3(N__9930),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10690),
            .sr(N__10616));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_10_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_10_4  (
            .in0(N__10970),
            .in1(N__10822),
            .in2(N__10765),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10690),
            .sr(N__10616));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_2  (
            .in0(N__10508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10457),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10385),
            .ce(),
            .sr(N__10607));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_0  (
            .in0(N__10827),
            .in1(N__10232),
            .in2(_gnd_net_),
            .in3(N__10926),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10716),
            .ce(N__10695),
            .sr(N__10643));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2  (
            .in0(N__10924),
            .in1(N__10034),
            .in2(_gnd_net_),
            .in3(N__10279),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10716),
            .ce(N__10695),
            .sr(N__10643));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_4  (
            .in0(N__10003),
            .in1(N__10231),
            .in2(_gnd_net_),
            .in3(N__10925),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10716),
            .ce(N__10695),
            .sr(N__10643));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_7  (
            .in0(N__10927),
            .in1(N__10776),
            .in2(_gnd_net_),
            .in3(N__10189),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10716),
            .ce(N__10695),
            .sr(N__10643));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_4  (
            .in0(N__10922),
            .in1(N__10120),
            .in2(_gnd_net_),
            .in3(N__10075),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10713),
            .ce(N__10694),
            .sr(N__10635));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_5  (
            .in0(N__10033),
            .in1(N__9997),
            .in2(_gnd_net_),
            .in3(N__10921),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10713),
            .ce(N__10694),
            .sr(N__10635));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_8_7  (
            .in0(N__9937),
            .in1(N__9900),
            .in2(_gnd_net_),
            .in3(N__10920),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10713),
            .ce(N__10694),
            .sr(N__10635));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_7_0  (
            .in0(N__10923),
            .in1(N__10826),
            .in2(_gnd_net_),
            .in3(N__10775),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10714),
            .ce(N__10696),
            .sr(N__10648));
endmodule // U712_TOP

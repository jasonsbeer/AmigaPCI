-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 12 2025 19:38:10

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TEAn : in std_logic;
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    TBIn : in std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__12664\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \N_267_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_266_i\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_0\ : std_logic;
signal \N_247_i\ : std_logic;
signal \N_249_i\ : std_logic;
signal \N_251_i\ : std_logic;
signal \N_253_i\ : std_logic;
signal \N_254_i\ : std_logic;
signal \N_252_i\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \N_264_i\ : std_logic;
signal \N_262_i\ : std_logic;
signal \N_258_i\ : std_logic;
signal \N_246_i\ : std_logic;
signal \N_248_i\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un2_D_LL_AMIGA_5\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un2_D_LM_AMIGA_6\ : std_logic;
signal \N_242_i\ : std_logic;
signal \N_260_i\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \N_239_i\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \N_263_i\ : std_logic;
signal \N_265_i\ : std_logic;
signal \N_257_i\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un2_D_LM_AMIGA_5\ : std_logic;
signal \N_250_i\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un2_D_LM_AMIGA_7\ : std_logic;
signal \N_238_i\ : std_logic;
signal \N_241_i\ : std_logic;
signal \N_261_i\ : std_logic;
signal \N_256_i\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un2_D_LM_AMIGA_2\ : std_logic;
signal \N_245_i\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un2_D_LM_AMIGA_4\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \N_259_i\ : std_logic;
signal \N_240_i\ : std_logic;
signal \N_243_i\ : std_logic;
signal \N_237_i\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un2_D_LL_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un2_D_LM_AMIGA_1\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un2_D_LM_AMIGA_3\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un2_D_LM_AMIGA_0\ : std_logic;
signal \N_268_i\ : std_logic;
signal \N_255_i\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \N_244_i\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un2_D_LL_AMIGA_3\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.N_67\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \BGn_c\ : std_logic;
signal \U111_CYCLE_SM.TS_DELAYZ0\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \LBENn_c_i_0\ : std_logic;
signal \U111_CYCLE_SM.N_33\ : std_logic;
signal \U111_CYCLE_SM.N_49\ : std_logic;
signal \U111_CYCLE_SM.N_75\ : std_logic;
signal \U111_CYCLE_SM.N_75_cascade_\ : std_logic;
signal \U111_CYCLE_SM.LATCH_EN_5\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \N_211_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \N_207_i\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un2_D_LL_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un2_D_LL_AMIGA_2\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \N_231_i\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un2_D_LL_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.N_60_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_46_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.N_39\ : std_logic;
signal \U111_CYCLE_SM.N_40\ : std_logic;
signal \U111_CYCLE_SM.N_40_cascade_\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.N_55_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_73\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \U111_CYCLE_SM.N_57_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.N_42\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \N_210_i\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \N_206_i\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \TAn_1_i\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un2_D_LL_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un2_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \U111_CYCLE_SM.N_40_i_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \N_224_i\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \N_216_i\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \N_219_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \N_220_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \N_234_i\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.N_44\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_g_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \N_232_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \N_223_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \N_205_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \N_212_i\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep31_i_ess\ : std_logic;
signal \N_236_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \N_227_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \N_218_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \N_209_i\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \N_233_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \N_235_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \N_222_i\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \N_230_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \N_215_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \N_226_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \N_229_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \N_214_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \N_217_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \N_213_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \N_228_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \N_225_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \N_208_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \N_221_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    A_AMIGA <= \A_AMIGA_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    \RnW_wire\ <= RnW;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__5291\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__12664\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__12664\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12648\,
            DIN => \N__12647\,
            DOUT => \N__12646\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12648\,
            PADOUT => \N__12647\,
            PADIN => \N__12646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12639\,
            DIN => \N__12638\,
            DOUT => \N__12637\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12639\,
            PADOUT => \N__12638\,
            PADIN => \N__12637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7982\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__7205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12630\,
            DIN => \N__12629\,
            DOUT => \N__12628\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12630\,
            PADOUT => \N__12629\,
            PADIN => \N__12628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4238\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__7613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12621\,
            DIN => \N__12620\,
            DOUT => \N__12619\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12621\,
            PADOUT => \N__12620\,
            PADIN => \N__12619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6392\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__8786\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12612\,
            DIN => \N__12611\,
            DOUT => \N__12610\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12612\,
            PADOUT => \N__12611\,
            PADIN => \N__12610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12603\,
            DIN => \N__12602\,
            DOUT => \N__12601\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12603\,
            PADOUT => \N__12602\,
            PADIN => \N__12601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4697\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__4463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12594\,
            DIN => \N__12593\,
            DOUT => \N__12592\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12594\,
            PADOUT => \N__12593\,
            PADIN => \N__12592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12585\,
            DIN => \N__12584\,
            DOUT => \N__12583\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12585\,
            PADOUT => \N__12584\,
            PADIN => \N__12583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4835\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__7967\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12576\,
            DIN => \N__12575\,
            DOUT => \N__12574\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12576\,
            PADOUT => \N__12575\,
            PADIN => \N__12574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11576\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__4763\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12567\,
            DIN => \N__12566\,
            DOUT => \N__12565\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12567\,
            PADOUT => \N__12566\,
            PADIN => \N__12565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6123\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12558\,
            DIN => \N__12557\,
            DOUT => \N__12556\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12558\,
            PADOUT => \N__12557\,
            PADIN => \N__12556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11678\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__8972\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12549\,
            DIN => \N__12548\,
            DOUT => \N__12547\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12549\,
            PADOUT => \N__12548\,
            PADIN => \N__12547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12540\,
            DIN => \N__12539\,
            DOUT => \N__12538\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12540\,
            PADOUT => \N__12539\,
            PADIN => \N__12538\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5675\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__8561\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12531\,
            DIN => \N__12530\,
            DOUT => \N__12529\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12531\,
            PADOUT => \N__12530\,
            PADIN => \N__12529\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10094\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12522\,
            DIN => \N__12521\,
            DOUT => \N__12520\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12522\,
            PADOUT => \N__12521\,
            PADIN => \N__12520\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12513\,
            DIN => \N__12512\,
            DOUT => \N__12511\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12513\,
            PADOUT => \N__12512\,
            PADIN => \N__12511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12504\,
            DIN => \N__12503\,
            DOUT => \N__12502\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12504\,
            PADOUT => \N__12503\,
            PADIN => \N__12502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10835\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__7877\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12495\,
            DIN => \N__12494\,
            DOUT => \N__12493\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12495\,
            PADOUT => \N__12494\,
            PADIN => \N__12493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8096\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__7514\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12486\,
            DIN => \N__12485\,
            DOUT => \N__12484\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12486\,
            PADOUT => \N__12485\,
            PADIN => \N__12484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4331\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__8924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12477\,
            DIN => \N__12476\,
            DOUT => \N__12475\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12477\,
            PADOUT => \N__12476\,
            PADIN => \N__12475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10751\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__5018\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12468\,
            DIN => \N__12467\,
            DOUT => \N__12466\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12468\,
            PADOUT => \N__12467\,
            PADIN => \N__12466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6248\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12459\,
            DIN => \N__12458\,
            DOUT => \N__12457\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12459\,
            PADOUT => \N__12458\,
            PADIN => \N__12457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10802\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__7736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12450\,
            DIN => \N__12449\,
            DOUT => \N__12448\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12450\,
            PADOUT => \N__12449\,
            PADIN => \N__12448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7703\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12441\,
            DIN => \N__12440\,
            DOUT => \N__12439\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12441\,
            PADOUT => \N__12440\,
            PADIN => \N__12439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4874\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__10649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12432\,
            DIN => \N__12431\,
            DOUT => \N__12430\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12432\,
            PADOUT => \N__12431\,
            PADIN => \N__12430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4445\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__5075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12423\,
            DIN => \N__12422\,
            DOUT => \N__12421\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12423\,
            PADOUT => \N__12422\,
            PADIN => \N__12421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12414\,
            DIN => \N__12413\,
            DOUT => \N__12412\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12414\,
            PADOUT => \N__12413\,
            PADIN => \N__12412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5159\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12405\,
            DIN => \N__12404\,
            DOUT => \N__12403\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12405\,
            PADOUT => \N__12404\,
            PADIN => \N__12403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5284\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12396\,
            DIN => \N__12395\,
            DOUT => \N__12394\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12396\,
            PADOUT => \N__12395\,
            PADIN => \N__12394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11369\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__5249\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12387\,
            DIN => \N__12386\,
            DOUT => \N__12385\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12387\,
            PADOUT => \N__12386\,
            PADIN => \N__12385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4139\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__11234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12378\,
            DIN => \N__12377\,
            DOUT => \N__12376\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12378\,
            PADOUT => \N__12377\,
            PADIN => \N__12376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4997\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__7760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12369\,
            DIN => \N__12368\,
            DOUT => \N__12367\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12369\,
            PADOUT => \N__12368\,
            PADIN => \N__12367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6665\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__7280\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12360\,
            DIN => \N__12359\,
            DOUT => \N__12358\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12360\,
            PADOUT => \N__12359\,
            PADIN => \N__12358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5495\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__5137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12351\,
            DIN => \N__12350\,
            DOUT => \N__12349\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12351\,
            PADOUT => \N__12350\,
            PADIN => \N__12349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12342\,
            DIN => \N__12341\,
            DOUT => \N__12340\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12342\,
            PADOUT => \N__12341\,
            PADIN => \N__12340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10781\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__5810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12333\,
            DIN => \N__12332\,
            DOUT => \N__12331\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12333\,
            PADOUT => \N__12332\,
            PADIN => \N__12331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11333\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__5216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12324\,
            DIN => \N__12323\,
            DOUT => \N__12322\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12324\,
            PADOUT => \N__12323\,
            PADIN => \N__12322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5483\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12315\,
            DIN => \N__12314\,
            DOUT => \N__12313\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12315\,
            PADOUT => \N__12314\,
            PADIN => \N__12313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4313\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__11435\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12306\,
            DIN => \N__12305\,
            DOUT => \N__12304\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12306\,
            PADOUT => \N__12305\,
            PADIN => \N__12304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4553\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__8603\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12297\,
            DIN => \N__12296\,
            DOUT => \N__12295\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12297\,
            PADOUT => \N__12296\,
            PADIN => \N__12295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12288\,
            DIN => \N__12287\,
            DOUT => \N__12286\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12288\,
            PADOUT => \N__12287\,
            PADIN => \N__12286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4271\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12279\,
            DIN => \N__12278\,
            DOUT => \N__12277\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12279\,
            PADOUT => \N__12278\,
            PADIN => \N__12277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11549\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__4970\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12270\,
            DIN => \N__12269\,
            DOUT => \N__12268\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12270\,
            PADOUT => \N__12269\,
            PADIN => \N__12268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10229\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__8633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12261\,
            DIN => \N__12260\,
            DOUT => \N__12259\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12261\,
            PADOUT => \N__12260\,
            PADIN => \N__12259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12252\,
            DIN => \N__12251\,
            DOUT => \N__12250\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12252\,
            PADOUT => \N__12251\,
            PADIN => \N__12250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4742\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__8858\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12243\,
            DIN => \N__12242\,
            DOUT => \N__12241\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12243\,
            PADOUT => \N__12242\,
            PADIN => \N__12241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12234\,
            DIN => \N__12233\,
            DOUT => \N__12232\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12234\,
            PADOUT => \N__12233\,
            PADIN => \N__12232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11606\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__9122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12225\,
            DIN => \N__12224\,
            DOUT => \N__12223\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12225\,
            PADOUT => \N__12224\,
            PADIN => \N__12223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4709\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__7817\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12216\,
            DIN => \N__12215\,
            DOUT => \N__12214\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12216\,
            PADOUT => \N__12215\,
            PADIN => \N__12214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4724\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__7913\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12207\,
            DIN => \N__12206\,
            DOUT => \N__12205\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12207\,
            PADOUT => \N__12206\,
            PADIN => \N__12205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10679\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__10289\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12198\,
            DIN => \N__12197\,
            DOUT => \N__12196\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12198\,
            PADOUT => \N__12197\,
            PADIN => \N__12196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12189\,
            DIN => \N__12188\,
            DOUT => \N__12187\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12189\,
            PADOUT => \N__12188\,
            PADIN => \N__12187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12180\,
            DIN => \N__12179\,
            DOUT => \N__12178\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12180\,
            PADOUT => \N__12179\,
            PADIN => \N__12178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11714\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__6632\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12171\,
            DIN => \N__12170\,
            DOUT => \N__12169\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12171\,
            PADOUT => \N__12170\,
            PADIN => \N__12169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4112\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__10610\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12162\,
            DIN => \N__12161\,
            DOUT => \N__12160\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12162\,
            PADOUT => \N__12161\,
            PADIN => \N__12160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10715\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__8117\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12153\,
            DIN => \N__12152\,
            DOUT => \N__12151\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12153\,
            PADOUT => \N__12152\,
            PADIN => \N__12151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12144\,
            DIN => \N__12143\,
            DOUT => \N__12142\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12144\,
            PADOUT => \N__12143\,
            PADIN => \N__12142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12135\,
            DIN => \N__12134\,
            DOUT => \N__12133\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12135\,
            PADOUT => \N__12134\,
            PADIN => \N__12133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4349\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__5381\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12126\,
            DIN => \N__12125\,
            DOUT => \N__12124\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12126\,
            PADOUT => \N__12125\,
            PADIN => \N__12124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12117\,
            DIN => \N__12116\,
            DOUT => \N__12115\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12117\,
            PADOUT => \N__12116\,
            PADIN => \N__12115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6133\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12108\,
            DIN => \N__12107\,
            DOUT => \N__12106\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12108\,
            PADOUT => \N__12107\,
            PADIN => \N__12106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8300\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__5183\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12099\,
            DIN => \N__12098\,
            DOUT => \N__12097\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12099\,
            PADOUT => \N__12098\,
            PADIN => \N__12097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4217\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__5996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12090\,
            DIN => \N__12089\,
            DOUT => \N__12088\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12090\,
            PADOUT => \N__12089\,
            PADIN => \N__12088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10556\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__4595\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12081\,
            DIN => \N__12080\,
            DOUT => \N__12079\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12081\,
            PADOUT => \N__12080\,
            PADIN => \N__12079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10523\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__7352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12072\,
            DIN => \N__12071\,
            DOUT => \N__12070\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12072\,
            PADOUT => \N__12071\,
            PADIN => \N__12070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4256\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__4531\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12063\,
            DIN => \N__12062\,
            DOUT => \N__12061\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12063\,
            PADOUT => \N__12062\,
            PADIN => \N__12061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4907\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__5846\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12054\,
            DIN => \N__12053\,
            DOUT => \N__12052\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12054\,
            PADOUT => \N__12053\,
            PADIN => \N__12052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10196\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__4664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12045\,
            DIN => \N__12044\,
            DOUT => \N__12043\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12045\,
            PADOUT => \N__12044\,
            PADIN => \N__12043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4163\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__10181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12036\,
            DIN => \N__12035\,
            DOUT => \N__12034\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12036\,
            PADOUT => \N__12035\,
            PADIN => \N__12034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4886\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__4367\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12027\,
            DIN => \N__12026\,
            DOUT => \N__12025\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12027\,
            PADOUT => \N__12026\,
            PADIN => \N__12025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4202\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__7577\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12018\,
            DIN => \N__12017\,
            DOUT => \N__12016\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12018\,
            PADOUT => \N__12017\,
            PADIN => \N__12016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7655\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__8321\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12009\,
            DIN => \N__12008\,
            DOUT => \N__12007\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12009\,
            PADOUT => \N__12008\,
            PADIN => \N__12007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12000\,
            DIN => \N__11999\,
            DOUT => \N__11998\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12000\,
            PADOUT => \N__11999\,
            PADIN => \N__11998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6557\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__6593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11991\,
            DIN => \N__11990\,
            DOUT => \N__11989\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11991\,
            PADOUT => \N__11990\,
            PADIN => \N__11989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11982\,
            DIN => \N__11981\,
            DOUT => \N__11980\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11982\,
            PADOUT => \N__11981\,
            PADIN => \N__11980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4100\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__11255\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11973\,
            DIN => \N__11972\,
            DOUT => \N__11971\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11973\,
            PADOUT => \N__11972\,
            PADIN => \N__11971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4928\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__4409\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11964\,
            DIN => \N__11963\,
            DOUT => \N__11962\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11964\,
            PADOUT => \N__11963\,
            PADIN => \N__11962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11955\,
            DIN => \N__11954\,
            DOUT => \N__11953\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11955\,
            PADOUT => \N__11954\,
            PADIN => \N__11953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11738\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__4808\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11946\,
            DIN => \N__11945\,
            DOUT => \N__11944\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11946\,
            PADOUT => \N__11945\,
            PADIN => \N__11944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10259\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__9050\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11937\,
            DIN => \N__11936\,
            DOUT => \N__11935\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11937\,
            PADOUT => \N__11936\,
            PADIN => \N__11935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8939\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__7433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11928\,
            DIN => \N__11927\,
            DOUT => \N__11926\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11928\,
            PADOUT => \N__11927\,
            PADIN => \N__11926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4574\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__5930\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11919\,
            DIN => \N__11918\,
            DOUT => \N__11917\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11919\,
            PADOUT => \N__11918\,
            PADIN => \N__11917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10580\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__6527\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11910\,
            DIN => \N__11909\,
            DOUT => \N__11908\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11910\,
            PADOUT => \N__11909\,
            PADIN => \N__11908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4856\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__11303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11901\,
            DIN => \N__11900\,
            DOUT => \N__11899\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11901\,
            PADOUT => \N__11900\,
            PADIN => \N__11899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11516\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__8711\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11892\,
            DIN => \N__11891\,
            DOUT => \N__11890\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11892\,
            PADOUT => \N__11891\,
            PADIN => \N__11890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6851\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11883\,
            DIN => \N__11882\,
            DOUT => \N__11881\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11883\,
            PADOUT => \N__11882\,
            PADIN => \N__11881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5039\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__5909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11874\,
            DIN => \N__11873\,
            DOUT => \N__11872\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11874\,
            PADOUT => \N__11873\,
            PADIN => \N__11872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11765\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__5537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11865\,
            DIN => \N__11864\,
            DOUT => \N__11863\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11865\,
            PADOUT => \N__11864\,
            PADIN => \N__11863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4082\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__10118\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11856\,
            DIN => \N__11855\,
            DOUT => \N__11854\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11856\,
            PADOUT => \N__11855\,
            PADIN => \N__11854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11847\,
            DIN => \N__11846\,
            DOUT => \N__11845\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11847\,
            PADOUT => \N__11846\,
            PADIN => \N__11845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11642\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__8480\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11838\,
            DIN => \N__11837\,
            DOUT => \N__11836\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11838\,
            PADOUT => \N__11837\,
            PADIN => \N__11836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5399\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__5309\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11829\,
            DIN => \N__11828\,
            DOUT => \N__11827\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11829\,
            PADOUT => \N__11828\,
            PADIN => \N__11827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__11402\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__7838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11820\,
            DIN => \N__11819\,
            DOUT => \N__11818\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11820\,
            PADOUT => \N__11819\,
            PADIN => \N__11818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5516\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__11486\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11811\,
            DIN => \N__11810\,
            DOUT => \N__11809\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11811\,
            PADOUT => \N__11810\,
            PADIN => \N__11809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10490\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__8399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11802\,
            DIN => \N__11801\,
            DOUT => \N__11800\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11802\,
            PADOUT => \N__11801\,
            PADIN => \N__11800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4793\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__10865\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2923\ : InMux
    port map (
            O => \N__11783\,
            I => \N__11780\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__2920\ : Sp12to4
    port map (
            O => \N__11774\,
            I => \N__11771\
        );

    \I__2919\ : Span12Mux_h
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__11768\,
            I => \READ_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__2917\ : IoInMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__2915\ : Span4Mux_s3_h
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__11753\,
            I => \N_221_i\
        );

    \I__2912\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11747\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__11747\,
            I => \N__11744\
        );

    \I__2910\ : Span12Mux_h
    port map (
            O => \N__11744\,
            I => \N__11741\
        );

    \I__2909\ : Odrv12
    port map (
            O => \N__11741\,
            I => \READ_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__2908\ : IoInMux
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__2906\ : Span12Mux_s8_h
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__2905\ : Odrv12
    port map (
            O => \N__11729\,
            I => \N_226_i\
        );

    \I__2904\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__2902\ : Span12Mux_s10_h
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__2901\ : Odrv12
    port map (
            O => \N__11717\,
            I => \READ_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__2900\ : IoInMux
    port map (
            O => \N__11714\,
            I => \N__11711\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__2898\ : Span4Mux_s3_h
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__2896\ : Sp12to4
    port map (
            O => \N__11702\,
            I => \N__11699\
        );

    \I__2895\ : Span12Mux_s9_h
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__2894\ : Span12Mux_v
    port map (
            O => \N__11696\,
            I => \N__11693\
        );

    \I__2893\ : Odrv12
    port map (
            O => \N__11693\,
            I => \N_229_i\
        );

    \I__2892\ : InMux
    port map (
            O => \N__11690\,
            I => \N__11687\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__11687\,
            I => \N__11684\
        );

    \I__2890\ : Span12Mux_s10_h
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__2889\ : Odrv12
    port map (
            O => \N__11681\,
            I => \READ_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__2888\ : IoInMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__2886\ : Span4Mux_s1_h
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__11666\,
            I => \N__11663\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__11660\,
            I => \N_214_i\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__2878\ : Sp12to4
    port map (
            O => \N__11648\,
            I => \N__11645\
        );

    \I__2877\ : Odrv12
    port map (
            O => \N__11645\,
            I => \READ_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__2876\ : IoInMux
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__2874\ : Span4Mux_s0_v
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__2871\ : Span4Mux_v
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__11624\,
            I => \N_217_i\
        );

    \I__2869\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2866\ : Sp12to4
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__11609\,
            I => \READ_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__2864\ : IoInMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__2862\ : Span4Mux_s2_h
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__2861\ : Span4Mux_h
    port map (
            O => \N__11597\,
            I => \N__11594\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__11594\,
            I => \N_213_i\
        );

    \I__2859\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__2857\ : Span12Mux_v
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__2856\ : Span12Mux_h
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__11579\,
            I => \READ_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__2854\ : IoInMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__2852\ : Span4Mux_s2_h
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__11564\,
            I => \N_228_i\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N__11555\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__11555\,
            I => \N__11552\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__11552\,
            I => \READ_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__2845\ : IoInMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__2843\ : IoSpan4Mux
    port map (
            O => \N__11543\,
            I => \N__11540\
        );

    \I__2842\ : IoSpan4Mux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__2841\ : Span4Mux_s1_h
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__11534\,
            I => \N_225_i\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__2836\ : Sp12to4
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__2835\ : Odrv12
    port map (
            O => \N__11519\,
            I => \READ_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__2834\ : IoInMux
    port map (
            O => \N__11516\,
            I => \N__11513\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__2832\ : Span12Mux_s7_v
    port map (
            O => \N__11510\,
            I => \N__11507\
        );

    \I__2831\ : Odrv12
    port map (
            O => \N__11507\,
            I => \N_208_i\
        );

    \I__2830\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__2826\ : Sp12to4
    port map (
            O => \N__11492\,
            I => \N__11489\
        );

    \I__2825\ : Odrv12
    port map (
            O => \N__11489\,
            I => \D_UM_040_in_7\
        );

    \I__2824\ : IoInMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11479\
        );

    \I__2822\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11476\
        );

    \I__2821\ : IoSpan4Mux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11476\,
            I => \N__11470\
        );

    \I__2819\ : Span4Mux_s3_h
    port map (
            O => \N__11473\,
            I => \N__11467\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__11470\,
            I => \N__11464\
        );

    \I__2817\ : Sp12to4
    port map (
            O => \N__11467\,
            I => \N__11461\
        );

    \I__2816\ : Sp12to4
    port map (
            O => \N__11464\,
            I => \N__11458\
        );

    \I__2815\ : Span12Mux_v
    port map (
            O => \N__11461\,
            I => \N__11455\
        );

    \I__2814\ : Span12Mux_v
    port map (
            O => \N__11458\,
            I => \N__11452\
        );

    \I__2813\ : Span12Mux_h
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__2812\ : Span12Mux_v
    port map (
            O => \N__11452\,
            I => \N__11446\
        );

    \I__2811\ : Span12Mux_h
    port map (
            O => \N__11449\,
            I => \N__11443\
        );

    \I__2810\ : Span12Mux_h
    port map (
            O => \N__11446\,
            I => \N__11440\
        );

    \I__2809\ : Odrv12
    port map (
            O => \N__11443\,
            I => \D_LL_040_in_7\
        );

    \I__2808\ : Odrv12
    port map (
            O => \N__11440\,
            I => \D_LL_040_in_7\
        );

    \I__2807\ : IoInMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11432\,
            I => \N__11429\
        );

    \I__2805\ : IoSpan4Mux
    port map (
            O => \N__11429\,
            I => \N__11426\
        );

    \I__2804\ : Span4Mux_s2_h
    port map (
            O => \N__11426\,
            I => \N__11423\
        );

    \I__2803\ : Span4Mux_h
    port map (
            O => \N__11423\,
            I => \N__11420\
        );

    \I__2802\ : Sp12to4
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__2801\ : Span12Mux_h
    port map (
            O => \N__11417\,
            I => \N__11414\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__11414\,
            I => \un1_D_UM_040_7\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11408\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__11408\,
            I => \N__11405\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__11405\,
            I => \READ_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__2796\ : IoInMux
    port map (
            O => \N__11402\,
            I => \N__11399\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11396\
        );

    \I__2794\ : Span4Mux_s1_h
    port map (
            O => \N__11396\,
            I => \N__11393\
        );

    \I__2793\ : Sp12to4
    port map (
            O => \N__11393\,
            I => \N__11390\
        );

    \I__2792\ : Span12Mux_s11_v
    port map (
            O => \N__11390\,
            I => \N__11387\
        );

    \I__2791\ : Odrv12
    port map (
            O => \N__11387\,
            I => \N_233_i\
        );

    \I__2790\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__2787\ : Sp12to4
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__11372\,
            I => \READ_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__2785\ : IoInMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__2783\ : Span4Mux_s3_h
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__2782\ : Sp12to4
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__2781\ : Span12Mux_s11_v
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__11354\,
            I => \N_235_i\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11345\
        );

    \I__2777\ : Span4Mux_v
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__2776\ : Sp12to4
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__2775\ : Span12Mux_h
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__11336\,
            I => \READ_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__2773\ : IoInMux
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11330\,
            I => \N__11327\
        );

    \I__2771\ : Span12Mux_s9_h
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__2770\ : Odrv12
    port map (
            O => \N__11324\,
            I => \N_222_i\
        );

    \I__2769\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11318\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__11306\,
            I => \D_UM_040_in_4\
        );

    \I__2763\ : IoInMux
    port map (
            O => \N__11303\,
            I => \N__11299\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__2759\ : Span4Mux_s2_h
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__11290\,
            I => \N__11284\
        );

    \I__2757\ : Span4Mux_v
    port map (
            O => \N__11287\,
            I => \N__11281\
        );

    \I__2756\ : Sp12to4
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__2755\ : Sp12to4
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__2754\ : Span12Mux_h
    port map (
            O => \N__11278\,
            I => \N__11272\
        );

    \I__2753\ : Span12Mux_h
    port map (
            O => \N__11275\,
            I => \N__11269\
        );

    \I__2752\ : Span12Mux_v
    port map (
            O => \N__11272\,
            I => \N__11266\
        );

    \I__2751\ : Span12Mux_h
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__2750\ : Span12Mux_v
    port map (
            O => \N__11266\,
            I => \N__11260\
        );

    \I__2749\ : Odrv12
    port map (
            O => \N__11263\,
            I => \D_LL_040_in_4\
        );

    \I__2748\ : Odrv12
    port map (
            O => \N__11260\,
            I => \D_LL_040_in_4\
        );

    \I__2747\ : IoInMux
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__2745\ : Span4Mux_s1_h
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__2744\ : Sp12to4
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__2743\ : Span12Mux_s7_v
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__2742\ : Span12Mux_h
    port map (
            O => \N__11240\,
            I => \N__11237\
        );

    \I__2741\ : Odrv12
    port map (
            O => \N__11237\,
            I => \un1_D_UM_040_4\
        );

    \I__2740\ : IoInMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__2738\ : IoSpan4Mux
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__2737\ : Span4Mux_s3_h
    port map (
            O => \N__11225\,
            I => \N__11221\
        );

    \I__2736\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11218\
        );

    \I__2735\ : Sp12to4
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11218\,
            I => \N__11212\
        );

    \I__2733\ : Span12Mux_v
    port map (
            O => \N__11215\,
            I => \N__11209\
        );

    \I__2732\ : Sp12to4
    port map (
            O => \N__11212\,
            I => \N__11206\
        );

    \I__2731\ : Span12Mux_h
    port map (
            O => \N__11209\,
            I => \N__11203\
        );

    \I__2730\ : Span12Mux_v
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__2729\ : Span12Mux_h
    port map (
            O => \N__11203\,
            I => \N__11197\
        );

    \I__2728\ : Span12Mux_v
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11197\,
            I => \D_LL_040_in_5\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11194\,
            I => \D_LL_040_in_5\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__2721\ : IoSpan4Mux
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__11174\,
            I => \D_UM_040_in_5\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11158\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11155\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11152\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11148\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11145\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11140\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11134\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11134\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11131\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11126\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11123\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11112\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11155\,
            I => \N__11112\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11108\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11105\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11148\,
            I => \N__11102\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11145\,
            I => \N__11099\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11094\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11094\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11140\,
            I => \N__11090\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11087\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11134\,
            I => \N__11083\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11131\,
            I => \N__11080\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11077\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11073\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11068\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11068\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11065\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11062\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11058\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11055\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11118\,
            I => \N__11052\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11049\
        );

    \I__2686\ : Span4Mux_v
    port map (
            O => \N__11112\,
            I => \N__11043\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11040\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__11108\,
            I => \N__11037\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11105\,
            I => \N__11034\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__11102\,
            I => \N__11031\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__11099\,
            I => \N__11026\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11094\,
            I => \N__11026\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11023\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__11090\,
            I => \N__11018\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11018\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11015\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__11083\,
            I => \N__11012\
        );

    \I__2674\ : Span4Mux_h
    port map (
            O => \N__11080\,
            I => \N__11007\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__11077\,
            I => \N__11007\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11004\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11073\,
            I => \N__11001\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__11068\,
            I => \N__10996\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11065\,
            I => \N__10996\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11062\,
            I => \N__10993\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11061\,
            I => \N__10990\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__10985\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__10985\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__10980\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11049\,
            I => \N__10980\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11048\,
            I => \N__10977\
        );

    \I__2661\ : InMux
    port map (
            O => \N__11047\,
            I => \N__10972\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11046\,
            I => \N__10972\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__11043\,
            I => \N__10967\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__10964\
        );

    \I__2657\ : Span4Mux_v
    port map (
            O => \N__11037\,
            I => \N__10959\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__11034\,
            I => \N__10959\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__11031\,
            I => \N__10954\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__11026\,
            I => \N__10954\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11023\,
            I => \N__10951\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__11018\,
            I => \N__10946\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__10946\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__11012\,
            I => \N__10939\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__11007\,
            I => \N__10939\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__10939\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__11001\,
            I => \N__10936\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__10996\,
            I => \N__10933\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__10993\,
            I => \N__10928\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10928\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__10985\,
            I => \N__10921\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__10980\,
            I => \N__10921\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10921\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10918\
        );

    \I__2639\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10915\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__10970\,
            I => \N__10912\
        );

    \I__2637\ : Sp12to4
    port map (
            O => \N__10967\,
            I => \N__10907\
        );

    \I__2636\ : Span12Mux_v
    port map (
            O => \N__10964\,
            I => \N__10907\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__10959\,
            I => \N__10900\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__10954\,
            I => \N__10900\
        );

    \I__2633\ : Span4Mux_v
    port map (
            O => \N__10951\,
            I => \N__10900\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__10946\,
            I => \N__10895\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__10939\,
            I => \N__10895\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__10936\,
            I => \N__10884\
        );

    \I__2629\ : Span4Mux_v
    port map (
            O => \N__10933\,
            I => \N__10884\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__10928\,
            I => \N__10884\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__10921\,
            I => \N__10884\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__10918\,
            I => \N__10884\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__10915\,
            I => \N__10881\
        );

    \I__2624\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10878\
        );

    \I__2623\ : Odrv12
    port map (
            O => \N__10907\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__10900\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__10895\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__10884\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__10881\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10878\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__2617\ : IoInMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__2615\ : Span12Mux_s6_v
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__2614\ : Span12Mux_h
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__10853\,
            I => \un1_D_UM_040_5\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__2609\ : Sp12to4
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__2608\ : Odrv12
    port map (
            O => \N__10838\,
            I => \READ_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__2607\ : IoInMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__2605\ : IoSpan4Mux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__2604\ : Span4Mux_s2_h
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__2603\ : Sp12to4
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__2602\ : Span12Mux_v
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__2601\ : Odrv12
    port map (
            O => \N__10817\,
            I => \N_230_i\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__10805\,
            I => \READ_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__2596\ : IoInMux
    port map (
            O => \N__10802\,
            I => \N__10799\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__2594\ : Odrv12
    port map (
            O => \N__10796\,
            I => \N_215_i\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__2591\ : Span12Mux_h
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__2590\ : Odrv12
    port map (
            O => \N__10784\,
            I => \READ_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__2589\ : IoInMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__2587\ : IoSpan4Mux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2586\ : Span4Mux_s2_v
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__10763\,
            I => \N_232_i\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__2580\ : Odrv12
    port map (
            O => \N__10754\,
            I => \READ_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__2579\ : IoInMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__2577\ : IoSpan4Mux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__2576\ : Span4Mux_s3_h
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2575\ : Span4Mux_v
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__10733\,
            I => \N_223_i\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__10718\,
            I => \READ_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__2567\ : IoInMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__2565\ : Span4Mux_s1_v
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__10697\,
            I => \N_205_i\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__10688\,
            I => \N__10685\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__10682\,
            I => \READ_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__2555\ : IoInMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__2553\ : Span4Mux_s3_v
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__2552\ : Sp12to4
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__2551\ : Span12Mux_s11_h
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__2550\ : Odrv12
    port map (
            O => \N__10664\,
            I => \N_212_i\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__2547\ : Span12Mux_h
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__10652\,
            I => \D_UM_040_in_2\
        );

    \I__2545\ : IoInMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2543\ : IoSpan4Mux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__2542\ : Span4Mux_s2_h
    port map (
            O => \N__10640\,
            I => \N__10636\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10633\
        );

    \I__2540\ : Sp12to4
    port map (
            O => \N__10636\,
            I => \N__10630\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10627\
        );

    \I__2538\ : Span12Mux_h
    port map (
            O => \N__10630\,
            I => \N__10624\
        );

    \I__2537\ : Span12Mux_v
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__2536\ : Span12Mux_h
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__2535\ : Span12Mux_v
    port map (
            O => \N__10621\,
            I => \N__10615\
        );

    \I__2534\ : Odrv12
    port map (
            O => \N__10618\,
            I => \D_LL_040_in_2\
        );

    \I__2533\ : Odrv12
    port map (
            O => \N__10615\,
            I => \D_LL_040_in_2\
        );

    \I__2532\ : IoInMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2530\ : Span4Mux_s2_h
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__2528\ : Sp12to4
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2526\ : Odrv12
    port map (
            O => \N__10592\,
            I => \un1_D_UM_040_2\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__10583\,
            I => \READ_CYCLE_ACTIVE_rep31_i_ess\
        );

    \I__2522\ : IoInMux
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__2520\ : Span12Mux_s10_h
    port map (
            O => \N__10574\,
            I => \N__10571\
        );

    \I__2519\ : Span12Mux_v
    port map (
            O => \N__10571\,
            I => \N__10568\
        );

    \I__2518\ : Odrv12
    port map (
            O => \N__10568\,
            I => \N_236_i\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10562\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__10562\,
            I => \N__10559\
        );

    \I__2515\ : Odrv12
    port map (
            O => \N__10559\,
            I => \READ_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__2514\ : IoInMux
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10553\,
            I => \N__10550\
        );

    \I__2512\ : IoSpan4Mux
    port map (
            O => \N__10550\,
            I => \N__10547\
        );

    \I__2511\ : Span4Mux_s2_h
    port map (
            O => \N__10547\,
            I => \N__10544\
        );

    \I__2510\ : Span4Mux_h
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__10541\,
            I => \N_227_i\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__10529\,
            I => \N__10526\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__10526\,
            I => \READ_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__2503\ : IoInMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10517\
        );

    \I__2501\ : Span4Mux_s0_v
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__2500\ : Sp12to4
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__2499\ : Span12Mux_s10_h
    port map (
            O => \N__10511\,
            I => \N__10508\
        );

    \I__2498\ : Odrv12
    port map (
            O => \N__10508\,
            I => \N_218_i\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10499\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__2494\ : Sp12to4
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__2493\ : Odrv12
    port map (
            O => \N__10493\,
            I => \READ_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__2492\ : IoInMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__2490\ : Span4Mux_s2_v
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__10475\,
            I => \N_209_i\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10468\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10468\,
            I => \N__10462\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10458\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__10462\,
            I => \N__10455\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10452\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__10458\,
            I => \N__10449\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__10455\,
            I => \N__10446\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10452\,
            I => \N__10443\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__10449\,
            I => \N__10440\
        );

    \I__2476\ : Sp12to4
    port map (
            O => \N__10446\,
            I => \N__10435\
        );

    \I__2475\ : Span12Mux_h
    port map (
            O => \N__10443\,
            I => \N__10435\
        );

    \I__2474\ : Span4Mux_h
    port map (
            O => \N__10440\,
            I => \N__10432\
        );

    \I__2473\ : Span12Mux_h
    port map (
            O => \N__10435\,
            I => \N__10429\
        );

    \I__2472\ : IoSpan4Mux
    port map (
            O => \N__10432\,
            I => \N__10426\
        );

    \I__2471\ : Odrv12
    port map (
            O => \N__10429\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__10426\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__10412\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10396\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10396\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10396\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10390\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10385\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10385\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10382\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10396\,
            I => \N__10376\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10371\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10371\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10368\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10360\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10360\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10360\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10357\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10354\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10351\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__10376\,
            I => \N__10343\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10371\,
            I => \N__10343\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10368\,
            I => \N__10343\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10340\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__10360\,
            I => \N__10331\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10357\,
            I => \N__10331\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10331\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10331\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10328\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__10343\,
            I => \N__10321\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10321\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__10331\,
            I => \N__10316\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10316\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10313\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__10326\,
            I => \N__10310\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__10321\,
            I => \N__10307\
        );

    \I__2432\ : Span4Mux_h
    port map (
            O => \N__10316\,
            I => \N__10304\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10301\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10298\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__10307\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__10304\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2427\ : Odrv12
    port map (
            O => \N__10301\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10298\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2425\ : IoInMux
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__2423\ : Span4Mux_s3_v
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__2421\ : Sp12to4
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__2420\ : Odrv12
    port map (
            O => \N__10274\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__2417\ : Span12Mux_h
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__2416\ : Odrv12
    port map (
            O => \N__10262\,
            I => \READ_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__2415\ : IoInMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__2413\ : IoSpan4Mux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__2412\ : Span4Mux_s0_h
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__2411\ : Sp12to4
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__2410\ : Odrv12
    port map (
            O => \N__10244\,
            I => \N_219_i\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10238\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__10235\,
            I => \N__10232\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__10232\,
            I => \READ_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__2405\ : IoInMux
    port map (
            O => \N__10229\,
            I => \N__10226\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__2403\ : Span4Mux_s1_h
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__2402\ : Sp12to4
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__2401\ : Span12Mux_s11_v
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__2400\ : Span12Mux_h
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__2399\ : Odrv12
    port map (
            O => \N__10211\,
            I => \N_220_i\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__2396\ : Span12Mux_h
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__2395\ : Odrv12
    port map (
            O => \N__10199\,
            I => \READ_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__2394\ : IoInMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__2392\ : Sp12to4
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__2391\ : Span12Mux_h
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__10184\,
            I => \N_234_i\
        );

    \I__2389\ : IoInMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__2387\ : IoSpan4Mux
    port map (
            O => \N__10175\,
            I => \N__10171\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10168\
        );

    \I__2385\ : IoSpan4Mux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__2383\ : Span4Mux_s2_h
    port map (
            O => \N__10165\,
            I => \N__10159\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__10162\,
            I => \N__10156\
        );

    \I__2381\ : Sp12to4
    port map (
            O => \N__10159\,
            I => \N__10153\
        );

    \I__2380\ : Sp12to4
    port map (
            O => \N__10156\,
            I => \N__10150\
        );

    \I__2379\ : Span12Mux_h
    port map (
            O => \N__10153\,
            I => \N__10147\
        );

    \I__2378\ : Span12Mux_h
    port map (
            O => \N__10150\,
            I => \N__10144\
        );

    \I__2377\ : Span12Mux_h
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__2376\ : Span12Mux_v
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__10141\,
            I => \D_LL_040_in_6\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__10138\,
            I => \D_LL_040_in_6\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__2371\ : Span4Mux_v
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__2370\ : Sp12to4
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__2369\ : Odrv12
    port map (
            O => \N__10121\,
            I => \D_UM_040_in_6\
        );

    \I__2368\ : IoInMux
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__2366\ : Span4Mux_s0_h
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2364\ : Sp12to4
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__2363\ : Span12Mux_v
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__2362\ : Span12Mux_h
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__2361\ : Odrv12
    port map (
            O => \N__10097\,
            I => \un1_D_UM_040_6\
        );

    \I__2360\ : IoInMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10087\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10078\
        );

    \I__2357\ : Span4Mux_s3_v
    port map (
            O => \N__10087\,
            I => \N__10074\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10066\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10066\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10066\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10059\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10059\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10059\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10052\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10052\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__10074\,
            I => \N__10044\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__10073\,
            I => \N__10035\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10032\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10059\,
            I => \N__10029\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10026\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10023\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10052\,
            I => \N__10020\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10015\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10015\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__10049\,
            I => \N__9996\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__10048\,
            I => \N__9993\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__10047\,
            I => \N__9989\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__10044\,
            I => \N__9985\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10043\,
            I => \N__9980\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10042\,
            I => \N__9980\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10041\,
            I => \N__9975\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10040\,
            I => \N__9975\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10039\,
            I => \N__9972\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10038\,
            I => \N__9969\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10035\,
            I => \N__9966\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__10032\,
            I => \N__9957\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__10029\,
            I => \N__9957\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10026\,
            I => \N__9957\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__9957\
        );

    \I__2324\ : Span4Mux_v
    port map (
            O => \N__10020\,
            I => \N__9952\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__9952\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10014\,
            I => \N__9949\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \N__9946\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__10012\,
            I => \N__9943\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__10011\,
            I => \N__9940\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10010\,
            I => \N__9931\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10009\,
            I => \N__9931\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10008\,
            I => \N__9931\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9914\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9914\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9914\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9914\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10003\,
            I => \N__9914\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10002\,
            I => \N__9914\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9914\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9914\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9901\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9901\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9901\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9901\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9901\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9901\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__9985\,
            I => \N__9884\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9884\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__9975\,
            I => \N__9884\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9972\,
            I => \N__9884\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9969\,
            I => \N__9884\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9881\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__9957\,
            I => \N__9874\
        );

    \I__2294\ : Span4Mux_h
    port map (
            O => \N__9952\,
            I => \N__9874\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9949\,
            I => \N__9874\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9865\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9865\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9865\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9865\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__9938\,
            I => \N__9861\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9931\,
            I => \N__9857\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9852\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9901\,
            I => \N__9852\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__9900\,
            I => \N__9847\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__9899\,
            I => \N__9843\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__9898\,
            I => \N__9831\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__9897\,
            I => \N__9827\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \N__9824\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__9895\,
            I => \N__9820\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__9884\,
            I => \N__9814\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__9881\,
            I => \N__9814\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__9874\,
            I => \N__9809\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9809\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9802\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9802\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9802\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__9857\,
            I => \N__9797\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9852\,
            I => \N__9797\
        );

    \I__2269\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9784\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9784\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9784\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9784\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9784\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9784\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9841\,
            I => \N__9767\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9767\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9767\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9767\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9767\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9767\
        );

    \I__2257\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9767\
        );

    \I__2256\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9767\
        );

    \I__2255\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9752\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9752\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9752\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9752\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9752\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9752\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9752\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__9814\,
            I => \N__9747\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9747\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9802\,
            I => \N__9744\
        );

    \I__2245\ : Sp12to4
    port map (
            O => \N__9797\,
            I => \N__9733\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9733\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9733\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9733\
        );

    \I__2241\ : Sp12to4
    port map (
            O => \N__9747\,
            I => \N__9733\
        );

    \I__2240\ : Span12Mux_v
    port map (
            O => \N__9744\,
            I => \N__9730\
        );

    \I__2239\ : Span12Mux_h
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__2238\ : Span12Mux_h
    port map (
            O => \N__9730\,
            I => \N__9724\
        );

    \I__2237\ : Odrv12
    port map (
            O => \N__9727\,
            I => \RnW_c\
        );

    \I__2236\ : Odrv12
    port map (
            O => \N__9724\,
            I => \RnW_c\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9710\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9710\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9710\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9710\,
            I => \N__9687\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9684\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9676\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9671\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9664\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9664\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9664\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9655\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9655\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9655\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9655\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9652\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9649\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9639\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9632\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9632\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9632\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9693\,
            I => \N__9627\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9627\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9622\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9622\
        );

    \I__2211\ : Span4Mux_v
    port map (
            O => \N__9687\,
            I => \N__9603\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9684\,
            I => \N__9603\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9598\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9598\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9591\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9591\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9591\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9676\,
            I => \N__9588\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9583\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9583\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9671\,
            I => \N__9564\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9559\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9559\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9554\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9649\,
            I => \N__9554\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9539\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9539\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9539\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9539\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9539\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9539\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9539\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9534\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9632\,
            I => \N__9534\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9531\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9528\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9515\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9515\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9515\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9515\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9515\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9515\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9498\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9498\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9498\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9498\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9498\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9498\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9498\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9498\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__9603\,
            I => \N__9487\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9487\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9487\
        );

    \I__2168\ : Span4Mux_h
    port map (
            O => \N__9588\,
            I => \N__9487\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9487\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9470\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9470\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9470\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9470\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9470\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9470\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9470\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9470\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9457\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9573\,
            I => \N__9457\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9457\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9457\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9457\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9457\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9454\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9451\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__9564\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__9559\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__9554\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9539\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__9534\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9531\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__9528\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9515\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9498\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__9487\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9470\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9457\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9454\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9451\,
            I => \U111_CYCLE_SM.N_44\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9413\
        );

    \I__2134\ : ClkMux
    port map (
            O => \N__9418\,
            I => \N__9317\
        );

    \I__2133\ : ClkMux
    port map (
            O => \N__9417\,
            I => \N__9317\
        );

    \I__2132\ : ClkMux
    port map (
            O => \N__9416\,
            I => \N__9317\
        );

    \I__2131\ : Glb2LocalMux
    port map (
            O => \N__9413\,
            I => \N__9317\
        );

    \I__2130\ : ClkMux
    port map (
            O => \N__9412\,
            I => \N__9317\
        );

    \I__2129\ : ClkMux
    port map (
            O => \N__9411\,
            I => \N__9317\
        );

    \I__2128\ : ClkMux
    port map (
            O => \N__9410\,
            I => \N__9317\
        );

    \I__2127\ : ClkMux
    port map (
            O => \N__9409\,
            I => \N__9317\
        );

    \I__2126\ : ClkMux
    port map (
            O => \N__9408\,
            I => \N__9317\
        );

    \I__2125\ : ClkMux
    port map (
            O => \N__9407\,
            I => \N__9317\
        );

    \I__2124\ : ClkMux
    port map (
            O => \N__9406\,
            I => \N__9317\
        );

    \I__2123\ : ClkMux
    port map (
            O => \N__9405\,
            I => \N__9317\
        );

    \I__2122\ : ClkMux
    port map (
            O => \N__9404\,
            I => \N__9317\
        );

    \I__2121\ : ClkMux
    port map (
            O => \N__9403\,
            I => \N__9317\
        );

    \I__2120\ : ClkMux
    port map (
            O => \N__9402\,
            I => \N__9317\
        );

    \I__2119\ : ClkMux
    port map (
            O => \N__9401\,
            I => \N__9317\
        );

    \I__2118\ : ClkMux
    port map (
            O => \N__9400\,
            I => \N__9317\
        );

    \I__2117\ : ClkMux
    port map (
            O => \N__9399\,
            I => \N__9317\
        );

    \I__2116\ : ClkMux
    port map (
            O => \N__9398\,
            I => \N__9317\
        );

    \I__2115\ : ClkMux
    port map (
            O => \N__9397\,
            I => \N__9317\
        );

    \I__2114\ : ClkMux
    port map (
            O => \N__9396\,
            I => \N__9317\
        );

    \I__2113\ : ClkMux
    port map (
            O => \N__9395\,
            I => \N__9317\
        );

    \I__2112\ : ClkMux
    port map (
            O => \N__9394\,
            I => \N__9317\
        );

    \I__2111\ : ClkMux
    port map (
            O => \N__9393\,
            I => \N__9317\
        );

    \I__2110\ : ClkMux
    port map (
            O => \N__9392\,
            I => \N__9317\
        );

    \I__2109\ : ClkMux
    port map (
            O => \N__9391\,
            I => \N__9317\
        );

    \I__2108\ : ClkMux
    port map (
            O => \N__9390\,
            I => \N__9317\
        );

    \I__2107\ : ClkMux
    port map (
            O => \N__9389\,
            I => \N__9317\
        );

    \I__2106\ : ClkMux
    port map (
            O => \N__9388\,
            I => \N__9317\
        );

    \I__2105\ : ClkMux
    port map (
            O => \N__9387\,
            I => \N__9317\
        );

    \I__2104\ : ClkMux
    port map (
            O => \N__9386\,
            I => \N__9317\
        );

    \I__2103\ : ClkMux
    port map (
            O => \N__9385\,
            I => \N__9317\
        );

    \I__2102\ : ClkMux
    port map (
            O => \N__9384\,
            I => \N__9317\
        );

    \I__2101\ : GlobalMux
    port map (
            O => \N__9317\,
            I => \CLK40\
        );

    \I__2100\ : CEMux
    port map (
            O => \N__9314\,
            I => \N__9257\
        );

    \I__2099\ : CEMux
    port map (
            O => \N__9313\,
            I => \N__9257\
        );

    \I__2098\ : CEMux
    port map (
            O => \N__9312\,
            I => \N__9257\
        );

    \I__2097\ : CEMux
    port map (
            O => \N__9311\,
            I => \N__9257\
        );

    \I__2096\ : CEMux
    port map (
            O => \N__9310\,
            I => \N__9257\
        );

    \I__2095\ : CEMux
    port map (
            O => \N__9309\,
            I => \N__9257\
        );

    \I__2094\ : CEMux
    port map (
            O => \N__9308\,
            I => \N__9257\
        );

    \I__2093\ : CEMux
    port map (
            O => \N__9307\,
            I => \N__9257\
        );

    \I__2092\ : CEMux
    port map (
            O => \N__9306\,
            I => \N__9257\
        );

    \I__2091\ : CEMux
    port map (
            O => \N__9305\,
            I => \N__9257\
        );

    \I__2090\ : CEMux
    port map (
            O => \N__9304\,
            I => \N__9257\
        );

    \I__2089\ : CEMux
    port map (
            O => \N__9303\,
            I => \N__9257\
        );

    \I__2088\ : CEMux
    port map (
            O => \N__9302\,
            I => \N__9257\
        );

    \I__2087\ : CEMux
    port map (
            O => \N__9301\,
            I => \N__9257\
        );

    \I__2086\ : CEMux
    port map (
            O => \N__9300\,
            I => \N__9257\
        );

    \I__2085\ : CEMux
    port map (
            O => \N__9299\,
            I => \N__9257\
        );

    \I__2084\ : CEMux
    port map (
            O => \N__9298\,
            I => \N__9257\
        );

    \I__2083\ : CEMux
    port map (
            O => \N__9297\,
            I => \N__9257\
        );

    \I__2082\ : CEMux
    port map (
            O => \N__9296\,
            I => \N__9257\
        );

    \I__2081\ : GlobalMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2080\ : gio2CtrlBuf
    port map (
            O => \N__9254\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9248\,
            I => \N__9221\
        );

    \I__2077\ : SRMux
    port map (
            O => \N__9247\,
            I => \N__9170\
        );

    \I__2076\ : SRMux
    port map (
            O => \N__9246\,
            I => \N__9170\
        );

    \I__2075\ : SRMux
    port map (
            O => \N__9245\,
            I => \N__9170\
        );

    \I__2074\ : SRMux
    port map (
            O => \N__9244\,
            I => \N__9170\
        );

    \I__2073\ : SRMux
    port map (
            O => \N__9243\,
            I => \N__9170\
        );

    \I__2072\ : SRMux
    port map (
            O => \N__9242\,
            I => \N__9170\
        );

    \I__2071\ : SRMux
    port map (
            O => \N__9241\,
            I => \N__9170\
        );

    \I__2070\ : SRMux
    port map (
            O => \N__9240\,
            I => \N__9170\
        );

    \I__2069\ : SRMux
    port map (
            O => \N__9239\,
            I => \N__9170\
        );

    \I__2068\ : SRMux
    port map (
            O => \N__9238\,
            I => \N__9170\
        );

    \I__2067\ : SRMux
    port map (
            O => \N__9237\,
            I => \N__9170\
        );

    \I__2066\ : SRMux
    port map (
            O => \N__9236\,
            I => \N__9170\
        );

    \I__2065\ : SRMux
    port map (
            O => \N__9235\,
            I => \N__9170\
        );

    \I__2064\ : SRMux
    port map (
            O => \N__9234\,
            I => \N__9170\
        );

    \I__2063\ : SRMux
    port map (
            O => \N__9233\,
            I => \N__9170\
        );

    \I__2062\ : SRMux
    port map (
            O => \N__9232\,
            I => \N__9170\
        );

    \I__2061\ : SRMux
    port map (
            O => \N__9231\,
            I => \N__9170\
        );

    \I__2060\ : SRMux
    port map (
            O => \N__9230\,
            I => \N__9170\
        );

    \I__2059\ : SRMux
    port map (
            O => \N__9229\,
            I => \N__9170\
        );

    \I__2058\ : SRMux
    port map (
            O => \N__9228\,
            I => \N__9170\
        );

    \I__2057\ : SRMux
    port map (
            O => \N__9227\,
            I => \N__9170\
        );

    \I__2056\ : SRMux
    port map (
            O => \N__9226\,
            I => \N__9170\
        );

    \I__2055\ : SRMux
    port map (
            O => \N__9225\,
            I => \N__9170\
        );

    \I__2054\ : SRMux
    port map (
            O => \N__9224\,
            I => \N__9170\
        );

    \I__2053\ : Glb2LocalMux
    port map (
            O => \N__9221\,
            I => \N__9170\
        );

    \I__2052\ : GlobalMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2051\ : gio2CtrlBuf
    port map (
            O => \N__9167\,
            I => \RESETn_c_i_g\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9161\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__9146\,
            I => \N__9141\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9138\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9135\
        );

    \I__2041\ : Sp12to4
    port map (
            O => \N__9141\,
            I => \N__9128\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9138\,
            I => \N__9128\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9135\,
            I => \N__9128\
        );

    \I__2038\ : Span12Mux_h
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__9125\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__2036\ : IoInMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__2034\ : IoSpan4Mux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2033\ : Span4Mux_s3_h
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__9104\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9098\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9091\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9087\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9084\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9081\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9078\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__9084\,
            I => \N__9075\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9081\,
            I => \N__9072\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__9078\,
            I => \N__9069\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9075\,
            I => \N__9064\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__9072\,
            I => \N__9064\
        );

    \I__2017\ : Sp12to4
    port map (
            O => \N__9069\,
            I => \N__9059\
        );

    \I__2016\ : Sp12to4
    port map (
            O => \N__9064\,
            I => \N__9059\
        );

    \I__2015\ : Span12Mux_h
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__2014\ : Span12Mux_v
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__9053\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__2012\ : IoInMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__2010\ : Span12Mux_s6_h
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__9041\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__9032\,
            I => \READ_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9021\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9018\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9015\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__9021\,
            I => \N__9012\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__9009\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9015\,
            I => \N__9006\
        );

    \I__1998\ : Sp12to4
    port map (
            O => \N__9012\,
            I => \N__9003\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__9009\,
            I => \N__9000\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__9006\,
            I => \N__8997\
        );

    \I__1995\ : Span12Mux_h
    port map (
            O => \N__9003\,
            I => \N__8994\
        );

    \I__1994\ : Sp12to4
    port map (
            O => \N__9000\,
            I => \N__8989\
        );

    \I__1993\ : Sp12to4
    port map (
            O => \N__8997\,
            I => \N__8989\
        );

    \I__1992\ : Span12Mux_v
    port map (
            O => \N__8994\,
            I => \N__8986\
        );

    \I__1991\ : Span12Mux_h
    port map (
            O => \N__8989\,
            I => \N__8983\
        );

    \I__1990\ : Odrv12
    port map (
            O => \N__8986\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__8983\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8975\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__1984\ : Span4Mux_s2_h
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__1983\ : Sp12to4
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__1982\ : Span12Mux_v
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__1981\ : Span12Mux_h
    port map (
            O => \N__8957\,
            I => \N__8954\
        );

    \I__1980\ : Odrv12
    port map (
            O => \N__8954\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__8942\,
            I => \READ_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__1975\ : IoInMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1973\ : Span12Mux_s2_h
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1972\ : Span12Mux_h
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1971\ : Odrv12
    port map (
            O => \N__8927\,
            I => \N_216_i\
        );

    \I__1970\ : IoInMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8921\,
            I => \N__8917\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__1967\ : Span4Mux_s3_h
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__1965\ : Span4Mux_h
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__1963\ : Sp12to4
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1962\ : Sp12to4
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__1961\ : Span12Mux_v
    port map (
            O => \N__8899\,
            I => \N__8893\
        );

    \I__1960\ : Span12Mux_v
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1959\ : Span12Mux_h
    port map (
            O => \N__8893\,
            I => \N__8885\
        );

    \I__1958\ : Span12Mux_v
    port map (
            O => \N__8890\,
            I => \N__8885\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8882\,
            I => \D_LM_040_in_1\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__1951\ : Sp12to4
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__1950\ : Span12Mux_h
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__1949\ : Odrv12
    port map (
            O => \N__8861\,
            I => \D_UU_040_in_1\
        );

    \I__1948\ : IoInMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8855\,
            I => \N__8852\
        );

    \I__1946\ : Span4Mux_s1_h
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__8837\,
            I => \un1_D_UU_040_1\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__8828\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8820\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8817\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8814\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8820\,
            I => \N__8811\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8808\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8805\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__8811\,
            I => \N__8800\
        );

    \I__1930\ : Span4Mux_v
    port map (
            O => \N__8808\,
            I => \N__8800\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__8805\,
            I => \N__8797\
        );

    \I__1928\ : Sp12to4
    port map (
            O => \N__8800\,
            I => \N__8792\
        );

    \I__1927\ : Sp12to4
    port map (
            O => \N__8797\,
            I => \N__8792\
        );

    \I__1926\ : Span12Mux_h
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__8789\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1924\ : IoInMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__1922\ : Span12Mux_s8_v
    port map (
            O => \N__8780\,
            I => \N__8777\
        );

    \I__1921\ : Odrv12
    port map (
            O => \N__8777\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__8768\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8757\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8754\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8751\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__8757\,
            I => \N__8748\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8754\,
            I => \N__8745\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8742\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__8748\,
            I => \N__8739\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__8745\,
            I => \N__8736\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__8742\,
            I => \N__8733\
        );

    \I__1907\ : Sp12to4
    port map (
            O => \N__8739\,
            I => \N__8728\
        );

    \I__1906\ : Sp12to4
    port map (
            O => \N__8736\,
            I => \N__8728\
        );

    \I__1905\ : Sp12to4
    port map (
            O => \N__8733\,
            I => \N__8725\
        );

    \I__1904\ : Span12Mux_h
    port map (
            O => \N__8728\,
            I => \N__8722\
        );

    \I__1903\ : Span12Mux_v
    port map (
            O => \N__8725\,
            I => \N__8719\
        );

    \I__1902\ : Span12Mux_v
    port map (
            O => \N__8722\,
            I => \N__8714\
        );

    \I__1901\ : Span12Mux_h
    port map (
            O => \N__8719\,
            I => \N__8714\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__8714\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1899\ : IoInMux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1897\ : IoSpan4Mux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__1896\ : IoSpan4Mux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1895\ : Span4Mux_s3_v
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__8690\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8683\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8679\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8676\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8673\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8679\,
            I => \N__8670\
        );

    \I__1886\ : Span12Mux_v
    port map (
            O => \N__8676\,
            I => \N__8665\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8665\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__8670\,
            I => \N__8662\
        );

    \I__1883\ : Span12Mux_v
    port map (
            O => \N__8665\,
            I => \N__8659\
        );

    \I__1882\ : Sp12to4
    port map (
            O => \N__8662\,
            I => \N__8656\
        );

    \I__1881\ : Span12Mux_h
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__1880\ : Span12Mux_h
    port map (
            O => \N__8656\,
            I => \N__8650\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__8653\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__8650\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__8636\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1873\ : IoInMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1871\ : Span12Mux_s3_h
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1870\ : Span12Mux_h
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1869\ : Odrv12
    port map (
            O => \N__8621\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1866\ : Span12Mux_s7_v
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1865\ : Span12Mux_h
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1864\ : Odrv12
    port map (
            O => \N__8606\,
            I => \D_UU_040_in_7\
        );

    \I__1863\ : IoInMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1861\ : IoSpan4Mux
    port map (
            O => \N__8597\,
            I => \N__8593\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8590\
        );

    \I__1859\ : Span4Mux_s2_h
    port map (
            O => \N__8593\,
            I => \N__8587\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8590\,
            I => \N__8584\
        );

    \I__1857\ : Sp12to4
    port map (
            O => \N__8587\,
            I => \N__8581\
        );

    \I__1856\ : Sp12to4
    port map (
            O => \N__8584\,
            I => \N__8578\
        );

    \I__1855\ : Span12Mux_h
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__1854\ : Span12Mux_s9_v
    port map (
            O => \N__8578\,
            I => \N__8572\
        );

    \I__1853\ : Span12Mux_h
    port map (
            O => \N__8575\,
            I => \N__8569\
        );

    \I__1852\ : Span12Mux_h
    port map (
            O => \N__8572\,
            I => \N__8566\
        );

    \I__1851\ : Odrv12
    port map (
            O => \N__8569\,
            I => \D_LM_040_in_7\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__8566\,
            I => \D_LM_040_in_7\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1847\ : Span4Mux_s2_v
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1844\ : Span12Mux_s11_h
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1843\ : Odrv12
    port map (
            O => \N__8543\,
            I => \un1_D_UU_040_7\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__8531\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8524\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8524\,
            I => \N__8518\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8514\
        );

    \I__1834\ : Span4Mux_h
    port map (
            O => \N__8518\,
            I => \N__8511\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8508\
        );

    \I__1832\ : Sp12to4
    port map (
            O => \N__8514\,
            I => \N__8505\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__8511\,
            I => \N__8500\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8500\
        );

    \I__1829\ : Span12Mux_v
    port map (
            O => \N__8505\,
            I => \N__8497\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8500\,
            I => \N__8494\
        );

    \I__1827\ : Span12Mux_h
    port map (
            O => \N__8497\,
            I => \N__8491\
        );

    \I__1826\ : Sp12to4
    port map (
            O => \N__8494\,
            I => \N__8488\
        );

    \I__1825\ : Span12Mux_v
    port map (
            O => \N__8491\,
            I => \N__8483\
        );

    \I__1824\ : Span12Mux_h
    port map (
            O => \N__8488\,
            I => \N__8483\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__8483\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1819\ : IoSpan4Mux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1818\ : IoSpan4Mux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1817\ : Span4Mux_s2_v
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__8459\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8449\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8445\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8449\,
            I => \N__8442\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8439\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8445\,
            I => \N__8436\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__8442\,
            I => \N__8431\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8439\,
            I => \N__8431\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8436\,
            I => \N__8428\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__8431\,
            I => \N__8425\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__1803\ : Sp12to4
    port map (
            O => \N__8425\,
            I => \N__8419\
        );

    \I__1802\ : Sp12to4
    port map (
            O => \N__8422\,
            I => \N__8416\
        );

    \I__1801\ : Span12Mux_h
    port map (
            O => \N__8419\,
            I => \N__8413\
        );

    \I__1800\ : Odrv12
    port map (
            O => \N__8416\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1799\ : Odrv12
    port map (
            O => \N__8413\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1796\ : Odrv12
    port map (
            O => \N__8402\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1795\ : IoInMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__1793\ : Span4Mux_s3_v
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1792\ : Span4Mux_h
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__8384\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__8375\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8368\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8365\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8362\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8359\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__8362\,
            I => \N__8356\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__8359\,
            I => \N__8353\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__8356\,
            I => \N__8349\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8353\,
            I => \N__8346\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8343\
        );

    \I__1777\ : Span12Mux_v
    port map (
            O => \N__8349\,
            I => \N__8340\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__8346\,
            I => \N__8337\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8334\
        );

    \I__1774\ : Span12Mux_h
    port map (
            O => \N__8340\,
            I => \N__8331\
        );

    \I__1773\ : Sp12to4
    port map (
            O => \N__8337\,
            I => \N__8326\
        );

    \I__1772\ : Span12Mux_v
    port map (
            O => \N__8334\,
            I => \N__8326\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8331\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__8326\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1769\ : IoInMux
    port map (
            O => \N__8321\,
            I => \N__8318\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8318\,
            I => \N__8315\
        );

    \I__1767\ : Span4Mux_s3_v
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__1766\ : Span4Mux_h
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__1764\ : Span4Mux_h
    port map (
            O => \N__8306\,
            I => \N__8303\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__8303\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1762\ : IoInMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1760\ : IoSpan4Mux
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1759\ : Span4Mux_s3_h
    port map (
            O => \N__8291\,
            I => \N__8288\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__1757\ : Span12Mux_h
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__8282\,
            I => \N_224_i\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8273\,
            I => \N__8268\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8265\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8262\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__8268\,
            I => \N__8255\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8255\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8255\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__8252\,
            I => \N__8249\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__8246\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8240\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1741\ : CEMux
    port map (
            O => \N__8237\,
            I => \N__8231\
        );

    \I__1740\ : CEMux
    port map (
            O => \N__8236\,
            I => \N__8228\
        );

    \I__1739\ : CEMux
    port map (
            O => \N__8235\,
            I => \N__8225\
        );

    \I__1738\ : CEMux
    port map (
            O => \N__8234\,
            I => \N__8222\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8231\,
            I => \U111_CYCLE_SM.N_40_i_0\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8228\,
            I => \U111_CYCLE_SM.N_40_i_0\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8225\,
            I => \U111_CYCLE_SM.N_40_i_0\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8222\,
            I => \U111_CYCLE_SM.N_40_i_0\
        );

    \I__1733\ : SRMux
    port map (
            O => \N__8213\,
            I => \N__8208\
        );

    \I__1732\ : SRMux
    port map (
            O => \N__8212\,
            I => \N__8205\
        );

    \I__1731\ : SRMux
    port map (
            O => \N__8211\,
            I => \N__8202\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8198\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8205\,
            I => \N__8195\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8192\
        );

    \I__1727\ : SRMux
    port map (
            O => \N__8201\,
            I => \N__8189\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__8198\,
            I => \N__8184\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__8195\,
            I => \N__8184\
        );

    \I__1724\ : Span4Mux_h
    port map (
            O => \N__8192\,
            I => \N__8179\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8189\,
            I => \N__8179\
        );

    \I__1722\ : Span4Mux_h
    port map (
            O => \N__8184\,
            I => \N__8176\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__8179\,
            I => \N__8173\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__8176\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__8173\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8165\,
            I => \N__8160\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8157\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8154\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8160\,
            I => \N__8151\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8146\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8154\,
            I => \N__8146\
        );

    \I__1711\ : Sp12to4
    port map (
            O => \N__8151\,
            I => \N__8143\
        );

    \I__1710\ : Sp12to4
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1709\ : Span12Mux_h
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1708\ : Span12Mux_v
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1707\ : Span12Mux_v
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1706\ : Span12Mux_h
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__8131\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1704\ : Odrv12
    port map (
            O => \N__8128\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8120\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8120\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1701\ : IoInMux
    port map (
            O => \N__8117\,
            I => \N__8114\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8114\,
            I => \N__8111\
        );

    \I__1699\ : Span4Mux_s2_v
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1697\ : Sp12to4
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1696\ : Span12Mux_s11_v
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__8099\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1694\ : IoInMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1692\ : Span4Mux_s3_h
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1690\ : Sp12to4
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1689\ : Span12Mux_s8_v
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__8078\,
            I => \N_206_i\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__8069\,
            I => \N__8065\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__8068\,
            I => \N__8062\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__8065\,
            I => \N__8059\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8056\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__8059\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8056\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8046\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8050\,
            I => \N__8043\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8040\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N__8037\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8034\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8030\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__8037\,
            I => \N__8025\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8025\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8022\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__8030\,
            I => \N__8019\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__8025\,
            I => \N__8016\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__8012\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__8019\,
            I => \N__8009\
        );

    \I__1666\ : Sp12to4
    port map (
            O => \N__8016\,
            I => \N__8006\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8003\
        );

    \I__1664\ : Span12Mux_v
    port map (
            O => \N__8012\,
            I => \N__7996\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__8009\,
            I => \N__7996\
        );

    \I__1662\ : Span12Mux_h
    port map (
            O => \N__8006\,
            I => \N__7996\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8003\,
            I => \N__7993\
        );

    \I__1660\ : Span12Mux_v
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7987\
        );

    \I__1658\ : Odrv12
    port map (
            O => \N__7990\,
            I => \LBENn_c\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__7987\,
            I => \LBENn_c\
        );

    \I__1656\ : IoInMux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1654\ : Span4Mux_s3_v
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__7970\,
            I => \TAn_1_i\
        );

    \I__1651\ : IoInMux
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1649\ : Span4Mux_s1_h
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1648\ : Sp12to4
    port map (
            O => \N__7958\,
            I => \N__7954\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7951\
        );

    \I__1646\ : Span12Mux_v
    port map (
            O => \N__7954\,
            I => \N__7948\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7945\
        );

    \I__1644\ : Span12Mux_h
    port map (
            O => \N__7948\,
            I => \N__7942\
        );

    \I__1643\ : Span12Mux_h
    port map (
            O => \N__7945\,
            I => \N__7939\
        );

    \I__1642\ : Span12Mux_h
    port map (
            O => \N__7942\,
            I => \N__7934\
        );

    \I__1641\ : Span12Mux_v
    port map (
            O => \N__7939\,
            I => \N__7934\
        );

    \I__1640\ : Odrv12
    port map (
            O => \N__7934\,
            I => \D_LM_040_in_4\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1636\ : Sp12to4
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__7916\,
            I => \D_UU_040_in_4\
        );

    \I__1633\ : IoInMux
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1631\ : Span4Mux_s2_v
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1629\ : Sp12to4
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1628\ : Odrv12
    port map (
            O => \N__7898\,
            I => \un1_D_UU_040_4\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1624\ : Sp12to4
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1623\ : Span12Mux_h
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__7880\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__1621\ : IoInMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1619\ : Span4Mux_s3_h
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__7868\,
            I => \N__7865\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__7865\,
            I => \N__7862\
        );

    \I__1616\ : Span12Mux_h
    port map (
            O => \N__7862\,
            I => \N__7859\
        );

    \I__1615\ : Odrv12
    port map (
            O => \N__7859\,
            I => \un2_D_LL_AMIGA_1\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7853\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1611\ : Sp12to4
    port map (
            O => \N__7847\,
            I => \N__7844\
        );

    \I__1610\ : Span12Mux_h
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__7841\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__1608\ : IoInMux
    port map (
            O => \N__7838\,
            I => \N__7835\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__1606\ : IoSpan4Mux
    port map (
            O => \N__7832\,
            I => \N__7829\
        );

    \I__1605\ : Span4Mux_s2_h
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1604\ : Sp12to4
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1603\ : Span12Mux_h
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__7820\,
            I => \un2_D_LL_AMIGA_4\
        );

    \I__1601\ : IoInMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7814\,
            I => \N__7810\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7807\
        );

    \I__1598\ : IoSpan4Mux
    port map (
            O => \N__7810\,
            I => \N__7804\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7807\,
            I => \N__7801\
        );

    \I__1596\ : Span4Mux_s2_h
    port map (
            O => \N__7804\,
            I => \N__7798\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7801\,
            I => \N__7795\
        );

    \I__1594\ : Sp12to4
    port map (
            O => \N__7798\,
            I => \N__7792\
        );

    \I__1593\ : Sp12to4
    port map (
            O => \N__7795\,
            I => \N__7789\
        );

    \I__1592\ : Span12Mux_h
    port map (
            O => \N__7792\,
            I => \N__7786\
        );

    \I__1591\ : Span12Mux_v
    port map (
            O => \N__7789\,
            I => \N__7783\
        );

    \I__1590\ : Span12Mux_h
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__1589\ : Span12Mux_h
    port map (
            O => \N__7783\,
            I => \N__7777\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__7780\,
            I => \D_LL_040_in_0\
        );

    \I__1587\ : Odrv12
    port map (
            O => \N__7777\,
            I => \D_LL_040_in_0\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7769\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__1584\ : Span12Mux_h
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1583\ : Odrv12
    port map (
            O => \N__7763\,
            I => \D_UM_040_in_0\
        );

    \I__1582\ : IoInMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1580\ : IoSpan4Mux
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1579\ : Span4Mux_s2_h
    port map (
            O => \N__7751\,
            I => \N__7748\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__7748\,
            I => \N__7745\
        );

    \I__1577\ : Span4Mux_h
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__7742\,
            I => \N__7739\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__7739\,
            I => \un1_D_UM_040_0\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7733\,
            I => \N__7730\
        );

    \I__1572\ : IoSpan4Mux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1571\ : Span4Mux_s3_h
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1570\ : Span4Mux_h
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__7718\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__1565\ : Glb2LocalMux
    port map (
            O => \N__7709\,
            I => \N__7706\
        );

    \I__1564\ : GlobalMux
    port map (
            O => \N__7706\,
            I => \CLK80\
        );

    \I__1563\ : IoInMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7696\
        );

    \I__1561\ : IoInMux
    port map (
            O => \N__7699\,
            I => \N__7693\
        );

    \I__1560\ : Span4Mux_s0_v
    port map (
            O => \N__7696\,
            I => \N__7690\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7693\,
            I => \N__7687\
        );

    \I__1558\ : Sp12to4
    port map (
            O => \N__7690\,
            I => \N__7684\
        );

    \I__1557\ : Span4Mux_s3_h
    port map (
            O => \N__7687\,
            I => \N__7681\
        );

    \I__1556\ : Span12Mux_h
    port map (
            O => \N__7684\,
            I => \N__7678\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7681\,
            I => \N__7675\
        );

    \I__1554\ : Span12Mux_v
    port map (
            O => \N__7678\,
            I => \N__7672\
        );

    \I__1553\ : Sp12to4
    port map (
            O => \N__7675\,
            I => \N__7669\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__7672\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7669\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__7658\,
            I => \READ_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__1547\ : IoInMux
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1545\ : IoSpan4Mux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1544\ : Span4Mux_s0_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1543\ : Sp12to4
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1542\ : Span12Mux_s11_v
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__7637\,
            I => \N_210_i\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1537\ : Sp12to4
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__1536\ : Span12Mux_h
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1535\ : Span12Mux_v
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__7616\,
            I => \D_UM_040_in_1\
        );

    \I__1533\ : IoInMux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1531\ : Span4Mux_s3_h
    port map (
            O => \N__7607\,
            I => \N__7603\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1529\ : Sp12to4
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7600\,
            I => \N__7594\
        );

    \I__1527\ : Span12Mux_v
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__1526\ : Span12Mux_v
    port map (
            O => \N__7594\,
            I => \N__7588\
        );

    \I__1525\ : Span12Mux_h
    port map (
            O => \N__7591\,
            I => \N__7583\
        );

    \I__1524\ : Span12Mux_v
    port map (
            O => \N__7588\,
            I => \N__7583\
        );

    \I__1523\ : Span12Mux_h
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__7580\,
            I => \D_LL_040_in_1\
        );

    \I__1521\ : IoInMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1519\ : Span4Mux_s3_h
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1518\ : Span4Mux_h
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__7559\,
            I => \un1_D_UM_040_1\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__7550\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7542\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7539\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7536\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7531\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7539\,
            I => \N__7531\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7536\,
            I => \N__7528\
        );

    \I__1505\ : Span12Mux_v
    port map (
            O => \N__7531\,
            I => \N__7525\
        );

    \I__1504\ : Span12Mux_v
    port map (
            O => \N__7528\,
            I => \N__7522\
        );

    \I__1503\ : Span12Mux_h
    port map (
            O => \N__7525\,
            I => \N__7519\
        );

    \I__1502\ : Odrv12
    port map (
            O => \N__7522\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__7519\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1500\ : IoInMux
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__1498\ : IoSpan4Mux
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__1497\ : Span4Mux_s3_h
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__1495\ : Sp12to4
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__1494\ : Span12Mux_h
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__1493\ : Odrv12
    port map (
            O => \N__7493\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7482\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7479\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7485\,
            I => \N__7476\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__7482\,
            I => \N__7471\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7479\,
            I => \N__7471\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7476\,
            I => \N__7468\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__7471\,
            I => \N__7465\
        );

    \I__1484\ : Span12Mux_v
    port map (
            O => \N__7468\,
            I => \N__7462\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7465\,
            I => \N__7459\
        );

    \I__1482\ : Span12Mux_h
    port map (
            O => \N__7462\,
            I => \N__7456\
        );

    \I__1481\ : Span4Mux_h
    port map (
            O => \N__7459\,
            I => \N__7453\
        );

    \I__1480\ : Span12Mux_v
    port map (
            O => \N__7456\,
            I => \N__7450\
        );

    \I__1479\ : Sp12to4
    port map (
            O => \N__7453\,
            I => \N__7447\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__7450\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1477\ : Odrv12
    port map (
            O => \N__7447\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__7436\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1473\ : IoInMux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__1471\ : Span4Mux_s2_h
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__7424\,
            I => \N__7421\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__1468\ : Sp12to4
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1467\ : Span12Mux_h
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1466\ : Odrv12
    port map (
            O => \N__7412\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7405\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7405\,
            I => \N__7398\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7402\,
            I => \N__7395\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7392\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7398\,
            I => \N__7389\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__7395\,
            I => \N__7384\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7384\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__7389\,
            I => \N__7381\
        );

    \I__1456\ : Sp12to4
    port map (
            O => \N__7384\,
            I => \N__7378\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__7381\,
            I => \N__7375\
        );

    \I__1454\ : Span12Mux_v
    port map (
            O => \N__7378\,
            I => \N__7372\
        );

    \I__1453\ : Span12Mux_v
    port map (
            O => \N__7375\,
            I => \N__7367\
        );

    \I__1452\ : Span12Mux_h
    port map (
            O => \N__7372\,
            I => \N__7367\
        );

    \I__1451\ : Odrv12
    port map (
            O => \N__7367\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__7355\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1446\ : IoInMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1444\ : Span4Mux_s2_v
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1443\ : Span4Mux_h
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1442\ : Span4Mux_h
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1441\ : Sp12to4
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__1440\ : Span12Mux_s8_v
    port map (
            O => \N__7334\,
            I => \N__7331\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__7331\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7325\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__1436\ : Odrv12
    port map (
            O => \N__7322\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7314\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7311\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7308\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7314\,
            I => \N__7305\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7302\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7299\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__7305\,
            I => \N__7296\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__7302\,
            I => \N__7291\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__7299\,
            I => \N__7291\
        );

    \I__1426\ : Sp12to4
    port map (
            O => \N__7296\,
            I => \N__7286\
        );

    \I__1425\ : Sp12to4
    port map (
            O => \N__7291\,
            I => \N__7286\
        );

    \I__1424\ : Span12Mux_h
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1423\ : Odrv12
    port map (
            O => \N__7283\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1422\ : IoInMux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1420\ : Span4Mux_s2_v
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1419\ : Sp12to4
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1418\ : Span12Mux_h
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1417\ : Odrv12
    port map (
            O => \N__7265\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__7256\,
            I => \READ_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \U111_CYCLE_SM.N_55_cascade_\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7243\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__7243\,
            I => \U111_CYCLE_SM.N_73\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7240\,
            I => \U111_CYCLE_SM.N_73\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7229\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7226\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7223\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7220\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7217\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7226\,
            I => \N__7212\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7212\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7220\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__7217\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__7212\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1397\ : IoInMux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1395\ : Span4Mux_s1_v
    port map (
            O => \N__7199\,
            I => \N__7194\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__7198\,
            I => \N__7190\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__7197\,
            I => \N__7185\
        );

    \I__1392\ : Span4Mux_v
    port map (
            O => \N__7194\,
            I => \N__7181\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7178\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7171\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7171\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7171\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7166\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7166\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7181\,
            I => \N__7163\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7178\,
            I => \N__7156\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7171\,
            I => \N__7156\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7166\,
            I => \N__7156\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__7163\,
            I => \N__7150\
        );

    \I__1380\ : Span4Mux_v
    port map (
            O => \N__7156\,
            I => \N__7150\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__7155\,
            I => \N__7147\
        );

    \I__1378\ : Sp12to4
    port map (
            O => \N__7150\,
            I => \N__7143\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7138\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7138\
        );

    \I__1375\ : Span12Mux_h
    port map (
            O => \N__7143\,
            I => \N__7133\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7138\,
            I => \N__7133\
        );

    \I__1373\ : Span12Mux_v
    port map (
            O => \N__7133\,
            I => \N__7130\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__7130\,
            I => \TACKn_in\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7127\,
            I => \N__7120\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7117\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7108\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7108\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7108\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7108\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7117\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7108\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7103\,
            I => \U111_CYCLE_SM.N_57_cascade_\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7097\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__7085\,
            I => \N__7078\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7075\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7083\,
            I => \N__7072\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7069\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7066\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__7078\,
            I => \N__7063\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7072\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7069\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7066\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7063\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7048\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__7040\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7045\,
            I => \N__7040\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__7040\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7031\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7028\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7025\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7022\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7031\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7028\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7025\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7022\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1330\ : Sp12to4
    port map (
            O => \N__7004\,
            I => \N__7000\
        );

    \I__1329\ : IoInMux
    port map (
            O => \N__7003\,
            I => \N__6997\
        );

    \I__1328\ : Span12Mux_h
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6991\
        );

    \I__1326\ : Span12Mux_v
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__1325\ : IoSpan4Mux
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__1324\ : Odrv12
    port map (
            O => \N__6988\,
            I => \TBIn_c\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6985\,
            I => \TBIn_c\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6972\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6969\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6972\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6955\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6952\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6955\,
            I => \U111_CYCLE_SM.N_42\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6952\,
            I => \U111_CYCLE_SM.N_42\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__6947\,
            I => \U111_CYCLE_SM.N_46_cascade_\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6936\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6927\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6927\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6927\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6927\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6924\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6936\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6927\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6924\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6910\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6910\,
            I => \N__6904\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6907\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__6904\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6896\,
            I => \U111_CYCLE_SM.N_39\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6888\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6883\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6883\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6888\,
            I => \U111_CYCLE_SM.N_40\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6883\,
            I => \U111_CYCLE_SM.N_40\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__6878\,
            I => \U111_CYCLE_SM.N_40_cascade_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6871\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6867\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6864\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6861\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6867\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__6864\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6861\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\
        );

    \I__1279\ : IoInMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6848\,
            I => \N__6844\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__6847\,
            I => \N__6838\
        );

    \I__1276\ : Span4Mux_s1_v
    port map (
            O => \N__6844\,
            I => \N__6832\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6825\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6825\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6825\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6820\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6820\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6815\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6815\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__6832\,
            I => \N__6812\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6807\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6807\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6815\,
            I => \N__6804\
        );

    \I__1264\ : Sp12to4
    port map (
            O => \N__6812\,
            I => \N__6801\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__6807\,
            I => \N__6798\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6804\,
            I => \N__6795\
        );

    \I__1261\ : Span12Mux_h
    port map (
            O => \N__6801\,
            I => \N__6792\
        );

    \I__1260\ : Sp12to4
    port map (
            O => \N__6798\,
            I => \N__6789\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__6795\,
            I => \N__6786\
        );

    \I__1258\ : Span12Mux_v
    port map (
            O => \N__6792\,
            I => \N__6779\
        );

    \I__1257\ : Span12Mux_h
    port map (
            O => \N__6789\,
            I => \N__6779\
        );

    \I__1256\ : Sp12to4
    port map (
            O => \N__6786\,
            I => \N__6779\
        );

    \I__1255\ : Span12Mux_v
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1254\ : Odrv12
    port map (
            O => \N__6776\,
            I => \TEAn_c\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6764\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6764\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6761\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6756\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6756\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6764\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6761\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6737\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6737\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6730\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6730\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6730\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6725\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6725\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6722\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6737\,
            I => \N__6719\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6730\,
            I => \N__6716\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6713\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6722\,
            I => \N__6710\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__6719\,
            I => \N__6704\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__6716\,
            I => \N__6704\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__6713\,
            I => \N__6701\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__6710\,
            I => \N__6698\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6695\
        );

    \I__1228\ : Sp12to4
    port map (
            O => \N__6704\,
            I => \N__6688\
        );

    \I__1227\ : Sp12to4
    port map (
            O => \N__6701\,
            I => \N__6688\
        );

    \I__1226\ : Sp12to4
    port map (
            O => \N__6698\,
            I => \N__6688\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6695\,
            I => \N__6685\
        );

    \I__1224\ : Span12Mux_h
    port map (
            O => \N__6688\,
            I => \N__6680\
        );

    \I__1223\ : Span12Mux_s7_h
    port map (
            O => \N__6685\,
            I => \N__6680\
        );

    \I__1222\ : Span12Mux_v
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1221\ : Odrv12
    port map (
            O => \N__6677\,
            I => \RESETn_c\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6668\,
            I => \READ_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__1217\ : IoInMux
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1215\ : Span12Mux_s8_v
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1214\ : Span12Mux_h
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__6653\,
            I => \N_207_i\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1209\ : Sp12to4
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1208\ : Span12Mux_h
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1207\ : Odrv12
    port map (
            O => \N__6635\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__1206\ : IoInMux
    port map (
            O => \N__6632\,
            I => \N__6629\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1204\ : Span4Mux_s2_h
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1203\ : Span4Mux_v
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__1202\ : Sp12to4
    port map (
            O => \N__6620\,
            I => \N__6617\
        );

    \I__1201\ : Span12Mux_h
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__1200\ : Odrv12
    port map (
            O => \N__6614\,
            I => \un2_D_LL_AMIGA_0\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1196\ : Sp12to4
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1195\ : Span12Mux_h
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1194\ : Odrv12
    port map (
            O => \N__6596\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__1193\ : IoInMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1191\ : IoSpan4Mux
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1190\ : IoSpan4Mux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1189\ : Span4Mux_s2_h
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1188\ : Sp12to4
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1187\ : Span12Mux_h
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__1186\ : Odrv12
    port map (
            O => \N__6572\,
            I => \un2_D_LL_AMIGA_2\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6560\,
            I => \READ_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__1181\ : IoInMux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1179\ : Span12Mux_s4_h
    port map (
            O => \N__6551\,
            I => \N__6548\
        );

    \I__1178\ : Span12Mux_h
    port map (
            O => \N__6548\,
            I => \N__6545\
        );

    \I__1177\ : Odrv12
    port map (
            O => \N__6545\,
            I => \N_231_i\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6536\
        );

    \I__1174\ : Span12Mux_v
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1173\ : Span12Mux_h
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__1172\ : Odrv12
    port map (
            O => \N__6530\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1169\ : IoSpan4Mux
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1168\ : Sp12to4
    port map (
            O => \N__6518\,
            I => \N__6515\
        );

    \I__1167\ : Span12Mux_s7_h
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1166\ : Span12Mux_v
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__6509\,
            I => \un2_D_LL_AMIGA_7\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6506\,
            I => \N__6503\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6495\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6492\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6489\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__6495\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6492\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6489\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6482\,
            I => \N__6478\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6475\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6469\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__6469\,
            I => \N__6462\
        );

    \I__1150\ : Span4Mux_v
    port map (
            O => \N__6466\,
            I => \N__6459\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6456\
        );

    \I__1148\ : Sp12to4
    port map (
            O => \N__6462\,
            I => \N__6449\
        );

    \I__1147\ : Sp12to4
    port map (
            O => \N__6459\,
            I => \N__6449\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6449\
        );

    \I__1145\ : Span12Mux_h
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1144\ : Span12Mux_v
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1143\ : Odrv12
    port map (
            O => \N__6443\,
            I => \PORTSIZE_c\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6437\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6437\,
            I => \N__6429\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6424\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6424\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6419\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6419\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6416\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__6429\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6424\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6419\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6416\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__6407\,
            I => \U111_CYCLE_SM.N_60_cascade_\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__6395\,
            I => \READ_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__1126\ : IoInMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1124\ : Span4Mux_s1_v
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__1123\ : Span4Mux_v
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1122\ : Sp12to4
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1121\ : Span12Mux_h
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1120\ : Odrv12
    port map (
            O => \N__6374\,
            I => \N_211_i\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__6371\,
            I => \U111_CYCLE_SM.N_75_cascade_\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6365\,
            I => \U111_CYCLE_SM.LATCH_EN_5\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__6362\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6352\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6349\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6342\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6356\,
            I => \N__6342\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6342\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6352\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6349\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6329\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6329\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1104\ : Span4Mux_h
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1102\ : Span12Mux_v
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1101\ : Span12Mux_h
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__6314\,
            I => \SIZ_c_1\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__6311\,
            I => \N__6307\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \N__6304\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6301\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6298\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6293\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6298\,
            I => \N__6293\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1090\ : Span12Mux_h
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__6281\,
            I => \SIZ_c_0\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__6272\,
            I => \WRITE_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__6263\,
            I => \WRITE_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__6251\,
            I => \WRITE_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__1078\ : IoInMux
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1076\ : Span4Mux_s3_v
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__6239\,
            I => \LBENn_c_i_0\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6233\,
            I => \U111_CYCLE_SM.N_33\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U111_CYCLE_SM.N_49\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6221\,
            I => \U111_CYCLE_SM.N_75\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1066\ : Span12Mux_h
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1065\ : Span12Mux_v
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__6206\,
            I => \TS_CPUn_c\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__1061\ : Span4Mux_h
    port map (
            O => \N__6197\,
            I => \N__6194\
        );

    \I__1060\ : Sp12to4
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1059\ : Span12Mux_h
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__6188\,
            I => \BGn_c\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6181\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6178\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6181\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6178\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1050\ : Span4Mux_h
    port map (
            O => \N__6164\,
            I => \N__6161\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6161\,
            I => \WRITE_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__1045\ : Span4Mux_h
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__6146\,
            I => \WRITE_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1041\ : Odrv12
    port map (
            O => \N__6137\,
            I => \WRITE_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__1040\ : IoInMux
    port map (
            O => \N__6134\,
            I => \N__6130\
        );

    \I__1039\ : IoInMux
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6127\,
            I => \N__6119\
        );

    \I__1036\ : Span4Mux_s2_v
    port map (
            O => \N__6124\,
            I => \N__6116\
        );

    \I__1035\ : IoInMux
    port map (
            O => \N__6123\,
            I => \N__6113\
        );

    \I__1034\ : IoInMux
    port map (
            O => \N__6122\,
            I => \N__6110\
        );

    \I__1033\ : IoSpan4Mux
    port map (
            O => \N__6119\,
            I => \N__6107\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__6116\,
            I => \N__6104\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6113\,
            I => \N__6101\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6098\
        );

    \I__1029\ : Span4Mux_s3_h
    port map (
            O => \N__6107\,
            I => \N__6095\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6104\,
            I => \N__6090\
        );

    \I__1027\ : Span4Mux_s2_v
    port map (
            O => \N__6101\,
            I => \N__6090\
        );

    \I__1026\ : IoSpan4Mux
    port map (
            O => \N__6098\,
            I => \N__6087\
        );

    \I__1025\ : Span4Mux_h
    port map (
            O => \N__6095\,
            I => \N__6084\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__6090\,
            I => \N__6081\
        );

    \I__1023\ : Span4Mux_s3_h
    port map (
            O => \N__6087\,
            I => \N__6078\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__6084\,
            I => \N__6075\
        );

    \I__1021\ : Span4Mux_v
    port map (
            O => \N__6081\,
            I => \N__6072\
        );

    \I__1020\ : Span4Mux_h
    port map (
            O => \N__6078\,
            I => \N__6069\
        );

    \I__1019\ : Span4Mux_h
    port map (
            O => \N__6075\,
            I => \N__6066\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__6072\,
            I => \N__6061\
        );

    \I__1017\ : Span4Mux_h
    port map (
            O => \N__6069\,
            I => \N__6061\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__6066\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__6061\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__6050\,
            I => \N__6047\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__6047\,
            I => \WRITE_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6038\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6038\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1007\ : Span12Mux_h
    port map (
            O => \N__6035\,
            I => \N__6031\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__1005\ : Odrv12
    port map (
            O => \N__6031\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6028\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1000\ : Span4Mux_h
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6011\,
            I => \U111_CYCLE_SM.N_67\
        );

    \I__998\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6004\
        );

    \I__997\ : InMux
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6004\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6001\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__994\ : IoInMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__992\ : IoSpan4Mux
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__991\ : Span4Mux_s2_h
    port map (
            O => \N__5987\,
            I => \N__5983\
        );

    \I__990\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__989\ : Span4Mux_v
    port map (
            O => \N__5983\,
            I => \N__5977\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5974\
        );

    \I__987\ : Sp12to4
    port map (
            O => \N__5977\,
            I => \N__5971\
        );

    \I__986\ : Sp12to4
    port map (
            O => \N__5974\,
            I => \N__5968\
        );

    \I__985\ : Span12Mux_s9_h
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__984\ : Span12Mux_v
    port map (
            O => \N__5968\,
            I => \N__5962\
        );

    \I__983\ : Span12Mux_h
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__982\ : Span12Mux_h
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__981\ : Odrv12
    port map (
            O => \N__5959\,
            I => \D_LM_040_in_5\
        );

    \I__980\ : Odrv12
    port map (
            O => \N__5956\,
            I => \D_LM_040_in_5\
        );

    \I__979\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5948\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5948\,
            I => \N__5945\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__976\ : Span4Mux_h
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__975\ : Sp12to4
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__974\ : Span12Mux_h
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__973\ : Odrv12
    port map (
            O => \N__5933\,
            I => \D_UU_040_in_5\
        );

    \I__972\ : IoInMux
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__970\ : Span4Mux_s3_h
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__5912\,
            I => \un1_D_UU_040_5\
        );

    \I__965\ : IoInMux
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__963\ : IoSpan4Mux
    port map (
            O => \N__5903\,
            I => \N__5899\
        );

    \I__962\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5896\
        );

    \I__961\ : IoSpan4Mux
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5896\,
            I => \N__5890\
        );

    \I__959\ : Span4Mux_s2_h
    port map (
            O => \N__5893\,
            I => \N__5887\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__5890\,
            I => \N__5884\
        );

    \I__957\ : Sp12to4
    port map (
            O => \N__5887\,
            I => \N__5881\
        );

    \I__956\ : Sp12to4
    port map (
            O => \N__5884\,
            I => \N__5878\
        );

    \I__955\ : Span12Mux_h
    port map (
            O => \N__5881\,
            I => \N__5873\
        );

    \I__954\ : Span12Mux_v
    port map (
            O => \N__5878\,
            I => \N__5873\
        );

    \I__953\ : Span12Mux_h
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__952\ : Odrv12
    port map (
            O => \N__5870\,
            I => \D_LM_040_in_3\
        );

    \I__951\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__948\ : Span4Mux_h
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__947\ : Sp12to4
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__946\ : Span12Mux_h
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__945\ : Odrv12
    port map (
            O => \N__5849\,
            I => \D_UU_040_in_3\
        );

    \I__944\ : IoInMux
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5840\
        );

    \I__942\ : IoSpan4Mux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__941\ : Sp12to4
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__940\ : Span12Mux_s6_v
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__939\ : Odrv12
    port map (
            O => \N__5831\,
            I => \un1_D_UU_040_3\
        );

    \I__938\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__936\ : Span4Mux_v
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__934\ : Span12Mux_h
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__933\ : Odrv12
    port map (
            O => \N__5813\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__932\ : IoInMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__930\ : IoSpan4Mux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__929\ : Span4Mux_s1_h
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__928\ : Span4Mux_v
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__927\ : Sp12to4
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__926\ : Span12Mux_s10_h
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__5789\,
            I => \un2_D_LL_AMIGA_3\
        );

    \I__924\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__921\ : Sp12to4
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5774\,
            I => \WRITE_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__919\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__916\ : Span4Mux_h
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__5759\,
            I => \WRITE_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__914\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5750\,
            I => \N__5747\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__5747\,
            I => \WRITE_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__910\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5735\,
            I => \WRITE_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__906\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__904\ : Span4Mux_h
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__902\ : Span4Mux_h
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__5717\,
            I => \WRITE_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__900\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__898\ : Span4Mux_v
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__5705\,
            I => \WRITE_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__896\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__5693\,
            I => \WRITE_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__892\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__890\ : Odrv12
    port map (
            O => \N__5684\,
            I => \WRITE_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__889\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5678\,
            I => \WRITE_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__887\ : IoInMux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__885\ : IoSpan4Mux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__884\ : Span4Mux_s1_v
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__882\ : Span12Mux_s9_v
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__881\ : Odrv12
    port map (
            O => \N__5657\,
            I => \N_244_i\
        );

    \I__880\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__5642\,
            I => \WRITE_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__875\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__5633\,
            I => \WRITE_CYCLE_ACTIVE_i_ess\
        );

    \I__872\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5624\,
            I => \WRITE_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__869\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__867\ : Span12Mux_s6_h
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__5612\,
            I => \WRITE_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__865\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__863\ : Span4Mux_h
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5597\,
            I => \WRITE_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__860\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__5585\,
            I => \WRITE_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__856\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__854\ : Sp12to4
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__853\ : Span12Mux_v
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__852\ : Odrv12
    port map (
            O => \N__5570\,
            I => \WRITE_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__851\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__848\ : Span4Mux_h
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__5555\,
            I => \WRITE_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__846\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__844\ : Span4Mux_h
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__5540\,
            I => \WRITE_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__841\ : IoInMux
    port map (
            O => \N__5537\,
            I => \N__5534\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__839\ : IoSpan4Mux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__5528\,
            I => \N__5525\
        );

    \I__837\ : Span12Mux_s7_h
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__836\ : Span12Mux_h
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__835\ : Odrv12
    port map (
            O => \N__5519\,
            I => \un2_D_LM_AMIGA_0\
        );

    \I__834\ : IoInMux
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__832\ : Span4Mux_s3_h
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__5504\,
            I => \N__5501\
        );

    \I__829\ : Span4Mux_h
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__5498\,
            I => \N_268_i\
        );

    \I__827\ : IoInMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__825\ : Span12Mux_s11_h
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__5486\,
            I => \N_255_i\
        );

    \I__823\ : IoInMux
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__821\ : IoSpan4Mux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__820\ : Span4Mux_s1_v
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__819\ : Sp12to4
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__818\ : Span12Mux_v
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__5465\,
            I => \TSn_c\
        );

    \I__816\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__814\ : Span12Mux_s8_h
    port map (
            O => \N__5456\,
            I => \N__5453\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__5453\,
            I => \WRITE_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__812\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__5441\,
            I => \WRITE_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__808\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__5429\,
            I => \WRITE_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__804\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__5414\,
            I => \WRITE_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__799\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__797\ : Span12Mux_h
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__5402\,
            I => \WRITE_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__795\ : IoInMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__793\ : Span4Mux_s2_v
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__5384\,
            I => \N_237_i\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__5381\,
            I => \N__5377\
        );

    \I__788\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5374\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5371\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5374\,
            I => \N__5368\
        );

    \I__785\ : IoSpan4Mux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__784\ : Span4Mux_v
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__783\ : IoSpan4Mux
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__782\ : Sp12to4
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__781\ : Span4Mux_s2_h
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__778\ : Span12Mux_v
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__777\ : Span12Mux_h
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__776\ : Span12Mux_v
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__775\ : Span12Mux_h
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__774\ : Odrv12
    port map (
            O => \N__5338\,
            I => \D_LM_040_in_0\
        );

    \I__773\ : Odrv12
    port map (
            O => \N__5335\,
            I => \D_LM_040_in_0\
        );

    \I__772\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__768\ : Sp12to4
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__767\ : Span12Mux_h
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__5312\,
            I => \D_UU_040_in_0\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__763\ : Span4Mux_s2_v
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__5294\,
            I => \un1_D_UU_040_0\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__757\ : IoSpan4Mux
    port map (
            O => \N__5285\,
            I => \N__5281\
        );

    \I__756\ : IoInMux
    port map (
            O => \N__5284\,
            I => \N__5278\
        );

    \I__755\ : IoSpan4Mux
    port map (
            O => \N__5281\,
            I => \N__5275\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5278\,
            I => \N__5272\
        );

    \I__753\ : IoSpan4Mux
    port map (
            O => \N__5275\,
            I => \N__5267\
        );

    \I__752\ : IoSpan4Mux
    port map (
            O => \N__5272\,
            I => \N__5267\
        );

    \I__751\ : Span4Mux_s3_v
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__5264\,
            I => \CONSTANT_ONE_NET\
        );

    \I__749\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__747\ : Span12Mux_v
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__5252\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__745\ : IoInMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__743\ : Span4Mux_s0_h
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__742\ : Sp12to4
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__741\ : Span12Mux_s11_v
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__740\ : Span12Mux_h
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__739\ : Odrv12
    port map (
            O => \N__5231\,
            I => \un2_D_LL_AMIGA_6\
        );

    \I__738\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__736\ : Span12Mux_h
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__5219\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__732\ : Span12Mux_s8_h
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__731\ : Span12Mux_h
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__5204\,
            I => \un2_D_LM_AMIGA_1\
        );

    \I__729\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5198\,
            I => \N__5195\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__726\ : Sp12to4
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__724\ : Odrv12
    port map (
            O => \N__5186\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__723\ : IoInMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5180\,
            I => \N__5177\
        );

    \I__721\ : IoSpan4Mux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__720\ : Span4Mux_s3_h
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__717\ : Sp12to4
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__716\ : Odrv12
    port map (
            O => \N__5162\,
            I => \un2_D_LM_AMIGA_3\
        );

    \I__715\ : IoInMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__713\ : IoSpan4Mux
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__712\ : Span4Mux_s3_v
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__711\ : Span4Mux_v
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__5144\,
            I => \LBENn_c_i\
        );

    \I__709\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__707\ : IoInMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5131\,
            I => \N__5125\
        );

    \I__704\ : Span4Mux_h
    port map (
            O => \N__5128\,
            I => \N__5122\
        );

    \I__703\ : Span12Mux_s5_h
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__5119\,
            I => \N__5113\
        );

    \I__700\ : Sp12to4
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__699\ : Span12Mux_v
    port map (
            O => \N__5113\,
            I => \N__5107\
        );

    \I__698\ : Span12Mux_h
    port map (
            O => \N__5110\,
            I => \N__5104\
        );

    \I__697\ : Span12Mux_h
    port map (
            O => \N__5107\,
            I => \N__5099\
        );

    \I__696\ : Span12Mux_v
    port map (
            O => \N__5104\,
            I => \N__5099\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__5099\,
            I => \D_LM_040_in_2\
        );

    \I__694\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__691\ : Span4Mux_h
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__689\ : Span12Mux_h
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__5078\,
            I => \D_UU_040_in_2\
        );

    \I__687\ : IoInMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__685\ : IoSpan4Mux
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__684\ : Span4Mux_s2_v
    port map (
            O => \N__5066\,
            I => \N__5063\
        );

    \I__683\ : Span4Mux_v
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__5060\,
            I => \un1_D_UU_040_2\
        );

    \I__681\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__679\ : Span4Mux_v
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__678\ : Sp12to4
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__677\ : Span12Mux_h
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__676\ : Odrv12
    port map (
            O => \N__5042\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__675\ : IoInMux
    port map (
            O => \N__5039\,
            I => \N__5036\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__673\ : Span12Mux_s5_h
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__5030\,
            I => \N_256_i\
        );

    \I__671\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5024\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__5021\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__668\ : IoInMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__666\ : Sp12to4
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__665\ : Span12Mux_s5_h
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__664\ : Span12Mux_h
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__663\ : Span12Mux_v
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__5000\,
            I => \un2_D_LM_AMIGA_2\
        );

    \I__661\ : IoInMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__659\ : Span12Mux_s8_h
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__4988\,
            I => \N_245_i\
        );

    \I__657\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__654\ : Sp12to4
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__653\ : Odrv12
    port map (
            O => \N__4973\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__652\ : IoInMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__650\ : IoSpan4Mux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__648\ : Span12Mux_s9_h
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__647\ : Span12Mux_h
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__4952\,
            I => \un2_D_LM_AMIGA_4\
        );

    \I__645\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__4937\,
            I => \WRITE_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__640\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4931\,
            I => \WRITE_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__638\ : IoInMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__636\ : IoSpan4Mux
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__635\ : Span4Mux_s2_h
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__634\ : Span4Mux_h
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__633\ : Span4Mux_h
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__4910\,
            I => \N_259_i\
        );

    \I__631\ : IoInMux
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__629\ : IoSpan4Mux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__628\ : IoSpan4Mux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__627\ : Span4Mux_s2_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__4889\,
            I => \N_240_i\
        );

    \I__624\ : IoInMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__622\ : Span12Mux_s7_v
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4877\,
            I => \N_243_i\
        );

    \I__620\ : IoInMux
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__618\ : Span4Mux_s2_h
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__617\ : Sp12to4
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__616\ : Span12Mux_s9_v
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__615\ : Odrv12
    port map (
            O => \N__4859\,
            I => \N_263_i\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__612\ : Span4Mux_s2_h
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__609\ : Span4Mux_h
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__4838\,
            I => \N_265_i\
        );

    \I__607\ : IoInMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__605\ : Span12Mux_s9_h
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__4826\,
            I => \N_257_i\
        );

    \I__603\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__599\ : Odrv12
    port map (
            O => \N__4811\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__598\ : IoInMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__596\ : Span12Mux_s10_h
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__595\ : Span12Mux_h
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__4796\,
            I => \un2_D_LM_AMIGA_5\
        );

    \I__593\ : IoInMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__591\ : Span12Mux_s10_v
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__590\ : Odrv12
    port map (
            O => \N__4784\,
            I => \N_250_i\
        );

    \I__589\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__585\ : Span4Mux_h
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__4766\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__583\ : IoInMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__581\ : IoSpan4Mux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__580\ : Span4Mux_s3_h
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__578\ : Span12Mux_s11_h
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__4745\,
            I => \un2_D_LM_AMIGA_7\
        );

    \I__576\ : IoInMux
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__574\ : IoSpan4Mux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__573\ : Span4Mux_s3_h
    port map (
            O => \N__4733\,
            I => \N__4730\
        );

    \I__572\ : Span4Mux_h
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__4727\,
            I => \N_238_i\
        );

    \I__570\ : IoInMux
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__568\ : Span4Mux_s3_v
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__4712\,
            I => \N_241_i\
        );

    \I__565\ : IoInMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__563\ : Span12Mux_s10_h
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__562\ : Odrv12
    port map (
            O => \N__4700\,
            I => \N_261_i\
        );

    \I__561\ : IoInMux
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__559\ : IoSpan4Mux
    port map (
            O => \N__4691\,
            I => \N__4688\
        );

    \I__558\ : Span4Mux_s1_h
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__557\ : Span4Mux_h
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__4682\,
            I => \N_248_i\
        );

    \I__555\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__552\ : Sp12to4
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__4667\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__550\ : IoInMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__548\ : Span4Mux_s2_h
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__546\ : Sp12to4
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__545\ : Span12Mux_s11_h
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__544\ : Span12Mux_h
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__4643\,
            I => \un2_D_LL_AMIGA_5\
        );

    \I__542\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__540\ : Span4Mux_h
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__539\ : Span4Mux_h
    port map (
            O => \N__4631\,
            I => \N__4627\
        );

    \I__538\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4624\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__4627\,
            I => \N__4621\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4618\
        );

    \I__535\ : Span12Mux_v
    port map (
            O => \N__4621\,
            I => \N__4613\
        );

    \I__534\ : Span12Mux_h
    port map (
            O => \N__4618\,
            I => \N__4613\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__4613\,
            I => \A_040_c_1\
        );

    \I__532\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__528\ : Odrv12
    port map (
            O => \N__4598\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__527\ : IoInMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__525\ : IoSpan4Mux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__524\ : Span4Mux_s0_h
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__523\ : Sp12to4
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__522\ : Span12Mux_h
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__4577\,
            I => \un2_D_LM_AMIGA_6\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__518\ : IoSpan4Mux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__517\ : IoSpan4Mux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__516\ : Span4Mux_s3_h
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__515\ : Span4Mux_h
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__4556\,
            I => \N_242_i\
        );

    \I__513\ : IoInMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__511\ : IoSpan4Mux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__510\ : Span4Mux_s3_h
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__509\ : Span4Mux_h
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__4538\,
            I => \N_260_i\
        );

    \I__507\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4528\
        );

    \I__505\ : IoInMux
    port map (
            O => \N__4531\,
            I => \N__4525\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4519\
        );

    \I__502\ : Sp12to4
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__501\ : Span4Mux_s2_h
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__500\ : Span12Mux_h
    port map (
            O => \N__4516\,
            I => \N__4510\
        );

    \I__499\ : Span4Mux_v
    port map (
            O => \N__4513\,
            I => \N__4507\
        );

    \I__498\ : Span12Mux_h
    port map (
            O => \N__4510\,
            I => \N__4504\
        );

    \I__497\ : Sp12to4
    port map (
            O => \N__4507\,
            I => \N__4501\
        );

    \I__496\ : Span12Mux_v
    port map (
            O => \N__4504\,
            I => \N__4498\
        );

    \I__495\ : Span12Mux_s11_h
    port map (
            O => \N__4501\,
            I => \N__4495\
        );

    \I__494\ : Span12Mux_v
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__493\ : Span12Mux_h
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__492\ : Odrv12
    port map (
            O => \N__4492\,
            I => \D_LL_040_in_3\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__4489\,
            I => \D_LL_040_in_3\
        );

    \I__490\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__486\ : Sp12to4
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__485\ : Span12Mux_h
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__484\ : Odrv12
    port map (
            O => \N__4466\,
            I => \D_UM_040_in_3\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__481\ : IoSpan4Mux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__480\ : Span4Mux_s2_h
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__479\ : Span4Mux_h
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__4448\,
            I => \un1_D_UM_040_3\
        );

    \I__477\ : IoInMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__475\ : Span4Mux_s3_v
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__474\ : Span4Mux_v
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__4433\,
            I => \N_239_i\
        );

    \I__472\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__470\ : Span4Mux_v
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__468\ : Span12Mux_h
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__4412\,
            I => \D_UU_040_in_6\
        );

    \I__465\ : IoInMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__463\ : Span4Mux_s2_h
    port map (
            O => \N__4403\,
            I => \N__4399\
        );

    \I__462\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4396\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__4399\,
            I => \N__4393\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__458\ : Sp12to4
    port map (
            O => \N__4390\,
            I => \N__4384\
        );

    \I__457\ : Span12Mux_h
    port map (
            O => \N__4387\,
            I => \N__4381\
        );

    \I__456\ : Span12Mux_s11_v
    port map (
            O => \N__4384\,
            I => \N__4378\
        );

    \I__455\ : Span12Mux_h
    port map (
            O => \N__4381\,
            I => \N__4375\
        );

    \I__454\ : Span12Mux_h
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__4375\,
            I => \D_LM_040_in_6\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__4372\,
            I => \D_LM_040_in_6\
        );

    \I__451\ : IoInMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__449\ : Span4Mux_s2_v
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__448\ : Span4Mux_h
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__4352\,
            I => \un1_D_UU_040_6\
        );

    \I__445\ : IoInMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__443\ : IoSpan4Mux
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__442\ : IoSpan4Mux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__441\ : Span4Mux_s3_h
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__4334\,
            I => \N_253_i\
        );

    \I__439\ : IoInMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__437\ : IoSpan4Mux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__436\ : Span4Mux_s3_h
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__4316\,
            I => \N_254_i\
        );

    \I__433\ : IoInMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__431\ : IoSpan4Mux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__430\ : Span4Mux_s3_h
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__4298\,
            I => \N_252_i\
        );

    \I__427\ : IoInMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4289\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__424\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__422\ : Span4Mux_h
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__4274\,
            I => \A_040_c_0\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__417\ : Span4Mux_s2_v
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__416\ : Span4Mux_v
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__4259\,
            I => \A_AMIGA_c_0\
        );

    \I__414\ : IoInMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__412\ : Span4Mux_s2_h
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__411\ : Span4Mux_v
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__410\ : Span4Mux_h
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__409\ : Odrv4
    port map (
            O => \N__4241\,
            I => \N_264_i\
        );

    \I__408\ : IoInMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__406\ : IoSpan4Mux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__405\ : IoSpan4Mux
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__404\ : Span4Mux_s2_h
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__403\ : Span4Mux_h
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__4220\,
            I => \N_262_i\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__399\ : Span4Mux_s2_h
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__4205\,
            I => \N_258_i\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__393\ : Span4Mux_s3_h
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__4190\,
            I => \N_246_i\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__389\ : Span4Mux_s0_v
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__388\ : Sp12to4
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__387\ : Span12Mux_h
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__386\ : Span12Mux_v
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__385\ : Span12Mux_v
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__4166\,
            I => \TAn_in\
        );

    \I__383\ : IoInMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__381\ : Span4Mux_s0_h
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__380\ : Span4Mux_h
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__379\ : Odrv4
    port map (
            O => \N__4151\,
            I => \N_267_i\
        );

    \I__378\ : IoInMux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__376\ : Odrv12
    port map (
            O => \N__4142\,
            I => \RESETn_c_i\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__373\ : Span4Mux_s1_h
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__371\ : Span4Mux_h
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__370\ : Odrv4
    port map (
            O => \N__4124\,
            I => \N_266_i\
        );

    \I__369\ : IoInMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__4115\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_0\
        );

    \I__366\ : IoInMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__364\ : Span4Mux_s3_h
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__363\ : Odrv4
    port map (
            O => \N__4103\,
            I => \N_247_i\
        );

    \I__362\ : IoInMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__360\ : IoSpan4Mux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__359\ : Span4Mux_s0_h
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__358\ : Span4Mux_h
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__4085\,
            I => \N_249_i\
        );

    \I__356\ : IoInMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__354\ : IoSpan4Mux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__353\ : Span4Mux_s3_v
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__352\ : Span4Mux_v
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__4067\,
            I => \N_251_i\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__348\ : Span4Mux_s0_h
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__347\ : Span4Mux_h
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__346\ : Span4Mux_h
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__345\ : Sp12to4
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__344\ : Span12Mux_v
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__343\ : Span12Mux_v
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__342\ : Span12Mux_h
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__4037\,
            I => \TCIn_c\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__9410\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4148\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4121\,
            GLOBALBUFFEROUTPUT => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5786\,
            lcout => \N_267_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6709\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_5_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5732\,
            lcout => \N_266_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9251\,
            in2 => \_gnd_net_\,
            in3 => \N__7094\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_2_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5621\,
            lcout => \N_247_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_4_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5690\,
            lcout => \N_249_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_6_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5771\,
            lcout => \N_251_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_0_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4949\,
            lcout => \N_253_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_1_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5462\,
            lcout => \N_254_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_7_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6143\,
            lcout => \N_252_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4630\,
            in2 => \_gnd_net_\,
            in3 => \N__6044\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6043\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4286\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_3_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_264_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_1_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5426\,
            lcout => \N_262_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_5_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5567\,
            lcout => \N_258_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_1_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6278\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_246_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_3_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_248_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11163\,
            in1 => \N__7409\,
            in2 => \_gnd_net_\,
            in3 => \N__4679\,
            lcout => \un2_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6465\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4640\,
            lcout => \U111_CYCLE_SM.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11118\,
            in1 => \N__8823\,
            in2 => \_gnd_net_\,
            in3 => \N__4610\,
            lcout => \un2_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_5_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6158\,
            lcout => \N_242_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_7_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_260_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11139\,
            in1 => \N__4535\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_2_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5552\,
            lcout => \N_239_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4430\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__11166\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_2_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_263_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_4_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5654\,
            lcout => \N_265_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_4_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4934\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_257_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8352\,
            in1 => \N__4823\,
            in2 => \_gnd_net_\,
            in3 => \N__11086\,
            lcout => \un2_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_5_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_250_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4781\,
            in1 => \N__10471\,
            in2 => \_gnd_net_\,
            in3 => \N__11117\,
            lcout => \un2_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_1_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_238_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_4_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_241_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_261_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5450\,
            lcout => \N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10971\,
            in1 => \N__7319\,
            in2 => \_gnd_net_\,
            in3 => \N__5027\,
            lcout => \un2_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5438\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_245_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11048\,
            in1 => \N__8452\,
            in2 => \_gnd_net_\,
            in3 => \N__4985\,
            lcout => \un2_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10077\,
            in2 => \_gnd_net_\,
            in3 => \N__9690\,
            lcout => \WRITE_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9409\,
            ce => \N__9297\,
            sr => \N__9225\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9691\,
            in1 => \_gnd_net_\,
            in2 => \N__10090\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9409\,
            ce => \N__9297\,
            sr => \N__9225\
        );

    \D_LM_AMIGA_iobuf_RNO_6_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5594\,
            lcout => \N_259_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_3_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_240_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_6_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6260\,
            lcout => \N_243_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_0_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5582\,
            lcout => \N_237_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5380\,
            in1 => \N__5330\,
            in2 => \_gnd_net_\,
            in3 => \N__11120\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5261\,
            in1 => \N__9095\,
            in2 => \_gnd_net_\,
            in3 => \N__11130\,
            lcout => \un2_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7545\,
            in1 => \N__5228\,
            in2 => \_gnd_net_\,
            in3 => \N__11046\,
            lcout => \un2_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8761\,
            in1 => \N__5201\,
            in2 => \_gnd_net_\,
            in3 => \N__11047\,
            lcout => \un2_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BUFENn_obuf_RNO_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8051\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__5096\,
            in2 => \_gnd_net_\,
            in3 => \N__11119\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5057\,
            in1 => \N__8168\,
            in2 => \_gnd_net_\,
            in3 => \N__11076\,
            lcout => \un2_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_7_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5639\,
            lcout => \N_268_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5630\,
            lcout => \N_255_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__6742\,
            in1 => \N__6007\,
            in2 => \N__8050\,
            in3 => \N__6185\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10002\,
            lcout => \WRITE_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9610\,
            lcout => \WRITE_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9615\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10000\,
            lcout => \READ_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9614\,
            lcout => \WRITE_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9611\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10004\,
            lcout => \WRITE_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9612\,
            lcout => \WRITE_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10006\,
            lcout => \WRITE_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10001\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9608\,
            lcout => \WRITE_CYCLE_ACTIVE_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => \N__9299\,
            sr => \N__9227\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9992\,
            in2 => \_gnd_net_\,
            in3 => \N__9571\,
            lcout => \WRITE_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9570\,
            in1 => \_gnd_net_\,
            in2 => \N__10047\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9999\,
            in2 => \_gnd_net_\,
            in3 => \N__9574\,
            lcout => \WRITE_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9573\,
            in1 => \_gnd_net_\,
            in2 => \N__10049\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9988\,
            in2 => \_gnd_net_\,
            in3 => \N__9569\,
            lcout => \WRITE_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9572\,
            in1 => \_gnd_net_\,
            in2 => \N__10048\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => \N__9301\,
            sr => \N__9231\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9850\,
            in2 => \_gnd_net_\,
            in3 => \N__9620\,
            lcout => \WRITE_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9842\,
            in2 => \_gnd_net_\,
            in3 => \N__9616\,
            lcout => \WRITE_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9617\,
            in1 => \_gnd_net_\,
            in2 => \N__9899\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9846\,
            in2 => \_gnd_net_\,
            in3 => \N__9618\,
            lcout => \WRITE_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9619\,
            in1 => \_gnd_net_\,
            in2 => \N__9900\,
            in3 => \_gnd_net_\,
            lcout => \WRITE_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9851\,
            in2 => \_gnd_net_\,
            in3 => \N__9621\,
            lcout => \WRITE_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => \N__9302\,
            sr => \N__9235\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10009\,
            lcout => \WRITE_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => \N__9304\,
            sr => \N__9238\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9681\,
            lcout => \WRITE_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => \N__9304\,
            sr => \N__9238\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10008\,
            lcout => \WRITE_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => \N__9304\,
            sr => \N__9238\
        );

    \D_UU_AMIGA_iobuf_RNO_7_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5681\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_244_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5986\,
            in1 => \N__5951\,
            in2 => \_gnd_net_\,
            in3 => \N__11144\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5902\,
            in1 => \N__5867\,
            in2 => \_gnd_net_\,
            in3 => \N__11143\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5828\,
            in1 => \N__7485\,
            in2 => \_gnd_net_\,
            in3 => \N__11111\,
            lcout => \un2_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \READ_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9418\,
            ce => \N__9307\,
            sr => \N__9236\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9719\,
            lcout => \READ_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9418\,
            ce => \N__9307\,
            sr => \N__9236\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10085\,
            lcout => \READ_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9418\,
            ce => \N__9307\,
            sr => \N__9236\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9696\,
            lcout => \READ_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9417\,
            ce => \N__9305\,
            sr => \N__9232\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9695\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10081\,
            lcout => \READ_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9417\,
            ce => \N__9305\,
            sr => \N__9232\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10083\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9694\,
            lcout => \WRITE_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9417\,
            ce => \N__9305\,
            sr => \N__9232\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10058\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \READ_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9416\,
            ce => \N__9303\,
            sr => \N__9228\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9422\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10057\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => \READ_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9412\,
            ce => \N__9300\,
            sr => \N__9224\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10050\,
            lcout => \READ_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9411\,
            ce => \N__9296\,
            sr => \N__9226\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9692\,
            lcout => \WRITE_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9411\,
            ce => \N__9296\,
            sr => \N__9226\
        );

    \U111_CYCLE_SM.A2_EN_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__6034\,
            in1 => \N__6224\,
            in2 => \_gnd_net_\,
            in3 => \N__6941\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__9229\
        );

    \U111_CYCLE_SM.TA_DIS_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101110010"
        )
    port map (
            in0 => \N__6436\,
            in1 => \N__6236\,
            in2 => \N__8068\,
            in3 => \N__6943\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__9229\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__6942\,
            in1 => \N__6023\,
            in2 => \N__10970\,
            in3 => \N__6435\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__9229\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__6368\,
            in1 => \N__6940\,
            in2 => \N__10326\,
            in3 => \N__6359\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__9229\
        );

    \U111_CYCLE_SM.TS_EN_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__6230\,
            in1 => \N__6008\,
            in2 => \N__6917\,
            in3 => \N__7250\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__9229\
        );

    \U111_CYCLE_SM.TS_DELAY_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6218\,
            lcout => \U111_CYCLE_SM.TS_DELAYZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9401\,
            ce => 'H',
            sr => \N__9233\
        );

    \U111_CYCLE_SM.TS_DELAY_RNI91BJ_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__6203\,
            in1 => \N__8049\,
            in2 => \_gnd_net_\,
            in3 => \N__6184\,
            lcout => \U111_CYCLE_SM.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9837\,
            lcout => \READ_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9575\,
            lcout => \WRITE_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9835\,
            lcout => \READ_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9579\,
            lcout => \READ_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9836\,
            lcout => \READ_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9577\,
            lcout => \WRITE_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9839\,
            lcout => \WRITE_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9578\,
            lcout => \WRITE_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => \N__9306\,
            sr => \N__9239\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10040\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \WRITE_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9388\,
            ce => \N__9308\,
            sr => \N__9241\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10041\,
            in2 => \_gnd_net_\,
            in3 => \N__9675\,
            lcout => \WRITE_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9388\,
            ce => \N__9308\,
            sr => \N__9241\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9683\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10043\,
            lcout => \READ_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9310\,
            sr => \N__9243\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9682\,
            lcout => \READ_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9310\,
            sr => \N__9243\
        );

    \LBENn_c_sbtinv_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8015\,
            lcout => \LBENn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10014\,
            in2 => \_gnd_net_\,
            in3 => \N__9707\,
            lcout => \READ_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9406\,
            ce => \N__9298\,
            sr => \N__9230\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__6481\,
            in1 => \N__6498\,
            in2 => \_gnd_net_\,
            in3 => \N__6432\,
            lcout => \U111_CYCLE_SM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6773\,
            in1 => \N__6836\,
            in2 => \N__7155\,
            in3 => \N__6939\,
            lcout => \U111_CYCLE_SM.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6835\,
            in1 => \N__7146\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => \U111_CYCLE_SM.N_75\,
            ltout => \U111_CYCLE_SM.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__6743\,
            in1 => \N__6358\,
            in2 => \N__6371\,
            in3 => \N__7037\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6893\,
            in1 => \N__6744\,
            in2 => \_gnd_net_\,
            in3 => \N__7234\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6875\,
            in2 => \_gnd_net_\,
            in3 => \N__7081\,
            lcout => \U111_CYCLE_SM.LATCH_EN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__6334\,
            in1 => \N__6356\,
            in2 => \N__6310\,
            in3 => \N__7036\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9397\,
            ce => 'H',
            sr => \N__9237\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI541Q_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7082\,
            in2 => \_gnd_net_\,
            in3 => \N__9567\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6891\,
            in2 => \N__6362\,
            in3 => \N__6976\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9397\,
            ce => 'H',
            sr => \N__9237\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010010"
        )
    port map (
            in0 => \N__7052\,
            in1 => \N__6355\,
            in2 => \N__6980\,
            in3 => \N__6892\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9397\,
            ce => 'H',
            sr => \N__9237\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__6357\,
            in1 => \N__6335\,
            in2 => \N__6311\,
            in3 => \N__6499\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9397\,
            ce => 'H',
            sr => \N__9237\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__6874\,
            in1 => \N__7084\,
            in2 => \N__10073\,
            in3 => \N__9568\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9393\,
            ce => 'H',
            sr => \N__9240\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9819\,
            in2 => \_gnd_net_\,
            in3 => \N__9642\,
            lcout => \READ_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9648\,
            in1 => \_gnd_net_\,
            in2 => \N__9898\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9823\,
            in2 => \_gnd_net_\,
            in3 => \N__9644\,
            lcout => \READ_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9645\,
            in1 => \_gnd_net_\,
            in2 => \N__9896\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9646\,
            in1 => \_gnd_net_\,
            in2 => \N__9897\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9830\,
            in2 => \_gnd_net_\,
            in3 => \N__9647\,
            lcout => \READ_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9643\,
            in1 => \_gnd_net_\,
            in2 => \N__9895\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => \N__9309\,
            sr => \N__9242\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9698\,
            lcout => \READ_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9386\,
            ce => \N__9311\,
            sr => \N__9244\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10039\,
            in2 => \_gnd_net_\,
            in3 => \N__9699\,
            lcout => \READ_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__9312\,
            sr => \N__9245\
        );

    \D_UU_040_iobuf_RNO_6_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6404\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9158\,
            in1 => \N__6650\,
            in2 => \_gnd_net_\,
            in3 => \N__11162\,
            lcout => \un2_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6611\,
            in1 => \N__8279\,
            in2 => \_gnd_net_\,
            in3 => \N__11161\,
            lcout => \un2_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_2_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6569\,
            lcout => \N_231_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6542\,
            in1 => \N__8687\,
            in2 => \_gnd_net_\,
            in3 => \N__11122\,
            lcout => \un2_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__7232\,
            in1 => \N__6506\,
            in2 => \N__6482\,
            in3 => \N__6440\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9408\,
            ce => 'H',
            sr => \N__9234\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__6433\,
            in1 => \N__7233\,
            in2 => \N__7197\,
            in3 => \N__6959\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__6745\,
            in1 => \N__6434\,
            in2 => \N__6407\,
            in3 => \N__6899\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__6770\,
            in1 => \_gnd_net_\,
            in2 => \N__6847\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__7184\,
            in1 => \N__6747\,
            in2 => \N__6947\,
            in3 => \N__6913\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6746\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6944\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_RNILNBJ_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6769\,
            in2 => \_gnd_net_\,
            in3 => \N__7035\,
            lcout => \U111_CYCLE_SM.N_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7126\,
            lcout => \U111_CYCLE_SM.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6842\,
            in2 => \N__7127\,
            in3 => \N__7189\,
            lcout => \U111_CYCLE_SM.N_40\,
            ltout => \U111_CYCLE_SM.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011111"
        )
    port map (
            in0 => \N__6749\,
            in1 => \_gnd_net_\,
            in2 => \N__6878\,
            in3 => \N__6870\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__7125\,
            in1 => \N__6841\,
            in2 => \N__6854\,
            in3 => \N__7188\,
            lcout => \U111_CYCLE_SM.N_40_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__6843\,
            in1 => \N__6771\,
            in2 => \_gnd_net_\,
            in3 => \N__7123\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110011"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__6748\,
            in2 => \N__7253\,
            in3 => \N__7246\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7235\,
            in1 => \N__6958\,
            in2 => \N__7198\,
            in3 => \N__7124\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__7083\,
            in1 => \N__9708\,
            in2 => \N__7103\,
            in3 => \N__7100\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100111111"
        )
    port map (
            in0 => \N__7051\,
            in1 => \N__7034\,
            in2 => \N__7013\,
            in3 => \N__6975\,
            lcout => \U111_CYCLE_SM.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7408\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7490\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8528\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => \N__8234\,
            sr => \N__8201\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_5_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7664\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_210_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7634\,
            in1 => \N__7606\,
            in2 => \_gnd_net_\,
            in3 => \N__11061\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10367\,
            in1 => \N__7556\,
            in2 => \_gnd_net_\,
            in3 => \N__7546\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7486\,
            in1 => \N__7442\,
            in2 => \_gnd_net_\,
            in3 => \N__10393\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7401\,
            in1 => \N__7364\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7328\,
            in1 => \N__7317\,
            in2 => \_gnd_net_\,
            in3 => \N__10395\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_1_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7262\,
            lcout => \N_206_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8033\,
            lcout => \TAn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7957\,
            in1 => \N__7931\,
            in2 => \_gnd_net_\,
            in3 => \N__11121\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11164\,
            in1 => \N__9029\,
            in2 => \_gnd_net_\,
            in3 => \N__7895\,
            lcout => \un2_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8527\,
            in1 => \N__7856\,
            in2 => \_gnd_net_\,
            in3 => \N__11165\,
            lcout => \un2_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7813\,
            in1 => \N__7772\,
            in2 => \_gnd_net_\,
            in3 => \N__11093\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8243\,
            in1 => \N__8272\,
            in2 => \_gnd_net_\,
            in3 => \N__10350\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8765\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9403\,
            ce => \N__8236\,
            sr => \N__8212\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9403\,
            ce => \N__8236\,
            sr => \N__8212\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9403\,
            ce => \N__8236\,
            sr => \N__8212\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9090\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__8235\,
            sr => \N__8211\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8372\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8456\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8164\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9024\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10472\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => \N__8237\,
            sr => \N__8213\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8163\,
            in1 => \N__8123\,
            in2 => \_gnd_net_\,
            in3 => \N__10380\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10403\,
            in1 => \N__8834\,
            in2 => \_gnd_net_\,
            in3 => \N__8824\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10405\,
            in1 => \N__8774\,
            in2 => \_gnd_net_\,
            in3 => \N__8760\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8686\,
            in1 => \N__8645\,
            in2 => \_gnd_net_\,
            in3 => \N__10404\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11167\,
            in1 => \N__8618\,
            in2 => \_gnd_net_\,
            in3 => \N__8596\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10407\,
            in1 => \N__8540\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8448\,
            in1 => \N__8408\,
            in2 => \_gnd_net_\,
            in3 => \N__10408\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10409\,
            in1 => \N__8381\,
            in2 => \_gnd_net_\,
            in3 => \N__8371\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9038\,
            lcout => \N_224_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10327\,
            in1 => \N__9164\,
            in2 => \_gnd_net_\,
            in3 => \N__9145\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__9094\,
            in2 => \_gnd_net_\,
            in3 => \N__10379\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9701\,
            in1 => \_gnd_net_\,
            in2 => \N__10011\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9399\,
            ce => \N__9313\,
            sr => \N__9246\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9939\,
            in2 => \_gnd_net_\,
            in3 => \N__9700\,
            lcout => \READ_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9399\,
            ce => \N__9313\,
            sr => \N__9246\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9702\,
            in1 => \_gnd_net_\,
            in2 => \N__10012\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9399\,
            ce => \N__9313\,
            sr => \N__9246\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9703\,
            in1 => \_gnd_net_\,
            in2 => \N__10013\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep31_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9399\,
            ce => \N__9313\,
            sr => \N__9246\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9025\,
            in1 => \N__8978\,
            in2 => \_gnd_net_\,
            in3 => \N__10381\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_3_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8951\,
            lcout => \N_216_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8920\,
            in1 => \N__8879\,
            in2 => \_gnd_net_\,
            in3 => \N__11168\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10461\,
            in1 => \N__10421\,
            in2 => \_gnd_net_\,
            in3 => \N__10406\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_6_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_219_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_7_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \N_220_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_5_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10208\,
            lcout => \N_234_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10174\,
            in1 => \N__10133\,
            in2 => \_gnd_net_\,
            in3 => \N__11129\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \_gnd_net_\,
            in3 => \N__9704\,
            lcout => \READ_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9407\,
            ce => \N__9314\,
            sr => \N__9247\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9705\,
            in1 => \_gnd_net_\,
            in2 => \N__9938\,
            in3 => \_gnd_net_\,
            lcout => \READ_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9407\,
            ce => \N__9314\,
            sr => \N__9247\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9864\,
            in2 => \_gnd_net_\,
            in3 => \N__9706\,
            lcout => \READ_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9407\,
            ce => \N__9314\,
            sr => \N__9247\
        );

    \D_LL_040_iobuf_RNO_3_LC_17_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_232_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_2_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10760\,
            lcout => \N_223_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_0_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10730\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_7_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10694\,
            lcout => \N_212_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10661\,
            in1 => \N__10639\,
            in2 => \_gnd_net_\,
            in3 => \N__11151\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_7_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_236_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_6_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_227_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_5_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10538\,
            lcout => \N_218_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_4_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10505\,
            lcout => \N_209_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11504\,
            in1 => \N__11482\,
            in2 => \_gnd_net_\,
            in3 => \N__11169\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_4_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_233_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_6_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_235_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_1_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_222_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11321\,
            in1 => \N__11302\,
            in2 => \_gnd_net_\,
            in3 => \N__11170\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11224\,
            in1 => \N__11189\,
            in2 => \_gnd_net_\,
            in3 => \N__11171\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_1_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_230_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_2_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10814\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_5_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_226_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_0_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11726\,
            lcout => \N_229_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_1_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_214_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_4_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11657\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_0_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11621\,
            lcout => \N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_7_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11591\,
            lcout => \N_228_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_4_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11561\,
            lcout => \N_225_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_3_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_208_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_0_LC_24_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11783\,
            lcout => \N_221_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

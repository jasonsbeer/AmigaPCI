-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 23 2024 17:07:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10049\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_172_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_187\ : std_logic;
signal \U712_REG_SM.N_173_0\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_66_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_92_cascade_\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_0\ : std_logic;
signal \U712_REG_SM.N_157_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_157_0\ : std_logic;
signal \U712_REG_SM.N_159_0_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_161_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_195\ : std_logic;
signal \U712_REG_SM.N_172_0\ : std_logic;
signal \U712_REG_SM.N_195_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.DS_EN_7_0\ : std_logic;
signal \U712_REG_SM.N_163_0\ : std_logic;
signal \U712_REG_SM.N_162_0\ : std_logic;
signal \U712_REG_SM.N_181\ : std_logic;
signal \U712_REG_SM.N_170_0_cascade_\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\ : std_logic;
signal \U712_CHIP_RAM.N_67_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_66_1\ : std_logic;
signal \U712_CHIP_RAM.N_58_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_170_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_159_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_START_2_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_169_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_167_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_161_0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_186_0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH6lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH6lt7\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_54_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_59\ : std_logic;
signal \U712_CHIP_RAM.N_59_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_74_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_tz_0\ : std_logic;
signal \U712_CHIP_RAM.N_81_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_92\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a3_0_1_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_55\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER46\ : std_logic;
signal \U712_CHIP_RAM.N_55_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_89\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_56\ : std_logic;
signal \U712_CHIP_RAM.N_43_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_54\ : std_logic;
signal \U712_CHIP_RAM.N_61\ : std_logic;
signal \U712_CHIP_RAM.N_60\ : std_logic;
signal \U712_CHIP_RAM.N_61_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_42\ : std_logic;
signal \U712_CHIP_RAM.N_13\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \N_517_i\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \U712_CHIP_RAM.REF_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.N_84\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_76_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_41_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_74\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\ : std_logic;
signal \U712_CHIP_RAM.N_88\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.N_77_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_58\ : std_logic;
signal \U712_CHIP_RAM.N_44\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_75\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_35\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE.LMBE_0\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DRDDIR_0_i\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_32\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.UMBE_0\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_4\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_31\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.REF_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_7\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE_0\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.N_38\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_34\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U712_CHIP_RAM.N_50_i_0_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3568\,
            RESETB => \N__6325\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10049\,
            DIN => \N__10048\,
            DOUT => \N__10047\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10049\,
            PADOUT => \N__10048\,
            PADIN => \N__10047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10040\,
            DIN => \N__10039\,
            DOUT => \N__10038\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10040\,
            PADOUT => \N__10039\,
            PADIN => \N__10038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10031\,
            DIN => \N__10030\,
            DOUT => \N__10029\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10031\,
            PADOUT => \N__10030\,
            PADIN => \N__10029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8689\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10022\,
            DIN => \N__10021\,
            DOUT => \N__10020\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10022\,
            PADOUT => \N__10021\,
            PADIN => \N__10020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6805\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10013\,
            DIN => \N__10012\,
            DOUT => \N__10011\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10013\,
            PADOUT => \N__10012\,
            PADIN => \N__10011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10004\,
            DIN => \N__10003\,
            DOUT => \N__10002\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10004\,
            PADOUT => \N__10003\,
            PADIN => \N__10002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9995\,
            DIN => \N__9994\,
            DOUT => \N__9993\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9995\,
            PADOUT => \N__9994\,
            PADIN => \N__9993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9986\,
            DIN => \N__9985\,
            DOUT => \N__9984\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9986\,
            PADOUT => \N__9985\,
            PADIN => \N__9984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9977\,
            DIN => \N__9976\,
            DOUT => \N__9975\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9977\,
            PADOUT => \N__9976\,
            PADIN => \N__9975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9968\,
            DIN => \N__9967\,
            DOUT => \N__9966\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9968\,
            PADOUT => \N__9967\,
            PADIN => \N__9966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9959\,
            DIN => \N__9958\,
            DOUT => \N__9957\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9959\,
            PADOUT => \N__9958\,
            PADIN => \N__9957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9950\,
            DIN => \N__9949\,
            DOUT => \N__9948\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9950\,
            PADOUT => \N__9949\,
            PADIN => \N__9948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3951\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9941\,
            DIN => \N__9940\,
            DOUT => \N__9939\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9941\,
            PADOUT => \N__9940\,
            PADIN => \N__9939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9932\,
            DIN => \N__9931\,
            DOUT => \N__9930\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9932\,
            PADOUT => \N__9931\,
            PADIN => \N__9930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9923\,
            DIN => \N__9922\,
            DOUT => \N__9921\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9923\,
            PADOUT => \N__9922\,
            PADIN => \N__9921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9914\,
            DIN => \N__9913\,
            DOUT => \N__9912\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9914\,
            PADOUT => \N__9913\,
            PADIN => \N__9912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9905\,
            DIN => \N__9904\,
            DOUT => \N__9903\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9905\,
            PADOUT => \N__9904\,
            PADIN => \N__9903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9896\,
            DIN => \N__9895\,
            DOUT => \N__9894\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9896\,
            PADOUT => \N__9895\,
            PADIN => \N__9894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7576\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9887\,
            DIN => \N__9886\,
            DOUT => \N__9885\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9887\,
            PADOUT => \N__9886\,
            PADIN => \N__9885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9878\,
            DIN => \N__9877\,
            DOUT => \N__9876\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9878\,
            PADOUT => \N__9877\,
            PADIN => \N__9876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8602\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9869\,
            DIN => \N__9868\,
            DOUT => \N__9867\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9869\,
            PADOUT => \N__9868\,
            PADIN => \N__9867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9860\,
            DIN => \N__9859\,
            DOUT => \N__9858\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9860\,
            PADOUT => \N__9859\,
            PADIN => \N__9858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9851\,
            DIN => \N__9850\,
            DOUT => \N__9849\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9851\,
            PADOUT => \N__9850\,
            PADIN => \N__9849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9842\,
            DIN => \N__9841\,
            DOUT => \N__9840\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9842\,
            PADOUT => \N__9841\,
            PADIN => \N__9840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9833\,
            DIN => \N__9832\,
            DOUT => \N__9831\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9833\,
            PADOUT => \N__9832\,
            PADIN => \N__9831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9824\,
            DIN => \N__9823\,
            DOUT => \N__9822\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9824\,
            PADOUT => \N__9823\,
            PADIN => \N__9822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9815\,
            DIN => \N__9814\,
            DOUT => \N__9813\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9815\,
            PADOUT => \N__9814\,
            PADIN => \N__9813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9806\,
            DIN => \N__9805\,
            DOUT => \N__9804\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9806\,
            PADOUT => \N__9805\,
            PADIN => \N__9804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9797\,
            DIN => \N__9796\,
            DOUT => \N__9795\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9797\,
            PADOUT => \N__9796\,
            PADIN => \N__9795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9788\,
            DIN => \N__9787\,
            DOUT => \N__9786\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9788\,
            PADOUT => \N__9787\,
            PADIN => \N__9786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9779\,
            DIN => \N__9778\,
            DOUT => \N__9777\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9779\,
            PADOUT => \N__9778\,
            PADIN => \N__9777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9770\,
            DIN => \N__9769\,
            DOUT => \N__9768\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9770\,
            PADOUT => \N__9769\,
            PADIN => \N__9768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7036\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9761\,
            DIN => \N__9760\,
            DOUT => \N__9759\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9761\,
            PADOUT => \N__9760\,
            PADIN => \N__9759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9752\,
            DIN => \N__9751\,
            DOUT => \N__9750\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9752\,
            PADOUT => \N__9751\,
            PADIN => \N__9750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9743\,
            DIN => \N__9742\,
            DOUT => \N__9741\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9743\,
            PADOUT => \N__9742\,
            PADIN => \N__9741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9734\,
            DIN => \N__9733\,
            DOUT => \N__9732\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9734\,
            PADOUT => \N__9733\,
            PADIN => \N__9732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9725\,
            DIN => \N__9724\,
            DOUT => \N__9723\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9725\,
            PADOUT => \N__9724\,
            PADIN => \N__9723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3604\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9716\,
            DIN => \N__9715\,
            DOUT => \N__9714\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9716\,
            PADOUT => \N__9715\,
            PADIN => \N__9714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5158\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9707\,
            DIN => \N__9706\,
            DOUT => \N__9705\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9707\,
            PADOUT => \N__9706\,
            PADIN => \N__9705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9698\,
            DIN => \N__9697\,
            DOUT => \N__9696\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9698\,
            PADOUT => \N__9697\,
            PADIN => \N__9696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9689\,
            DIN => \N__9688\,
            DOUT => \N__9687\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9689\,
            PADOUT => \N__9688\,
            PADIN => \N__9687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9680\,
            DIN => \N__9679\,
            DOUT => \N__9678\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9680\,
            PADOUT => \N__9679\,
            PADIN => \N__9678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9671\,
            DIN => \N__9670\,
            DOUT => \N__9669\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9671\,
            PADOUT => \N__9670\,
            PADIN => \N__9669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3619\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9662\,
            DIN => \N__9661\,
            DOUT => \N__9660\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9662\,
            PADOUT => \N__9661\,
            PADIN => \N__9660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9653\,
            DIN => \N__9652\,
            DOUT => \N__9651\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9653\,
            PADOUT => \N__9652\,
            PADIN => \N__9651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4636\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9644\,
            DIN => \N__9643\,
            DOUT => \N__9642\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9644\,
            PADOUT => \N__9643\,
            PADIN => \N__9642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9635\,
            DIN => \N__9634\,
            DOUT => \N__9633\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9635\,
            PADOUT => \N__9634\,
            PADIN => \N__9633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9626\,
            DIN => \N__9625\,
            DOUT => \N__9624\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9626\,
            PADOUT => \N__9625\,
            PADIN => \N__9624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9617\,
            DIN => \N__9616\,
            DOUT => \N__9615\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9617\,
            PADOUT => \N__9616\,
            PADIN => \N__9615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9608\,
            DIN => \N__9607\,
            DOUT => \N__9606\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9608\,
            PADOUT => \N__9607\,
            PADIN => \N__9606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7015\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9599\,
            DIN => \N__9598\,
            DOUT => \N__9597\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9599\,
            PADOUT => \N__9598\,
            PADIN => \N__9597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9590\,
            DIN => \N__9589\,
            DOUT => \N__9588\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9590\,
            PADOUT => \N__9589\,
            PADIN => \N__9588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9581\,
            DIN => \N__9580\,
            DOUT => \N__9579\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9581\,
            PADOUT => \N__9580\,
            PADIN => \N__9579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9572\,
            DIN => \N__9571\,
            DOUT => \N__9570\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9572\,
            PADOUT => \N__9571\,
            PADIN => \N__9570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6343\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9563\,
            DIN => \N__9562\,
            DOUT => \N__9561\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9563\,
            PADOUT => \N__9562\,
            PADIN => \N__9561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9554\,
            DIN => \N__9553\,
            DOUT => \N__9552\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9554\,
            PADOUT => \N__9553\,
            PADIN => \N__9552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4635\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9545\,
            DIN => \N__9544\,
            DOUT => \N__9543\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9545\,
            PADOUT => \N__9544\,
            PADIN => \N__9543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9536\,
            DIN => \N__9535\,
            DOUT => \N__9534\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9536\,
            PADOUT => \N__9535\,
            PADIN => \N__9534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9527\,
            DIN => \N__9526\,
            DOUT => \N__9525\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9527\,
            PADOUT => \N__9526\,
            PADIN => \N__9525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6931\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9518\,
            DIN => \N__9517\,
            DOUT => \N__9516\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9518\,
            PADOUT => \N__9517\,
            PADIN => \N__9516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9509\,
            DIN => \N__9508\,
            DOUT => \N__9507\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9509\,
            PADOUT => \N__9508\,
            PADIN => \N__9507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6907\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9500\,
            DIN => \N__9499\,
            DOUT => \N__9498\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9500\,
            PADOUT => \N__9499\,
            PADIN => \N__9498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7360\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9491\,
            DIN => \N__9490\,
            DOUT => \N__9489\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9491\,
            PADOUT => \N__9490\,
            PADIN => \N__9489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9482\,
            DIN => \N__9481\,
            DOUT => \N__9480\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9482\,
            PADOUT => \N__9481\,
            PADIN => \N__9480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9473\,
            DIN => \N__9472\,
            DOUT => \N__9471\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9473\,
            PADOUT => \N__9472\,
            PADIN => \N__9471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9464\,
            DIN => \N__9463\,
            DOUT => \N__9462\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9464\,
            PADOUT => \N__9463\,
            PADIN => \N__9462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9455\,
            DIN => \N__9454\,
            DOUT => \N__9453\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9455\,
            PADOUT => \N__9454\,
            PADIN => \N__9453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9446\,
            DIN => \N__9445\,
            DOUT => \N__9444\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9446\,
            PADOUT => \N__9445\,
            PADIN => \N__9444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9437\,
            DIN => \N__9436\,
            DOUT => \N__9435\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9437\,
            PADOUT => \N__9436\,
            PADIN => \N__9435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8854\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9428\,
            DIN => \N__9427\,
            DOUT => \N__9426\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9428\,
            PADOUT => \N__9427\,
            PADIN => \N__9426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5794\,
            DIN0 => OPEN,
            DOUT0 => \N__3745\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9419\,
            DIN => \N__9418\,
            DOUT => \N__9417\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9419\,
            PADOUT => \N__9418\,
            PADIN => \N__9417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9410\,
            DIN => \N__9409\,
            DOUT => \N__9408\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9410\,
            PADOUT => \N__9409\,
            PADIN => \N__9408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9401\,
            DIN => \N__9400\,
            DOUT => \N__9399\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9401\,
            PADOUT => \N__9400\,
            PADIN => \N__9399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9392\,
            DIN => \N__9391\,
            DOUT => \N__9390\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9392\,
            PADOUT => \N__9391\,
            PADIN => \N__9390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9383\,
            DIN => \N__9382\,
            DOUT => \N__9381\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9383\,
            PADOUT => \N__9382\,
            PADIN => \N__9381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9374\,
            DIN => \N__9373\,
            DOUT => \N__9372\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9374\,
            PADOUT => \N__9373\,
            PADIN => \N__9372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9365\,
            DIN => \N__9364\,
            DOUT => \N__9363\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9365\,
            PADOUT => \N__9364\,
            PADIN => \N__9363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9356\,
            DIN => \N__9355\,
            DOUT => \N__9354\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9356\,
            PADOUT => \N__9355\,
            PADIN => \N__9354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9347\,
            DIN => \N__9346\,
            DOUT => \N__9345\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9347\,
            PADOUT => \N__9346\,
            PADIN => \N__9345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7474\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9338\,
            DIN => \N__9337\,
            DOUT => \N__9336\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9338\,
            PADOUT => \N__9337\,
            PADIN => \N__9336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2223\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9315\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9312\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9309\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9306\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__9309\,
            I => \N__9303\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__9306\,
            I => \N__9300\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__9303\,
            I => \N__9297\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__9300\,
            I => \N__9294\
        );

    \I__2215\ : Sp12to4
    port map (
            O => \N__9297\,
            I => \N__9289\
        );

    \I__2214\ : Sp12to4
    port map (
            O => \N__9294\,
            I => \N__9289\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__9289\,
            I => \DRA_c_8\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__9286\,
            I => \N__9283\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9280\,
            I => \N__9277\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__9277\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9271\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9261\
        );

    \I__2206\ : ClkMux
    port map (
            O => \N__9270\,
            I => \N__9142\
        );

    \I__2205\ : ClkMux
    port map (
            O => \N__9269\,
            I => \N__9142\
        );

    \I__2204\ : ClkMux
    port map (
            O => \N__9268\,
            I => \N__9142\
        );

    \I__2203\ : ClkMux
    port map (
            O => \N__9267\,
            I => \N__9142\
        );

    \I__2202\ : ClkMux
    port map (
            O => \N__9266\,
            I => \N__9142\
        );

    \I__2201\ : ClkMux
    port map (
            O => \N__9265\,
            I => \N__9142\
        );

    \I__2200\ : ClkMux
    port map (
            O => \N__9264\,
            I => \N__9142\
        );

    \I__2199\ : Glb2LocalMux
    port map (
            O => \N__9261\,
            I => \N__9142\
        );

    \I__2198\ : ClkMux
    port map (
            O => \N__9260\,
            I => \N__9142\
        );

    \I__2197\ : ClkMux
    port map (
            O => \N__9259\,
            I => \N__9142\
        );

    \I__2196\ : ClkMux
    port map (
            O => \N__9258\,
            I => \N__9142\
        );

    \I__2195\ : ClkMux
    port map (
            O => \N__9257\,
            I => \N__9142\
        );

    \I__2194\ : ClkMux
    port map (
            O => \N__9256\,
            I => \N__9142\
        );

    \I__2193\ : ClkMux
    port map (
            O => \N__9255\,
            I => \N__9142\
        );

    \I__2192\ : ClkMux
    port map (
            O => \N__9254\,
            I => \N__9142\
        );

    \I__2191\ : ClkMux
    port map (
            O => \N__9253\,
            I => \N__9142\
        );

    \I__2190\ : ClkMux
    port map (
            O => \N__9252\,
            I => \N__9142\
        );

    \I__2189\ : ClkMux
    port map (
            O => \N__9251\,
            I => \N__9142\
        );

    \I__2188\ : ClkMux
    port map (
            O => \N__9250\,
            I => \N__9142\
        );

    \I__2187\ : ClkMux
    port map (
            O => \N__9249\,
            I => \N__9142\
        );

    \I__2186\ : ClkMux
    port map (
            O => \N__9248\,
            I => \N__9142\
        );

    \I__2185\ : ClkMux
    port map (
            O => \N__9247\,
            I => \N__9142\
        );

    \I__2184\ : ClkMux
    port map (
            O => \N__9246\,
            I => \N__9142\
        );

    \I__2183\ : ClkMux
    port map (
            O => \N__9245\,
            I => \N__9142\
        );

    \I__2182\ : ClkMux
    port map (
            O => \N__9244\,
            I => \N__9142\
        );

    \I__2181\ : ClkMux
    port map (
            O => \N__9243\,
            I => \N__9142\
        );

    \I__2180\ : ClkMux
    port map (
            O => \N__9242\,
            I => \N__9142\
        );

    \I__2179\ : ClkMux
    port map (
            O => \N__9241\,
            I => \N__9142\
        );

    \I__2178\ : ClkMux
    port map (
            O => \N__9240\,
            I => \N__9142\
        );

    \I__2177\ : ClkMux
    port map (
            O => \N__9239\,
            I => \N__9142\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9238\,
            I => \N__9142\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9237\,
            I => \N__9142\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9236\,
            I => \N__9142\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9235\,
            I => \N__9142\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9234\,
            I => \N__9142\
        );

    \I__2171\ : ClkMux
    port map (
            O => \N__9233\,
            I => \N__9142\
        );

    \I__2170\ : ClkMux
    port map (
            O => \N__9232\,
            I => \N__9142\
        );

    \I__2169\ : ClkMux
    port map (
            O => \N__9231\,
            I => \N__9142\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9230\,
            I => \N__9142\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9229\,
            I => \N__9142\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9228\,
            I => \N__9142\
        );

    \I__2165\ : ClkMux
    port map (
            O => \N__9227\,
            I => \N__9142\
        );

    \I__2164\ : GlobalMux
    port map (
            O => \N__9142\,
            I => \CLK80_OUT\
        );

    \I__2163\ : CEMux
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__9136\,
            I => \N__9131\
        );

    \I__2161\ : CEMux
    port map (
            O => \N__9135\,
            I => \N__9128\
        );

    \I__2160\ : CEMux
    port map (
            O => \N__9134\,
            I => \N__9124\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9131\,
            I => \N__9121\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9128\,
            I => \N__9118\
        );

    \I__2157\ : CEMux
    port map (
            O => \N__9127\,
            I => \N__9115\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9124\,
            I => \N__9112\
        );

    \I__2155\ : Span4Mux_h
    port map (
            O => \N__9121\,
            I => \N__9109\
        );

    \I__2154\ : Span4Mux_h
    port map (
            O => \N__9118\,
            I => \N__9104\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9104\
        );

    \I__2152\ : Span4Mux_h
    port map (
            O => \N__9112\,
            I => \N__9101\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__9109\,
            I => \U712_CHIP_RAM.N_50_i_0_0\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__9104\,
            I => \U712_CHIP_RAM.N_50_i_0_0\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__9101\,
            I => \U712_CHIP_RAM.N_50_i_0_0\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9082\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9075\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9075\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9075\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9072\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9069\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9066\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9063\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9060\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9057\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9047\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9075\,
            I => \N__9044\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9072\,
            I => \N__9030\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9023\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9020\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9017\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9010\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__8998\
        );

    \I__2130\ : SRMux
    port map (
            O => \N__9056\,
            I => \N__8908\
        );

    \I__2129\ : SRMux
    port map (
            O => \N__9055\,
            I => \N__8908\
        );

    \I__2128\ : SRMux
    port map (
            O => \N__9054\,
            I => \N__8908\
        );

    \I__2127\ : SRMux
    port map (
            O => \N__9053\,
            I => \N__8908\
        );

    \I__2126\ : SRMux
    port map (
            O => \N__9052\,
            I => \N__8908\
        );

    \I__2125\ : SRMux
    port map (
            O => \N__9051\,
            I => \N__8908\
        );

    \I__2124\ : SRMux
    port map (
            O => \N__9050\,
            I => \N__8908\
        );

    \I__2123\ : Glb2LocalMux
    port map (
            O => \N__9047\,
            I => \N__8908\
        );

    \I__2122\ : Glb2LocalMux
    port map (
            O => \N__9044\,
            I => \N__8908\
        );

    \I__2121\ : SRMux
    port map (
            O => \N__9043\,
            I => \N__8908\
        );

    \I__2120\ : SRMux
    port map (
            O => \N__9042\,
            I => \N__8908\
        );

    \I__2119\ : SRMux
    port map (
            O => \N__9041\,
            I => \N__8908\
        );

    \I__2118\ : SRMux
    port map (
            O => \N__9040\,
            I => \N__8908\
        );

    \I__2117\ : SRMux
    port map (
            O => \N__9039\,
            I => \N__8908\
        );

    \I__2116\ : SRMux
    port map (
            O => \N__9038\,
            I => \N__8908\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__9037\,
            I => \N__8908\
        );

    \I__2114\ : SRMux
    port map (
            O => \N__9036\,
            I => \N__8908\
        );

    \I__2113\ : SRMux
    port map (
            O => \N__9035\,
            I => \N__8908\
        );

    \I__2112\ : SRMux
    port map (
            O => \N__9034\,
            I => \N__8908\
        );

    \I__2111\ : SRMux
    port map (
            O => \N__9033\,
            I => \N__8908\
        );

    \I__2110\ : Glb2LocalMux
    port map (
            O => \N__9030\,
            I => \N__8908\
        );

    \I__2109\ : SRMux
    port map (
            O => \N__9029\,
            I => \N__8908\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__9028\,
            I => \N__8908\
        );

    \I__2107\ : SRMux
    port map (
            O => \N__9027\,
            I => \N__8908\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__9026\,
            I => \N__8908\
        );

    \I__2105\ : Glb2LocalMux
    port map (
            O => \N__9023\,
            I => \N__8908\
        );

    \I__2104\ : Glb2LocalMux
    port map (
            O => \N__9020\,
            I => \N__8908\
        );

    \I__2103\ : Glb2LocalMux
    port map (
            O => \N__9017\,
            I => \N__8908\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__9016\,
            I => \N__8908\
        );

    \I__2101\ : SRMux
    port map (
            O => \N__9015\,
            I => \N__8908\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__9014\,
            I => \N__8908\
        );

    \I__2099\ : SRMux
    port map (
            O => \N__9013\,
            I => \N__8908\
        );

    \I__2098\ : Glb2LocalMux
    port map (
            O => \N__9010\,
            I => \N__8908\
        );

    \I__2097\ : SRMux
    port map (
            O => \N__9009\,
            I => \N__8908\
        );

    \I__2096\ : SRMux
    port map (
            O => \N__9008\,
            I => \N__8908\
        );

    \I__2095\ : SRMux
    port map (
            O => \N__9007\,
            I => \N__8908\
        );

    \I__2094\ : SRMux
    port map (
            O => \N__9006\,
            I => \N__8908\
        );

    \I__2093\ : SRMux
    port map (
            O => \N__9005\,
            I => \N__8908\
        );

    \I__2092\ : SRMux
    port map (
            O => \N__9004\,
            I => \N__8908\
        );

    \I__2091\ : SRMux
    port map (
            O => \N__9003\,
            I => \N__8908\
        );

    \I__2090\ : SRMux
    port map (
            O => \N__9002\,
            I => \N__8908\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__9001\,
            I => \N__8908\
        );

    \I__2088\ : Glb2LocalMux
    port map (
            O => \N__8998\,
            I => \N__8908\
        );

    \I__2087\ : SRMux
    port map (
            O => \N__8997\,
            I => \N__8908\
        );

    \I__2086\ : GlobalMux
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__2085\ : gio2CtrlBuf
    port map (
            O => \N__8905\,
            I => \RESETn_c_i_g\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__8902\,
            I => \N__8898\
        );

    \I__2083\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8895\
        );

    \I__2082\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8891\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8888\
        );

    \I__2080\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8885\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8882\
        );

    \I__2078\ : Span4Mux_v
    port map (
            O => \N__8888\,
            I => \N__8877\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__8885\,
            I => \N__8877\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__8882\,
            I => \N__8874\
        );

    \I__2075\ : Sp12to4
    port map (
            O => \N__8877\,
            I => \N__8871\
        );

    \I__2074\ : Sp12to4
    port map (
            O => \N__8874\,
            I => \N__8868\
        );

    \I__2073\ : Span12Mux_v
    port map (
            O => \N__8871\,
            I => \N__8865\
        );

    \I__2072\ : Span12Mux_h
    port map (
            O => \N__8868\,
            I => \N__8862\
        );

    \I__2071\ : Span12Mux_h
    port map (
            O => \N__8865\,
            I => \N__8857\
        );

    \I__2070\ : Span12Mux_v
    port map (
            O => \N__8862\,
            I => \N__8857\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__8857\,
            I => \CASUn_c\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8851\,
            I => \N__8848\
        );

    \I__2066\ : Span12Mux_s2_h
    port map (
            O => \N__8848\,
            I => \N__8845\
        );

    \I__2065\ : Span12Mux_h
    port map (
            O => \N__8845\,
            I => \N__8842\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__8842\,
            I => \CUUBEn_c\
        );

    \I__2063\ : IoInMux
    port map (
            O => \N__8839\,
            I => \N__8836\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__2061\ : IoSpan4Mux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__2060\ : IoSpan4Mux
    port map (
            O => \N__8830\,
            I => \N__8827\
        );

    \I__2059\ : Sp12to4
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__2058\ : Span12Mux_s7_h
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__2057\ : Odrv12
    port map (
            O => \N__8821\,
            I => \WEn_c\
        );

    \I__2056\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8806\
        );

    \I__2055\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8803\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \N__8800\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__8815\,
            I => \N__8797\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__8814\,
            I => \N__8794\
        );

    \I__2051\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8787\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8787\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__8811\,
            I => \N__8784\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \N__8781\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__8809\,
            I => \N__8778\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8772\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8803\,
            I => \N__8772\
        );

    \I__2044\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8769\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8764\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8764\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8761\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__8792\,
            I => \N__8758\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__8787\,
            I => \N__8754\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8751\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8748\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8743\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8743\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__8772\,
            I => \N__8734\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8769\,
            I => \N__8734\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8734\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8734\
        );

    \I__2030\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8729\
        );

    \I__2029\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8726\
        );

    \I__2028\ : Span4Mux_h
    port map (
            O => \N__8754\,
            I => \N__8723\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8720\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8715\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8743\,
            I => \N__8715\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__8734\,
            I => \N__8712\
        );

    \I__2023\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8707\
        );

    \I__2022\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8707\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8729\,
            I => \N__8704\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8726\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__8723\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__8720\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__8715\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__8712\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__8707\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__8704\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2013\ : IoInMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__2011\ : Span4Mux_s3_v
    port map (
            O => \N__8683\,
            I => \N__8680\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__8680\,
            I => \N__8677\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__8677\,
            I => \N__8674\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__8674\,
            I => \CASn_c\
        );

    \I__2007\ : IoInMux
    port map (
            O => \N__8671\,
            I => \N__8668\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8668\,
            I => \N__8665\
        );

    \I__2005\ : IoSpan4Mux
    port map (
            O => \N__8665\,
            I => \N__8662\
        );

    \I__2004\ : Span4Mux_s0_v
    port map (
            O => \N__8662\,
            I => \N__8659\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__8659\,
            I => \N__8656\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__8656\,
            I => \N__8653\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__8653\,
            I => \RASn_c\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8645\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8642\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__8648\,
            I => \N__8638\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8635\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8632\
        );

    \I__1995\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8628\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8625\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__8635\,
            I => \N__8622\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__8632\,
            I => \N__8619\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8616\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8628\,
            I => \N__8613\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8625\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8622\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__8619\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8616\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__8613\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1984\ : IoInMux
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1982\ : Span12Mux_s8_v
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__8593\,
            I => \CRCSn_c\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8587\,
            I => \U712_CHIP_RAM.N_38\
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1976\ : IoSpan4Mux
    port map (
            O => \N__8578\,
            I => \N__8575\
        );

    \I__1975\ : Span4Mux_s3_h
    port map (
            O => \N__8575\,
            I => \N__8572\
        );

    \I__1974\ : Sp12to4
    port map (
            O => \N__8572\,
            I => \N__8569\
        );

    \I__1973\ : Span12Mux_h
    port map (
            O => \N__8569\,
            I => \N__8566\
        );

    \I__1972\ : Odrv12
    port map (
            O => \N__8566\,
            I => \CMA_c_7\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8560\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__1969\ : Sp12to4
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1968\ : Span12Mux_v
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1967\ : Span12Mux_h
    port map (
            O => \N__8551\,
            I => \N__8548\
        );

    \I__1966\ : Odrv12
    port map (
            O => \N__8548\,
            I => \A_c_17\
        );

    \I__1965\ : IoInMux
    port map (
            O => \N__8545\,
            I => \N__8542\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8542\,
            I => \N__8539\
        );

    \I__1963\ : Span4Mux_s2_h
    port map (
            O => \N__8539\,
            I => \N__8536\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__8536\,
            I => \N__8533\
        );

    \I__1961\ : Sp12to4
    port map (
            O => \N__8533\,
            I => \N__8530\
        );

    \I__1960\ : Span12Mux_h
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__8527\,
            I => \CMA_c_8\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8520\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8517\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8511\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8517\,
            I => \N__8511\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8508\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__8511\,
            I => \N__8503\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8503\
        );

    \I__1951\ : Sp12to4
    port map (
            O => \N__8503\,
            I => \N__8500\
        );

    \I__1950\ : Span12Mux_v
    port map (
            O => \N__8500\,
            I => \N__8497\
        );

    \I__1949\ : Span12Mux_h
    port map (
            O => \N__8497\,
            I => \N__8494\
        );

    \I__1948\ : Odrv12
    port map (
            O => \N__8494\,
            I => \RAS0n_c\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8485\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8485\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__8485\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8476\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8476\,
            I => \N__8473\
        );

    \I__1941\ : Sp12to4
    port map (
            O => \N__8473\,
            I => \N__8470\
        );

    \I__1940\ : Span12Mux_v
    port map (
            O => \N__8470\,
            I => \N__8467\
        );

    \I__1939\ : Span12Mux_h
    port map (
            O => \N__8467\,
            I => \N__8464\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__8464\,
            I => \A_c_19\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__8461\,
            I => \N__8456\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__8460\,
            I => \N__8451\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8438\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8438\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8438\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8438\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8435\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8432\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__8449\,
            I => \N__8428\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__8448\,
            I => \N__8424\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__8447\,
            I => \N__8417\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8410\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8435\,
            I => \N__8410\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8407\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8404\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8401\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8398\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8395\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8392\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8385\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8385\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8385\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8382\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__8416\,
            I => \N__8373\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8366\
        );

    \I__1912\ : Span4Mux_h
    port map (
            O => \N__8410\,
            I => \N__8363\
        );

    \I__1911\ : Span4Mux_h
    port map (
            O => \N__8407\,
            I => \N__8346\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8346\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8346\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8398\,
            I => \N__8346\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8395\,
            I => \N__8346\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8392\,
            I => \N__8346\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8346\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8346\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8341\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8341\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8338\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8329\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8329\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8329\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8329\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8326\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8321\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8321\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8318\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8315\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__8363\,
            I => \N__8312\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__8346\,
            I => \N__8309\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8302\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8302\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8302\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8326\,
            I => \CPU_CYCLEm\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8321\,
            I => \CPU_CYCLEm\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8318\,
            I => \CPU_CYCLEm\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__8315\,
            I => \CPU_CYCLEm\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__8312\,
            I => \CPU_CYCLEm\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__8309\,
            I => \CPU_CYCLEm\
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__8302\,
            I => \CPU_CYCLEm\
        );

    \I__1879\ : IoInMux
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1877\ : IoSpan4Mux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1876\ : IoSpan4Mux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1875\ : Span4Mux_s0_h
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1874\ : Sp12to4
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1873\ : Odrv12
    port map (
            O => \N__8269\,
            I => \CMA_c_9\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8256\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8253\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8250\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8244\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8241\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8234\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8234\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8234\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8256\,
            I => \N__8231\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8253\,
            I => \N__8226\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8226\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8223\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8216\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8247\,
            I => \N__8216\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8244\,
            I => \N__8211\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8241\,
            I => \N__8211\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8208\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__8231\,
            I => \N__8201\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__8226\,
            I => \N__8201\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8201\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8197\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8194\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8191\
        );

    \I__1849\ : Span4Mux_h
    port map (
            O => \N__8211\,
            I => \N__8184\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__8208\,
            I => \N__8184\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__8201\,
            I => \N__8184\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8181\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8178\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8194\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8191\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8184\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__8178\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__8161\,
            I => \U712_CHIP_RAM.N_34\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \N__8150\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__8157\,
            I => \N__8147\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8143\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8136\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8132\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8129\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8126\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8121\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8121\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8143\,
            I => \N__8118\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8142\,
            I => \N__8115\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8108\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8108\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8105\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8136\,
            I => \N__8102\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8099\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8132\,
            I => \N__8096\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8129\,
            I => \N__8093\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8084\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8084\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__8118\,
            I => \N__8084\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8084\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8081\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8078\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8075\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8070\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__8102\,
            I => \N__8070\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8099\,
            I => \N__8061\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__8096\,
            I => \N__8061\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__8093\,
            I => \N__8061\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8084\,
            I => \N__8061\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8058\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8078\,
            I => \N__8055\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__8075\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__8070\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__8061\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8058\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__8055\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1798\ : IoInMux
    port map (
            O => \N__8044\,
            I => \N__8041\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8038\
        );

    \I__1796\ : Span4Mux_s1_h
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1794\ : Span12Mux_s8_v
    port map (
            O => \N__8032\,
            I => \N__8029\
        );

    \I__1793\ : Span12Mux_h
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__8026\,
            I => \CMA_c_3\
        );

    \I__1791\ : CEMux
    port map (
            O => \N__8023\,
            I => \N__8015\
        );

    \I__1790\ : CEMux
    port map (
            O => \N__8022\,
            I => \N__8012\
        );

    \I__1789\ : CEMux
    port map (
            O => \N__8021\,
            I => \N__8009\
        );

    \I__1788\ : CEMux
    port map (
            O => \N__8020\,
            I => \N__8006\
        );

    \I__1787\ : CEMux
    port map (
            O => \N__8019\,
            I => \N__8003\
        );

    \I__1786\ : CEMux
    port map (
            O => \N__8018\,
            I => \N__8000\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__7997\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8012\,
            I => \N__7992\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__7992\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8006\,
            I => \N__7989\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8003\,
            I => \N__7986\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8000\,
            I => \N__7979\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__7997\,
            I => \N__7979\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__7992\,
            I => \N__7979\
        );

    \I__1777\ : Span4Mux_h
    port map (
            O => \N__7989\,
            I => \N__7976\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__7986\,
            I => \N__7973\
        );

    \I__1775\ : Sp12to4
    port map (
            O => \N__7979\,
            I => \N__7970\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__7976\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__7973\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__7970\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7960\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__7960\,
            I => \N__7956\
        );

    \I__1769\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7953\
        );

    \I__1768\ : Sp12to4
    port map (
            O => \N__7956\,
            I => \N__7948\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7948\
        );

    \I__1766\ : Span12Mux_v
    port map (
            O => \N__7948\,
            I => \N__7945\
        );

    \I__1765\ : Span12Mux_h
    port map (
            O => \N__7945\,
            I => \N__7942\
        );

    \I__1764\ : Odrv12
    port map (
            O => \N__7942\,
            I => \RAS1n_c\
        );

    \I__1763\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7935\
        );

    \I__1762\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7932\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__7935\,
            I => \N__7927\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7927\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__7927\,
            I => \U712_CHIP_RAM.REF_SYNCZ0Z_0\
        );

    \I__1758\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7921\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__7921\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_7\
        );

    \I__1756\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7915\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__1754\ : Span12Mux_v
    port map (
            O => \N__7912\,
            I => \N__7909\
        );

    \I__1753\ : Span12Mux_h
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__7906\,
            I => \A_c_18\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1749\ : Span12Mux_v
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__1748\ : Span12Mux_h
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1747\ : Odrv12
    port map (
            O => \N__7891\,
            I => \A_c_16\
        );

    \I__1746\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7884\
        );

    \I__1745\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7881\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__7884\,
            I => \N__7878\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7875\
        );

    \I__1742\ : Sp12to4
    port map (
            O => \N__7878\,
            I => \N__7872\
        );

    \I__1741\ : Span12Mux_h
    port map (
            O => \N__7875\,
            I => \N__7869\
        );

    \I__1740\ : Span12Mux_v
    port map (
            O => \N__7872\,
            I => \N__7866\
        );

    \I__1739\ : Span12Mux_v
    port map (
            O => \N__7869\,
            I => \N__7861\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__7866\,
            I => \N__7861\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__7861\,
            I => \DRA_c_2\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__7849\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7842\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7839\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7842\,
            I => \N__7834\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7839\,
            I => \N__7834\
        );

    \I__1728\ : Sp12to4
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__1727\ : Span12Mux_v
    port map (
            O => \N__7831\,
            I => \N__7828\
        );

    \I__1726\ : Span12Mux_h
    port map (
            O => \N__7828\,
            I => \N__7825\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__7825\,
            I => \DRA_c_5\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7819\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7819\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1722\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7812\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7809\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7812\,
            I => \N__7806\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7803\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__7806\,
            I => \N__7800\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__7803\,
            I => \N__7797\
        );

    \I__1716\ : Sp12to4
    port map (
            O => \N__7800\,
            I => \N__7792\
        );

    \I__1715\ : Sp12to4
    port map (
            O => \N__7797\,
            I => \N__7792\
        );

    \I__1714\ : Span12Mux_h
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__1713\ : Span12Mux_v
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__7786\,
            I => \DRA_c_4\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7780\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7780\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7774\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7774\,
            I => \N__7770\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7767\
        );

    \I__1706\ : Span12Mux_v
    port map (
            O => \N__7770\,
            I => \N__7764\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__7767\,
            I => \N__7761\
        );

    \I__1704\ : Span12Mux_v
    port map (
            O => \N__7764\,
            I => \N__7758\
        );

    \I__1703\ : Span12Mux_h
    port map (
            O => \N__7761\,
            I => \N__7755\
        );

    \I__1702\ : Span12Mux_h
    port map (
            O => \N__7758\,
            I => \N__7752\
        );

    \I__1701\ : Span12Mux_v
    port map (
            O => \N__7755\,
            I => \N__7749\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__7752\,
            I => \DRA_c_1\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__7749\,
            I => \DRA_c_1\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7741\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7741\,
            I => \N__7738\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__7738\,
            I => \N__7735\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__7735\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7729\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__7729\,
            I => \N__7725\
        );

    \I__1692\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7722\
        );

    \I__1691\ : Sp12to4
    port map (
            O => \N__7725\,
            I => \N__7717\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7717\
        );

    \I__1689\ : Span12Mux_v
    port map (
            O => \N__7717\,
            I => \N__7714\
        );

    \I__1688\ : Span12Mux_h
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__7711\,
            I => \DRA_c_3\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7705\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7702\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__7702\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7693\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__7693\,
            I => \N__7690\
        );

    \I__1680\ : Span4Mux_h
    port map (
            O => \N__7690\,
            I => \N__7687\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__7687\,
            I => \U712_BYTE_ENABLE.UUBE_0\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7681\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__7678\,
            I => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7672\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7666\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7666\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7660\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7660\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7654\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7647\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7644\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7639\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7639\
        );

    \I__1663\ : Sp12to4
    port map (
            O => \N__7639\,
            I => \N__7636\
        );

    \I__1662\ : Span12Mux_v
    port map (
            O => \N__7636\,
            I => \N__7633\
        );

    \I__1661\ : Span12Mux_h
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__1660\ : Odrv12
    port map (
            O => \N__7630\,
            I => \DRA_c_6\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7624\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7624\,
            I => \N__7621\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__7621\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7615\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7615\,
            I => \N__7611\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7608\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7611\,
            I => \N__7603\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7608\,
            I => \N__7603\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1650\ : Sp12to4
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1649\ : Span12Mux_h
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1648\ : Odrv12
    port map (
            O => \N__7594\,
            I => \DRA_c_7\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7588\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__7585\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7579\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7579\,
            I => \U712_CHIP_RAM.N_31\
        );

    \I__1642\ : IoInMux
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7570\
        );

    \I__1640\ : Span4Mux_s3_v
    port map (
            O => \N__7570\,
            I => \N__7567\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7567\,
            I => \N__7564\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__7558\,
            I => \CMA_c_0\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7551\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7548\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7551\,
            I => \N__7543\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7548\,
            I => \N__7543\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1630\ : Sp12to4
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__1629\ : Span12Mux_h
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1628\ : Span12Mux_v
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__7531\,
            I => \DRA_c_0\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__1624\ : Span4Mux_h
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__7519\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7513\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1620\ : CEMux
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7502\
        );

    \I__1618\ : CEMux
    port map (
            O => \N__7506\,
            I => \N__7499\
        );

    \I__1617\ : CEMux
    port map (
            O => \N__7505\,
            I => \N__7496\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__7502\,
            I => \N__7491\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7499\,
            I => \N__7491\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7488\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__7491\,
            I => \N__7485\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__7488\,
            I => \N__7482\
        );

    \I__1611\ : Span4Mux_h
    port map (
            O => \N__7485\,
            I => \N__7479\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__7482\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__7479\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1608\ : IoInMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1606\ : IoSpan4Mux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1605\ : IoSpan4Mux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1604\ : Span4Mux_s2_h
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1603\ : Sp12to4
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__7456\,
            I => \CMA_c_5\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7450\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7444\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7444\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_4\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1595\ : Sp12to4
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1594\ : Span12Mux_v
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1593\ : Span12Mux_h
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__7426\,
            I => \A_c_14\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__7423\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7417\,
            I => \N__7414\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1586\ : Sp12to4
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1585\ : Span12Mux_h
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1584\ : Odrv12
    port map (
            O => \N__7402\,
            I => \A_c_7\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7396\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7390\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7390\,
            I => \N__7387\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__7387\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7381\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7381\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7375\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7375\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7369\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__7363\,
            I => \U712_BYTE_ENABLE.UMBE_0\
        );

    \I__1570\ : IoInMux
    port map (
            O => \N__7360\,
            I => \N__7357\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1568\ : Span4Mux_s2_h
    port map (
            O => \N__7354\,
            I => \N__7351\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1566\ : Span12Mux_v
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__7345\,
            I => \N__7342\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__7342\,
            I => \CUMBEn_c\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7334\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__7338\,
            I => \N__7331\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7328\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7334\,
            I => \N__7325\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7322\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7328\,
            I => \N__7319\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__7325\,
            I => \N__7314\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7322\,
            I => \N__7314\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7319\,
            I => \N__7308\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__7314\,
            I => \N__7308\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7305\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__7308\,
            I => \REG_CYCLEm\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7305\,
            I => \REG_CYCLEm\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7292\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7292\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7289\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7286\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7292\,
            I => \N__7277\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7289\,
            I => \N__7277\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7277\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7274\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7270\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__7277\,
            I => \N__7265\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7265\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7262\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7259\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__7265\,
            I => \DMA_CYCLEm\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7262\,
            I => \DMA_CYCLEm\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__7259\,
            I => \DMA_CYCLEm\
        );

    \I__1534\ : IoInMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1532\ : Span4Mux_s1_v
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__7243\,
            I => \N__7240\
        );

    \I__1530\ : Sp12to4
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1529\ : Span12Mux_s7_h
    port map (
            O => \N__7237\,
            I => \N__7234\
        );

    \I__1528\ : Span12Mux_v
    port map (
            O => \N__7234\,
            I => \N__7231\
        );

    \I__1527\ : Odrv12
    port map (
            O => \N__7231\,
            I => \DRDENn_c\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7224\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7221\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7224\,
            I => \N__7218\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7221\,
            I => \N__7215\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__7218\,
            I => \N__7211\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7215\,
            I => \N__7208\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7205\
        );

    \I__1519\ : Sp12to4
    port map (
            O => \N__7211\,
            I => \N__7202\
        );

    \I__1518\ : Sp12to4
    port map (
            O => \N__7208\,
            I => \N__7199\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7205\,
            I => \N__7196\
        );

    \I__1516\ : Span12Mux_v
    port map (
            O => \N__7202\,
            I => \N__7193\
        );

    \I__1515\ : Span12Mux_h
    port map (
            O => \N__7199\,
            I => \N__7190\
        );

    \I__1514\ : Span12Mux_h
    port map (
            O => \N__7196\,
            I => \N__7187\
        );

    \I__1513\ : Span12Mux_h
    port map (
            O => \N__7193\,
            I => \N__7182\
        );

    \I__1512\ : Span12Mux_v
    port map (
            O => \N__7190\,
            I => \N__7182\
        );

    \I__1511\ : Span12Mux_v
    port map (
            O => \N__7187\,
            I => \N__7179\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__7182\,
            I => \CASLn_c\
        );

    \I__1509\ : Odrv12
    port map (
            O => \N__7179\,
            I => \CASLn_c\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7170\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7170\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7167\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7159\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7159\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7147\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7142\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7142\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7138\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7131\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7131\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7131\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7147\,
            I => \N__7128\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7125\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7122\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7138\,
            I => \N__7119\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7116\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__7128\,
            I => \N__7109\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__7125\,
            I => \N__7109\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7109\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__7119\,
            I => \N__7103\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__7116\,
            I => \N__7103\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__7109\,
            I => \N__7100\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7097\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7103\,
            I => \N__7094\
        );

    \I__1482\ : Sp12to4
    port map (
            O => \N__7100\,
            I => \N__7089\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7097\,
            I => \N__7089\
        );

    \I__1480\ : Sp12to4
    port map (
            O => \N__7094\,
            I => \N__7084\
        );

    \I__1479\ : Span12Mux_v
    port map (
            O => \N__7089\,
            I => \N__7084\
        );

    \I__1478\ : Span12Mux_h
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__1477\ : Odrv12
    port map (
            O => \N__7081\,
            I => \RESETn_c\
        );

    \I__1476\ : IoInMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1474\ : Span12Mux_s7_v
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1473\ : Odrv12
    port map (
            O => \N__7069\,
            I => \RESETn_c_i\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__7066\,
            I => \N__7062\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7059\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7056\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7050\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7050\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7047\
        );

    \I__1466\ : Odrv12
    port map (
            O => \N__7050\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7047\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7039\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__1462\ : IoInMux
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7033\,
            I => \N__7030\
        );

    \I__1460\ : Span4Mux_s3_h
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1458\ : Span12Mux_s8_v
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__1457\ : Span12Mux_h
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__1456\ : Odrv12
    port map (
            O => \N__7018\,
            I => \CMA_c_6\
        );

    \I__1455\ : IoInMux
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__7009\
        );

    \I__1453\ : IoSpan4Mux
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__1452\ : Sp12to4
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__1451\ : Span12Mux_s9_v
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__7000\,
            I => \CMA_c_10\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1447\ : Span12Mux_h
    port map (
            O => \N__6991\,
            I => \N__6988\
        );

    \I__1446\ : Span12Mux_v
    port map (
            O => \N__6988\,
            I => \N__6985\
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__6985\,
            I => \A_c_3\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__6976\,
            I => \N__6973\
        );

    \I__1441\ : Sp12to4
    port map (
            O => \N__6973\,
            I => \N__6970\
        );

    \I__1440\ : Span12Mux_h
    port map (
            O => \N__6970\,
            I => \N__6967\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__6967\,
            I => \A_c_10\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6958\,
            I => \N__6954\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6957\,
            I => \N__6951\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__6954\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6951\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__6946\,
            I => \N__6943\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6940\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6940\,
            I => \N__6937\
        );

    \I__1429\ : Span12Mux_h
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__1428\ : Odrv12
    port map (
            O => \N__6934\,
            I => \U712_BYTE_ENABLE.LMBE_0\
        );

    \I__1427\ : IoInMux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1425\ : IoSpan4Mux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1424\ : Span4Mux_s2_v
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1423\ : Span4Mux_v
    port map (
            O => \N__6919\,
            I => \N__6916\
        );

    \I__1422\ : Sp12to4
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1421\ : Span12Mux_h
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__6910\,
            I => \CLMBEn_c\
        );

    \I__1419\ : IoInMux
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__1417\ : Span4Mux_s2_v
    port map (
            O => \N__6901\,
            I => \N__6897\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6894\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__6897\,
            I => \N__6891\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6888\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__6891\,
            I => \N__6884\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__6888\,
            I => \N__6881\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6878\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__6884\,
            I => \DBDIR_c\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__6881\,
            I => \DBDIR_c\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6878\,
            I => \DBDIR_c\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__6871\,
            I => \N__6868\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6863\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__6867\,
            I => \N__6860\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6856\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6853\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6860\,
            I => \N__6848\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6848\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6845\
        );

    \I__1399\ : Span4Mux_v
    port map (
            O => \N__6853\,
            I => \N__6839\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6848\,
            I => \N__6839\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__6845\,
            I => \N__6836\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6833\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__6839\,
            I => \N__6830\
        );

    \I__1394\ : Sp12to4
    port map (
            O => \N__6836\,
            I => \N__6825\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6833\,
            I => \N__6825\
        );

    \I__1392\ : Sp12to4
    port map (
            O => \N__6830\,
            I => \N__6822\
        );

    \I__1391\ : Span12Mux_h
    port map (
            O => \N__6825\,
            I => \N__6819\
        );

    \I__1390\ : Span12Mux_h
    port map (
            O => \N__6822\,
            I => \N__6816\
        );

    \I__1389\ : Span12Mux_v
    port map (
            O => \N__6819\,
            I => \N__6813\
        );

    \I__1388\ : Span12Mux_v
    port map (
            O => \N__6816\,
            I => \N__6810\
        );

    \I__1387\ : Odrv12
    port map (
            O => \N__6813\,
            I => \RnW_c\
        );

    \I__1386\ : Odrv12
    port map (
            O => \N__6810\,
            I => \RnW_c\
        );

    \I__1385\ : IoInMux
    port map (
            O => \N__6805\,
            I => \N__6802\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6802\,
            I => \N__6799\
        );

    \I__1383\ : IoSpan4Mux
    port map (
            O => \N__6799\,
            I => \N__6796\
        );

    \I__1382\ : IoSpan4Mux
    port map (
            O => \N__6796\,
            I => \N__6793\
        );

    \I__1381\ : Sp12to4
    port map (
            O => \N__6793\,
            I => \N__6790\
        );

    \I__1380\ : Span12Mux_s7_h
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__1379\ : Span12Mux_v
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__6784\,
            I => \DRDDIR_0_i\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6778\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6778\,
            I => \N__6775\
        );

    \I__1375\ : Span12Mux_v
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__1374\ : Span12Mux_h
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1373\ : Odrv12
    port map (
            O => \N__6769\,
            I => \A_c_9\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__6766\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6760\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6760\,
            I => \N__6757\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__6757\,
            I => \N__6754\
        );

    \I__1368\ : Span12Mux_v
    port map (
            O => \N__6754\,
            I => \N__6751\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__6751\,
            I => \N__6748\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__6748\,
            I => \A_c_2\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6742\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6742\,
            I => \U712_CHIP_RAM.N_32\
        );

    \I__1363\ : IoInMux
    port map (
            O => \N__6739\,
            I => \N__6736\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1361\ : Span12Mux_s4_v
    port map (
            O => \N__6733\,
            I => \N__6730\
        );

    \I__1360\ : Odrv12
    port map (
            O => \N__6730\,
            I => \CMA_c_1\
        );

    \I__1359\ : IoInMux
    port map (
            O => \N__6727\,
            I => \N__6724\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6721\
        );

    \I__1357\ : Span4Mux_s1_v
    port map (
            O => \N__6721\,
            I => \N__6717\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6714\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__6717\,
            I => \N__6710\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6707\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6704\
        );

    \I__1352\ : Span4Mux_v
    port map (
            O => \N__6710\,
            I => \N__6701\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__6707\,
            I => \N__6696\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6704\,
            I => \N__6696\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__6701\,
            I => \N__6690\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__6696\,
            I => \N__6690\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6687\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6690\,
            I => \DBENn_c\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6687\,
            I => \DBENn_c\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__6682\,
            I => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0_cascade_\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1341\ : Span12Mux_s11_v
    port map (
            O => \N__6673\,
            I => \N__6670\
        );

    \I__1340\ : Span12Mux_h
    port map (
            O => \N__6670\,
            I => \N__6667\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__6667\,
            I => \A_c_11\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6658\,
            I => \N__6655\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1334\ : Sp12to4
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1333\ : Span12Mux_v
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1332\ : Span12Mux_h
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6643\,
            I => \A_c_4\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6637\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1326\ : Span12Mux_v
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1325\ : Span12Mux_h
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1324\ : Odrv12
    port map (
            O => \N__6622\,
            I => \A_c_15\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6613\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__1317\ : Span12Mux_h
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__6598\,
            I => \A_c_8\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6591\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6588\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6591\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6588\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1309\ : Span12Mux_s10_v
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1308\ : Span12Mux_h
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__6571\,
            I => \A_c_13\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1303\ : Sp12to4
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1302\ : Span12Mux_v
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__1301\ : Span12Mux_h
    port map (
            O => \N__6553\,
            I => \N__6550\
        );

    \I__1300\ : Odrv12
    port map (
            O => \N__6550\,
            I => \A_c_6\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6544\,
            I => \U712_CHIP_RAM.N_35\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6538\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6538\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_6\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6532\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6532\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__1289\ : Span12Mux_h
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__6514\,
            I => \A_c_12\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1284\ : Span12Mux_v
    port map (
            O => \N__6502\,
            I => \N__6499\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__6499\,
            I => \N__6496\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__6496\,
            I => \A_c_5\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6486\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6486\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6483\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6486\,
            I => \U712_CHIP_RAM.N_75\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6483\,
            I => \U712_CHIP_RAM.N_75\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__6472\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6459\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6456\
        );

    \I__1269\ : Span4Mux_v
    port map (
            O => \N__6459\,
            I => \N__6453\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6456\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__6453\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__6448\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6441\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6438\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6441\,
            I => \N__6434\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6438\,
            I => \N__6431\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6428\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__6434\,
            I => \N__6425\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__6431\,
            I => \N__6422\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6428\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__6425\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__6422\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__6415\,
            I => \N__6410\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__6414\,
            I => \N__6407\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6404\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6398\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6398\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6404\,
            I => \N__6395\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6392\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6389\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__6395\,
            I => \N__6386\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6392\,
            I => \N__6383\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__6389\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__6386\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__6383\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6370\,
            I => \TACK_EN_i_ess\
        );

    \I__1239\ : CEMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__6358\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6346\,
            I => \U712_BYTE_ENABLE.LLBE_0\
        );

    \I__1231\ : IoInMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1229\ : IoSpan4Mux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__1228\ : Span4Mux_s0_v
    port map (
            O => \N__6334\,
            I => \N__6331\
        );

    \I__1227\ : Sp12to4
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__6328\,
            I => \CLLBEn_c\
        );

    \I__1225\ : IoInMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1223\ : Span12Mux_s6_v
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1222\ : Odrv12
    port map (
            O => \N__6316\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1221\ : IoInMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1219\ : Span4Mux_s0_v
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1217\ : Span4Mux_v
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__6298\,
            I => \CMA_c_2\
        );

    \I__1215\ : IoInMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1213\ : IoSpan4Mux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1212\ : IoSpan4Mux
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__1211\ : Span4Mux_s3_h
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__6277\,
            I => \CMA_c_4\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6271\,
            I => \N__6263\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6260\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6255\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6255\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6252\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6266\,
            I => \N__6247\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__6263\,
            I => \N__6242\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6260\,
            I => \N__6242\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6237\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6252\,
            I => \N__6237\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__6251\,
            I => \N__6232\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6228\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6225\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__6242\,
            I => \N__6222\
        );

    \I__1193\ : Span4Mux_h
    port map (
            O => \N__6237\,
            I => \N__6219\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6214\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6214\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6209\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6209\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6228\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6225\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__6219\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6209\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6192\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6189\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6192\,
            I => \U712_CHIP_RAM.N_41_i\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6189\,
            I => \U712_CHIP_RAM.N_41_i\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6181\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6175\,
            I => \U712_CHIP_RAM.N_74\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__6172\,
            I => \N__6167\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6159\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6156\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6147\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6140\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6140\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6140\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6137\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6134\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6159\,
            I => \N__6129\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6156\,
            I => \N__6129\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6124\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6124\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6115\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6115\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6115\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6115\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6147\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6140\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6137\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6134\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6129\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6124\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6115\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6097\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6097\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6087\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6087\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6084\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6087\,
            I => \U712_CHIP_RAM.N_88\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6084\,
            I => \U712_CHIP_RAM.N_88\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6067\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6067\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6067\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6067\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6067\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6064\,
            I => \U712_CHIP_RAM.N_77_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6054\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6054\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6048\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6054\,
            I => \N__6045\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6038\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6038\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6038\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6048\,
            I => \N__6017\
        );

    \I__1129\ : Span4Mux_v
    port map (
            O => \N__6045\,
            I => \N__6012\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__6012\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6009\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6006\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6035\,
            I => \N__5999\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6034\,
            I => \N__5999\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6033\,
            I => \N__5999\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6032\,
            I => \N__5990\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6031\,
            I => \N__5990\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6030\,
            I => \N__5990\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6029\,
            I => \N__5990\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6028\,
            I => \N__5981\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6027\,
            I => \N__5981\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6026\,
            I => \N__5981\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6025\,
            I => \N__5981\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6024\,
            I => \N__5976\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6023\,
            I => \N__5976\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6022\,
            I => \N__5969\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6021\,
            I => \N__5969\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6020\,
            I => \N__5969\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__6012\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6006\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5999\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5990\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5981\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5976\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1098\ : Span4Mux_v
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__5941\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \N__5934\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5937\,
            I => \N__5931\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5928\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5925\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5928\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5925\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5916\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__5919\,
            I => \N__5912\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5905\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5897\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5897\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5897\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5890\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5885\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5885\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__5905\,
            I => \N__5882\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5879\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5876\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5871\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5871\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5866\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5866\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5890\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5885\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__5882\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5879\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__5876\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5871\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5866\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5848\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__5845\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__5842\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5836\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5836\,
            I => \N__5833\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__1060\ : Sp12to4
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__1059\ : Span12Mux_h
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__1058\ : Span12Mux_v
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1057\ : Odrv12
    port map (
            O => \N__5821\,
            I => \DBRn_c\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5813\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5810\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5807\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5804\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5801\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5807\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__5804\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__5801\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1048\ : IoInMux
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__1046\ : IoSpan4Mux
    port map (
            O => \N__5788\,
            I => \N__5785\
        );

    \I__1045\ : Span4Mux_s2_h
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__1044\ : Sp12to4
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1043\ : Span12Mux_h
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1042\ : Odrv12
    port map (
            O => \N__5776\,
            I => \N_517_i\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5770\,
            I => \N__5766\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5763\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__5766\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5763\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5754\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5751\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5754\,
            I => \N__5748\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5751\,
            I => \N__5745\
        );

    \I__1032\ : Span4Mux_v
    port map (
            O => \N__5748\,
            I => \N__5741\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__5745\,
            I => \N__5738\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5735\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__5741\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__5738\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5735\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1026\ : IoInMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__1024\ : IoSpan4Mux
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__1023\ : Span4Mux_s3_v
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__1022\ : Sp12to4
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__1021\ : Span12Mux_v
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__5710\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5704\,
            I => \U712_CHIP_RAM.REF_SYNCZ0Z_1\
        );

    \I__1017\ : SRMux
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5692\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__5683\,
            I => \U712_CHIP_RAM.N_84\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5670\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5667\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5663\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5660\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__5673\,
            I => \N__5657\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5670\,
            I => \N__5651\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5667\,
            I => \N__5651\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5648\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5645\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5642\
        );

    \I__999\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5639\
        );

    \I__998\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5636\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__5651\,
            I => \N__5631\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5631\
        );

    \I__995\ : Span4Mux_h
    port map (
            O => \N__5645\,
            I => \N__5628\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__5642\,
            I => \N__5623\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5623\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5636\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__5631\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__5628\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__5623\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__5614\,
            I => \U712_CHIP_RAM.N_76_cascade_\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__5611\,
            I => \N__5606\
        );

    \I__986\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5602\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__5609\,
            I => \N__5599\
        );

    \I__984\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5596\
        );

    \I__983\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5593\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5602\,
            I => \N__5590\
        );

    \I__981\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5587\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5596\,
            I => \N__5584\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5581\
        );

    \I__978\ : Span4Mux_v
    port map (
            O => \N__5590\,
            I => \N__5578\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__5584\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__5581\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__5578\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__973\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5566\,
            I => \U712_CHIP_RAM.N_55\
        );

    \I__971\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5553\
        );

    \I__969\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5550\
        );

    \I__968\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5543\
        );

    \I__967\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5543\
        );

    \I__966\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5543\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__5553\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5550\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__5536\,
            I => \U712_CHIP_RAM.N_55_cascade_\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \N__5529\
        );

    \I__960\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5526\
        );

    \I__959\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5523\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5526\,
            I => \N__5519\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5516\
        );

    \I__956\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5513\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__5519\,
            I => \N__5508\
        );

    \I__954\ : Span4Mux_h
    port map (
            O => \N__5516\,
            I => \N__5508\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5505\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__5508\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_a3_0\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__5505\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_a3_0\
        );

    \I__950\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5496\
        );

    \I__949\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5490\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5487\
        );

    \I__947\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5484\
        );

    \I__946\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5481\
        );

    \I__945\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5478\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5490\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__5487\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5484\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5481\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \N__5463\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__5466\,
            I => \N__5456\
        );

    \I__937\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5448\
        );

    \I__936\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5448\
        );

    \I__935\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5445\
        );

    \I__934\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5442\
        );

    \I__933\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5439\
        );

    \I__932\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5436\
        );

    \I__931\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5431\
        );

    \I__930\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5431\
        );

    \I__929\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5428\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5425\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5445\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5442\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5439\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5431\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5428\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__5425\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__920\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5406\
        );

    \I__919\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5403\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5406\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5403\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5398\,
            I => \U712_CHIP_RAM.N_43_cascade_\
        );

    \I__915\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__5394\,
            I => \N__5386\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5393\,
            I => \N__5382\
        );

    \I__912\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5378\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5375\
        );

    \I__910\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5368\
        );

    \I__909\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5368\
        );

    \I__908\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5368\
        );

    \I__907\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5365\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5378\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5368\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__902\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5353\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__900\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5343\
        );

    \I__899\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5343\
        );

    \I__898\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5340\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5343\,
            I => \U712_CHIP_RAM.N_60\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5340\,
            I => \U712_CHIP_RAM.N_60\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \U712_CHIP_RAM.N_61_cascade_\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__5332\,
            I => \N__5329\
        );

    \I__893\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5324\
        );

    \I__892\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5316\
        );

    \I__891\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5316\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5324\,
            I => \N__5313\
        );

    \I__889\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5310\
        );

    \I__888\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5307\
        );

    \I__887\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5304\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5316\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__885\ : Odrv4
    port map (
            O => \N__5313\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5310\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5307\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5304\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__5293\,
            I => \N__5288\
        );

    \I__880\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5281\
        );

    \I__879\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5281\
        );

    \I__878\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5281\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5281\,
            I => \U712_CHIP_RAM.N_13\
        );

    \I__876\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5275\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5275\,
            I => \N__5271\
        );

    \I__874\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5268\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__5271\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5268\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5263\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\
        );

    \I__870\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5257\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__867\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5247\
        );

    \I__866\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5243\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5247\,
            I => \N__5240\
        );

    \I__864\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5237\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5243\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__5240\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__860\ : IoInMux
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5224\
        );

    \I__858\ : IoSpan4Mux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__857\ : Span4Mux_s3_h
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__856\ : Span4Mux_h
    port map (
            O => \N__5218\,
            I => \N__5215\
        );

    \I__855\ : Sp12to4
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__854\ : Span12Mux_h
    port map (
            O => \N__5212\,
            I => \N__5208\
        );

    \I__853\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5205\
        );

    \I__852\ : Odrv12
    port map (
            O => \N__5208\,
            I => \CLK_EN_c\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5205\,
            I => \CLK_EN_c\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__5200\,
            I => \U712_CHIP_RAM.N_74_cascade_\
        );

    \I__849\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5194\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_tz_0\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5191\,
            I => \U712_CHIP_RAM.N_81_cascade_\
        );

    \I__846\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__5182\,
            I => \N__5179\
        );

    \I__843\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5176\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5176\,
            I => \N__5172\
        );

    \I__841\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5169\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__5172\,
            I => \N__5166\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5169\,
            I => \U712_CHIP_RAM.N_92\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5166\,
            I => \U712_CHIP_RAM.N_92\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a3_0_1_3_cascade_\
        );

    \I__836\ : IoInMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__834\ : Span4Mux_s3_v
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__833\ : Sp12to4
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__832\ : Span12Mux_s11_h
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__831\ : Span12Mux_v
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__830\ : Odrv12
    port map (
            O => \N__5140\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__829\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5133\
        );

    \I__828\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5130\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5130\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__5127\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__824\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5118\
        );

    \I__823\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5115\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5118\,
            I => \N__5112\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__5112\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__819\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5103\
        );

    \I__818\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5100\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5100\,
            I => \U712_CHIP_RAM.REFRESH6lto2\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.REFRESH6lto2\
        );

    \I__814\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5089\,
            I => \N__5086\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__5086\,
            I => \U712_CHIP_RAM.REFRESH6lt7\
        );

    \I__811\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5079\
        );

    \I__810\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5076\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5079\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5076\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__806\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5062\
        );

    \I__805\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5062\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__802\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5051\
        );

    \I__801\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5048\
        );

    \I__800\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5045\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5048\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5045\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__796\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5031\
        );

    \I__795\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5031\
        );

    \I__794\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5028\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5023\,
            I => \N__5019\
        );

    \I__790\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__789\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5016\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5013\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__786\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5002\
        );

    \I__785\ : InMux
    port map (
            O => \N__5007\,
            I => \N__4997\
        );

    \I__784\ : InMux
    port map (
            O => \N__5006\,
            I => \N__4997\
        );

    \I__783\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4994\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5002\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4997\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4994\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__4987\,
            I => \U712_CHIP_RAM.N_54_cascade_\
        );

    \I__778\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4977\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__4980\,
            I => \N__4973\
        );

    \I__775\ : Span4Mux_h
    port map (
            O => \N__4977\,
            I => \N__4970\
        );

    \I__774\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4967\
        );

    \I__773\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4964\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4970\,
            I => \U712_CHIP_RAM.N_59\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4967\,
            I => \U712_CHIP_RAM.N_59\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4964\,
            I => \U712_CHIP_RAM.N_59\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__4957\,
            I => \U712_CHIP_RAM.N_59_cascade_\
        );

    \I__768\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__4948\,
            I => \U712_REG_SM.N_170_0\
        );

    \I__765\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4941\
        );

    \I__764\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4936\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4933\
        );

    \I__762\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4928\
        );

    \I__761\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4928\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4936\,
            I => \N__4925\
        );

    \I__759\ : Span4Mux_h
    port map (
            O => \N__4933\,
            I => \N__4922\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4928\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__4925\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__4922\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \N__4910\
        );

    \I__754\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4907\
        );

    \I__753\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4902\
        );

    \I__752\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4902\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4907\,
            I => \N__4899\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4902\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__4899\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__4894\,
            I => \N__4889\
        );

    \I__747\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4886\
        );

    \I__746\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4881\
        );

    \I__745\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4881\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4886\,
            I => \N__4878\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4881\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__4878\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__741\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4870\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_1\
        );

    \I__739\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4864\,
            I => \N__4861\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__4861\,
            I => \N__4858\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__4858\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__4855\,
            I => \N__4851\
        );

    \I__734\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4846\
        );

    \I__733\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4846\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__731\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4839\
        );

    \I__730\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4836\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4839\,
            I => \U712_REG_SM.N_169_0\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4836\,
            I => \U712_REG_SM.N_169_0\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__726\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4824\
        );

    \I__725\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4820\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4824\,
            I => \N__4817\
        );

    \I__723\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4814\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4820\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__4817\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__718\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4799\
        );

    \I__717\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4794\
        );

    \I__716\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4794\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4799\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4794\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4780\
        );

    \I__712\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4780\
        );

    \I__711\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4780\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4780\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__709\ : IoInMux
    port map (
            O => \N__4777\,
            I => \N__4773\
        );

    \I__708\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4770\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4773\,
            I => \N__4767\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4764\
        );

    \I__705\ : Span4Mux_s3_h
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__704\ : Span12Mux_h
    port map (
            O => \N__4764\,
            I => \N__4758\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__4761\,
            I => \N__4755\
        );

    \I__702\ : Span12Mux_v
    port map (
            O => \N__4758\,
            I => \N__4752\
        );

    \I__701\ : Span12Mux_v
    port map (
            O => \N__4755\,
            I => \N__4749\
        );

    \I__700\ : Odrv12
    port map (
            O => \N__4752\,
            I => \C1_c\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__4749\,
            I => \C1_c\
        );

    \I__698\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4739\
        );

    \I__697\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4736\
        );

    \I__696\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4733\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4739\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4733\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__692\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4718\
        );

    \I__691\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4715\
        );

    \I__690\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4712\
        );

    \I__689\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4707\
        );

    \I__688\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4707\
        );

    \I__687\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4704\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4712\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4707\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4704\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__4693\,
            I => \N__4688\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__4692\,
            I => \N__4685\
        );

    \I__679\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4678\
        );

    \I__678\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4675\
        );

    \I__677\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4672\
        );

    \I__676\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4665\
        );

    \I__675\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4665\
        );

    \I__674\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4665\
        );

    \I__673\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4662\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4678\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4675\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4672\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4665\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4662\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__667\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4646\
        );

    \I__666\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4641\
        );

    \I__665\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4641\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4646\,
            I => \U712_REG_SM.N_161_0\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4641\,
            I => \U712_REG_SM.N_161_0\
        );

    \I__662\ : IoInMux
    port map (
            O => \N__4636\,
            I => \N__4632\
        );

    \I__661\ : IoInMux
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4632\,
            I => \N__4626\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4623\
        );

    \I__658\ : Span4Mux_s2_v
    port map (
            O => \N__4626\,
            I => \N__4620\
        );

    \I__657\ : Span4Mux_s2_v
    port map (
            O => \N__4623\,
            I => \N__4617\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__4620\,
            I => \N__4614\
        );

    \I__655\ : Span4Mux_h
    port map (
            O => \N__4617\,
            I => \N__4611\
        );

    \I__654\ : Sp12to4
    port map (
            O => \N__4614\,
            I => \N__4608\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__4611\,
            I => \N__4605\
        );

    \I__652\ : Span12Mux_s8_v
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__651\ : Sp12to4
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__650\ : Span12Mux_h
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__649\ : Span12Mux_v
    port map (
            O => \N__4599\,
            I => \N__4593\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__4596\,
            I => \ASn_c\
        );

    \I__647\ : Odrv12
    port map (
            O => \N__4593\,
            I => \ASn_c\
        );

    \I__646\ : CEMux
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_REG_SM.N_186_0\
        );

    \I__644\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__4576\,
            I => \N__4572\
        );

    \I__641\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__4572\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4569\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__4564\,
            I => \U712_CHIP_RAM.N_58_cascade_\
        );

    \I__637\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4555\
        );

    \I__636\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4555\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\
        );

    \I__634\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4549\,
            I => \N__4546\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__4546\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_0\
        );

    \I__631\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4534\
        );

    \I__630\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4534\
        );

    \I__629\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4534\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4534\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__4531\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\
        );

    \I__626\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4524\
        );

    \I__625\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4521\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4524\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__622\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__619\ : Sp12to4
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__618\ : Span12Mux_h
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__617\ : Span12Mux_v
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__4498\,
            I => \C3_c\
        );

    \I__615\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4491\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__4494\,
            I => \N__4486\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4491\,
            I => \N__4483\
        );

    \I__612\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4478\
        );

    \I__611\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4478\
        );

    \I__610\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4475\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__4483\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4478\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4475\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__4468\,
            I => \U712_CHIP_RAM.N_67_cascade_\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__4465\,
            I => \N__4461\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__4464\,
            I => \N__4457\
        );

    \I__603\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4454\
        );

    \I__602\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4449\
        );

    \I__601\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4449\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4454\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4449\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\
        );

    \I__598\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4441\,
            I => \U712_CHIP_RAM.DBENn_7_0_0\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4438\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__4435\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4_cascade_\
        );

    \I__594\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4429\,
            I => \U712_CHIP_RAM.N_66_1\
        );

    \I__592\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4421\
        );

    \I__591\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4418\
        );

    \I__590\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4415\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4421\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4418\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4415\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__585\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4398\
        );

    \I__584\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4395\
        );

    \I__583\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4392\
        );

    \I__582\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4387\
        );

    \I__581\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4387\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4398\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4395\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4392\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4387\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__576\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4375\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4375\,
            I => \U712_REG_SM.N_181\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__4372\,
            I => \U712_REG_SM.N_170_0_cascade_\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__572\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4359\
        );

    \I__571\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4359\
        );

    \I__570\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4356\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4356\,
            I => \N__4349\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__4353\,
            I => \N__4346\
        );

    \I__566\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4343\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__4349\,
            I => \N__4340\
        );

    \I__564\ : Sp12to4
    port map (
            O => \N__4346\,
            I => \N__4333\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4333\
        );

    \I__562\ : Sp12to4
    port map (
            O => \N__4340\,
            I => \N__4333\
        );

    \I__561\ : Span12Mux_h
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__560\ : Span12Mux_v
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__4327\,
            I => \SIZ_c_1\
        );

    \I__558\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4317\
        );

    \I__557\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4317\
        );

    \I__556\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4314\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4310\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4307\
        );

    \I__553\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4304\
        );

    \I__552\ : Span4Mux_h
    port map (
            O => \N__4310\,
            I => \N__4297\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__4307\,
            I => \N__4297\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4297\
        );

    \I__549\ : Span4Mux_h
    port map (
            O => \N__4297\,
            I => \N__4294\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__4291\,
            I => \N__4288\
        );

    \I__546\ : Span4Mux_h
    port map (
            O => \N__4288\,
            I => \N__4285\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__4285\,
            I => \A_c_1\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__4282\,
            I => \N__4278\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \N__4273\
        );

    \I__542\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4268\
        );

    \I__541\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4261\
        );

    \I__540\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4261\
        );

    \I__539\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4261\
        );

    \I__538\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4256\
        );

    \I__537\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4256\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4251\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4261\,
            I => \N__4251\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N__4246\
        );

    \I__533\ : Sp12to4
    port map (
            O => \N__4251\,
            I => \N__4246\
        );

    \I__532\ : Span12Mux_v
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4243\,
            I => \A_c_0\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4240\,
            I => \N__4236\
        );

    \I__529\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4227\
        );

    \I__528\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4227\
        );

    \I__527\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4224\
        );

    \I__526\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4217\
        );

    \I__525\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4217\
        );

    \I__524\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4217\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4227\,
            I => \N__4210\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4224\,
            I => \N__4210\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4217\,
            I => \N__4210\
        );

    \I__520\ : Sp12to4
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__519\ : Span12Mux_v
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__4204\,
            I => \SIZ_c_0\
        );

    \I__517\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4198\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4198\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4195\,
            I => \U712_REG_SM.N_159_0_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4183\
        );

    \I__513\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4183\
        );

    \I__512\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4180\
        );

    \I__511\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4175\
        );

    \I__510\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4175\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4183\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4180\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4175\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__505\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4161\
        );

    \I__504\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4154\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4161\,
            I => \N__4151\
        );

    \I__502\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4146\
        );

    \I__501\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4146\
        );

    \I__500\ : InMux
    port map (
            O => \N__4158\,
            I => \N__4143\
        );

    \I__499\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4140\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4154\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__4151\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4146\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4143\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4140\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4129\,
            I => \U712_REG_SM.N_161_0_cascade_\
        );

    \I__492\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4123\,
            I => \U712_REG_SM.N_195\
        );

    \I__490\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4117\,
            I => \U712_REG_SM.N_172_0\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__4114\,
            I => \U712_REG_SM.N_195_cascade_\
        );

    \I__487\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__4105\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__4102\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__482\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4093\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__4090\,
            I => \U712_REG_SM.DS_EN_7_0\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__4087\,
            I => \U712_CHIP_RAM.N_92_cascade_\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__477\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4077\
        );

    \I__476\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4074\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4077\,
            I => \REG_TACK\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4074\,
            I => \REG_TACK\
        );

    \I__473\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4065\
        );

    \I__472\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4062\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4065\,
            I => \CPU_TACKm\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4062\,
            I => \CPU_TACKm\
        );

    \I__469\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4054\,
            I => \N__4051\
        );

    \I__467\ : Span4Mux_v
    port map (
            O => \N__4051\,
            I => \N__4047\
        );

    \I__466\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4044\
        );

    \I__465\ : Sp12to4
    port map (
            O => \N__4047\,
            I => \N__4039\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4044\,
            I => \N__4039\
        );

    \I__463\ : Span12Mux_h
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__462\ : Span12Mux_v
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__461\ : Odrv12
    port map (
            O => \N__4033\,
            I => \AWEn_c\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4030\,
            I => \N__4027\
        );

    \I__459\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__4021\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_0\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__4018\,
            I => \U712_REG_SM.N_157_0_cascade_\
        );

    \I__455\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4011\
        );

    \I__454\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4008\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4011\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4008\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__451\ : IoInMux
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4000\,
            I => \N__3997\
        );

    \I__449\ : Span12Mux_s8_v
    port map (
            O => \N__3997\,
            I => \N__3994\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__3994\,
            I => \VBENn_c\
        );

    \I__447\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3988\,
            I => \N__3984\
        );

    \I__445\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3981\
        );

    \I__444\ : Span4Mux_v
    port map (
            O => \N__3984\,
            I => \N__3978\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3981\,
            I => \N__3975\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__441\ : Span12Mux_h
    port map (
            O => \N__3975\,
            I => \N__3969\
        );

    \I__440\ : Sp12to4
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__439\ : Span12Mux_v
    port map (
            O => \N__3969\,
            I => \N__3963\
        );

    \I__438\ : Span12Mux_v
    port map (
            O => \N__3966\,
            I => \N__3960\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__3963\,
            I => \TSn_c\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__3960\,
            I => \TSn_c\
        );

    \I__435\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3952\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3952\,
            I => \N__3948\
        );

    \I__433\ : IoInMux
    port map (
            O => \N__3951\,
            I => \N__3945\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__3948\,
            I => \N__3942\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3939\
        );

    \I__430\ : Span12Mux_v
    port map (
            O => \N__3942\,
            I => \N__3936\
        );

    \I__429\ : IoSpan4Mux
    port map (
            O => \N__3939\,
            I => \N__3933\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__3936\,
            I => \RAMENn_c\
        );

    \I__427\ : Odrv4
    port map (
            O => \N__3933\,
            I => \RAMENn_c\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3928\,
            I => \U712_CHIP_RAM.N_66_1_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3925\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0_0_cascade_\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__3922\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\
        );

    \I__423\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3915\
        );

    \I__422\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3912\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3915\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3912\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__3907\,
            I => \U712_REG_SM.N_172_0_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U712_REG_SM.N_187\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3898\,
            I => \N__3894\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__3897\,
            I => \N__3891\
        );

    \I__414\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3885\
        );

    \I__413\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3880\
        );

    \I__412\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3880\
        );

    \I__411\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3875\
        );

    \I__410\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3875\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3885\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3880\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3875\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__406\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3865\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3865\,
            I => \U712_REG_SM.UDS_OUT_2_0_0\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3862\,
            I => \N__3859\
        );

    \I__403\ : InMux
    port map (
            O => \N__3859\,
            I => \N__3856\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3856\,
            I => \U712_REG_SM.LDS_OUT_2_0_0\
        );

    \I__401\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3849\
        );

    \I__400\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3846\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3849\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3846\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__397\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3837\
        );

    \I__396\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3834\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3837\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3834\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__3829\,
            I => \N__3825\
        );

    \I__392\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3822\
        );

    \I__391\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3819\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3822\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3819\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__388\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3802\
        );

    \I__387\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3802\
        );

    \I__386\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3802\
        );

    \I__385\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3802\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3802\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__382\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3789\
        );

    \I__381\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3789\
        );

    \I__380\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3786\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3789\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3786\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__377\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3775\
        );

    \I__375\ : Span4Mux_v
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__374\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3762\
        );

    \I__373\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3762\
        );

    \I__372\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3762\
        );

    \I__371\ : Span4Mux_h
    port map (
            O => \N__3769\,
            I => \N__3757\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3762\,
            I => \N__3757\
        );

    \I__369\ : Span4Mux_v
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__368\ : Sp12to4
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__367\ : Span12Mux_h
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__3748\,
            I => \CLK40_OUT_i\
        );

    \I__365\ : IoInMux
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__363\ : IoSpan4Mux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__362\ : Span4Mux_s1_h
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__361\ : Sp12to4
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__360\ : Span12Mux_v
    port map (
            O => \N__3730\,
            I => \N__3726\
        );

    \I__359\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3723\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3726\,
            I => \TACK_OUTn\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3723\,
            I => \TACK_OUTn\
        );

    \I__356\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3709\
        );

    \I__355\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3709\
        );

    \I__354\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3709\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3709\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__351\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__349\ : Span4Mux_v
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__348\ : Span4Mux_h
    port map (
            O => \N__3694\,
            I => \N__3691\
        );

    \I__347\ : Sp12to4
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3688\,
            I => \REGSPACEn_c\
        );

    \I__345\ : InMux
    port map (
            O => \N__3685\,
            I => \N__3679\
        );

    \I__344\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3679\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3679\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__342\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3664\
        );

    \I__341\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3664\
        );

    \I__340\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3664\
        );

    \I__339\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3664\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3664\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__337\ : InMux
    port map (
            O => \N__3661\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__336\ : InMux
    port map (
            O => \N__3658\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__335\ : InMux
    port map (
            O => \N__3655\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__334\ : InMux
    port map (
            O => \N__3652\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__333\ : InMux
    port map (
            O => \N__3649\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__332\ : ClkMux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__331\ : GlobalMux
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__330\ : gio2CtrlBuf
    port map (
            O => \N__3640\,
            I => \C1_c_g\
        );

    \I__329\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3634\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__327\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3627\
        );

    \I__326\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3624\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3627\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__3624\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__321\ : Span4Mux_s2_v
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__320\ : Span4Mux_v
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__319\ : Odrv4
    port map (
            O => \N__3607\,
            I => \CLK80_OUT_i_i\
        );

    \I__318\ : IoInMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__316\ : Span4Mux_s2_h
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__315\ : Span4Mux_h
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__314\ : Odrv4
    port map (
            O => \N__3592\,
            I => \CLK40_OUT_i_i\
        );

    \I__313\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3586\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3586\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__311\ : InMux
    port map (
            O => \N__3583\,
            I => \bfn_7_3_0_\
        );

    \I__310\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3577\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__308\ : InMux
    port map (
            O => \N__3574\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__307\ : InMux
    port map (
            O => \N__3571\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__306\ : IoInMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__3565\,
            I => \N__3562\
        );

    \I__304\ : IoSpan4Mux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__303\ : Span4Mux_s2_v
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__302\ : Sp12to4
    port map (
            O => \N__3556\,
            I => \N__3553\
        );

    \I__301\ : Span12Mux_v
    port map (
            O => \N__3553\,
            I => \N__3550\
        );

    \I__300\ : Odrv12
    port map (
            O => \N__3550\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7078\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4777\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9274\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3794\,
            in2 => \_gnd_net_\,
            in3 => \N__3630\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100101110"
        )
    port map (
            in0 => \N__5744\,
            in1 => \N__3904\,
            in2 => \N__4099\,
            in3 => \N__4111\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9269\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3589\,
            in2 => \_gnd_net_\,
            in3 => \N__3583\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3580\,
            in2 => \_gnd_net_\,
            in3 => \N__3574\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5106\,
            in2 => \_gnd_net_\,
            in3 => \N__3571\,
            lcout => \U712_CHIP_RAM.REFRESH6lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__3661\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5136\,
            in2 => \_gnd_net_\,
            in3 => \N__3658\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3841\,
            in2 => \_gnd_net_\,
            in3 => \N__3655\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3853\,
            in2 => \_gnd_net_\,
            in3 => \N__3652\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3828\,
            in2 => \_gnd_net_\,
            in3 => \N__3649\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3646\,
            ce => 'H',
            sr => \N__5701\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__3637\,
            in1 => \N__3811\,
            in2 => \N__6414\,
            in3 => \N__6462\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3774\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110001000"
        )
    port map (
            in0 => \N__3772\,
            in1 => \N__3814\,
            in2 => \N__6415\,
            in3 => \N__6437\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3795\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__3813\,
            in1 => \N__3729\,
            in2 => \N__3799\,
            in3 => \N__3773\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4827\,
            in1 => \N__3890\,
            in2 => \_gnd_net_\,
            in3 => \N__4842\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__3674\,
            in1 => \N__3717\,
            in2 => \N__3897\,
            in3 => \N__3919\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__3716\,
            in1 => \N__3684\,
            in2 => \N__3898\,
            in3 => \N__3675\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__3673\,
            in1 => \N__4126\,
            in2 => \N__4408\,
            in3 => \N__3718\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__3991\,
            in1 => \N__3676\,
            in2 => \N__3706\,
            in3 => \N__3685\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.C3_SYNC_2_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4164\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3918\,
            in1 => \N__4188\,
            in2 => \_gnd_net_\,
            in3 => \N__4157\,
            lcout => \U712_REG_SM.N_172_0\,
            ltout => \U712_REG_SM.N_172_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4425\,
            in2 => \N__3907\,
            in3 => \N__4404\,
            lcout => \U712_REG_SM.N_173_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4015\,
            in1 => \N__4823\,
            in2 => \N__4168\,
            in3 => \N__4189\,
            lcout => \U712_REG_SM.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__3868\,
            in1 => \N__5769\,
            in2 => \N__6867\,
            in3 => \N__3889\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9270\,
            ce => 'H',
            sr => \N__9014\
        );

    \U712_REG_SM.LDS_OUT_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001010"
        )
    port map (
            in0 => \N__3888\,
            in1 => \N__6859\,
            in2 => \N__3862\,
            in3 => \N__4575\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9270\,
            ce => 'H',
            sr => \N__9014\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4234\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNO_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4276\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100100010"
        )
    port map (
            in0 => \N__4364\,
            in1 => \N__4313\,
            in2 => \N__4281\,
            in3 => \N__4232\,
            lcout => \U712_BYTE_ENABLE.LLBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3852\,
            in1 => \N__3840\,
            in2 => \N__3829\,
            in3 => \N__5092\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9237\,
            ce => 'H',
            sr => \N__9055\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8372\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000101110"
        )
    port map (
            in0 => \N__5250\,
            in1 => \N__5532\,
            in2 => \N__4030\,
            in3 => \N__5327\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110001"
        )
    port map (
            in0 => \N__3987\,
            in1 => \N__3955\,
            in2 => \N__5609\,
            in3 => \N__8371\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__4057\,
            in1 => \N__6887\,
            in2 => \N__5533\,
            in3 => \N__5328\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__6060\,
            in1 => \N__8370\,
            in2 => \N__5680\,
            in3 => \N__4460\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__5676\,
            in1 => \N__7273\,
            in2 => \N__4464\,
            in3 => \N__6061\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0U9V_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__5894\,
            in1 => \_gnd_net_\,
            in2 => \N__6251\,
            in3 => \N__5559\,
            lcout => \U712_CHIP_RAM.N_66_1\,
            ltout => \U712_CHIP_RAM.N_66_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6051\,
            in2 => \N__3928\,
            in3 => \N__6171\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__6052\,
            in1 => \N__4984\,
            in2 => \N__3925\,
            in3 => \N__5499\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__8369\,
            in1 => \N__4069\,
            in2 => \N__3922\,
            in3 => \N__6053\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9255\,
            ce => 'H',
            sr => \N__9040\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5893\,
            in2 => \_gnd_net_\,
            in3 => \N__6231\,
            lcout => \U712_CHIP_RAM.N_92\,
            ltout => \U712_CHIP_RAM.N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__5460\,
            in1 => \N__6250\,
            in2 => \N__4087\,
            in3 => \N__4201\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9255\,
            ce => 'H',
            sr => \N__9040\
        );

    \U712_REG_SM.REG_TACK_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111000"
        )
    port map (
            in0 => \N__4893\,
            in1 => \N__4914\,
            in2 => \N__4084\,
            in3 => \N__4944\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9255\,
            ce => 'H',
            sr => \N__9040\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4080\,
            in2 => \_gnd_net_\,
            in3 => \N__4068\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__4050\,
            in1 => \N__5675\,
            in2 => \N__6871\,
            in3 => \N__5605\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4681\,
            in1 => \N__4527\,
            in2 => \N__4494\,
            in3 => \N__4721\,
            lcout => \U712_REG_SM.N_157_0\,
            ltout => \U712_REG_SM.N_157_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4160\,
            in2 => \N__4018\,
            in3 => \N__4192\,
            lcout => \U712_REG_SM.N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__5674\,
            in1 => \N__7284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4014\,
            in1 => \N__4159\,
            in2 => \_gnd_net_\,
            in3 => \N__4191\,
            lcout => \U712_REG_SM.N_159_0\,
            ltout => \U712_REG_SM.N_159_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5278\,
            in2 => \N__4195\,
            in3 => \N__5818\,
            lcout => \U712_REG_SM.N_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4190\,
            in2 => \_gnd_net_\,
            in3 => \N__4158\,
            lcout => \U712_REG_SM.N_161_0\,
            ltout => \U712_REG_SM.N_161_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4742\,
            in1 => \N__4723\,
            in2 => \N__4129\,
            in3 => \N__4683\,
            lcout => \U712_REG_SM.N_195\,
            ltout => \U712_REG_SM.N_195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__4120\,
            in1 => \N__4424\,
            in2 => \N__4114\,
            in3 => \N__4403\,
            lcout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\,
            ltout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9088\,
            in1 => \_gnd_net_\,
            in2 => \N__4102\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4528\,
            in2 => \_gnd_net_\,
            in3 => \N__4489\,
            lcout => \U712_REG_SM.N_162_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__4490\,
            in1 => \N__6844\,
            in2 => \_gnd_net_\,
            in3 => \N__4684\,
            lcout => \U712_REG_SM.DS_EN_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4722\,
            in2 => \_gnd_net_\,
            in3 => \N__4682\,
            lcout => \U712_REG_SM.N_163_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4402\,
            in1 => \N__4724\,
            in2 => \N__4692\,
            in3 => \N__4650\,
            lcout => \U712_REG_SM.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4649\,
            in1 => \N__4426\,
            in2 => \_gnd_net_\,
            in3 => \N__4401\,
            lcout => \U712_REG_SM.N_170_0\,
            ltout => \U712_REG_SM.N_170_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__4945\,
            in1 => \N__4378\,
            in2 => \N__4372\,
            in3 => \N__4743\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9268\,
            ce => 'H',
            sr => \N__9006\
        );

    \U712_BYTE_ENABLE.LMBE_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__4271\,
            in1 => \N__4323\,
            in2 => \N__4240\,
            in3 => \N__4365\,
            lcout => \U712_BYTE_ENABLE.LMBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__4324\,
            in1 => \N__4239\,
            in2 => \N__4369\,
            in3 => \N__4272\,
            lcout => \U712_BYTE_ENABLE.UUBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010110001000"
        )
    port map (
            in0 => \N__4352\,
            in1 => \N__4322\,
            in2 => \N__4282\,
            in3 => \N__4235\,
            lcout => \U712_BYTE_ENABLE.UMBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110001011100"
        )
    port map (
            in0 => \N__4444\,
            in1 => \N__6695\,
            in2 => \N__4465\,
            in3 => \N__6059\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__9051\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6035\,
            in1 => \N__6166\,
            in2 => \_gnd_net_\,
            in3 => \N__5392\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__9094\,
            in1 => \N__5007\,
            in2 => \N__5059\,
            in3 => \N__5083\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6034\,
            in1 => \N__6164\,
            in2 => \N__4980\,
            in3 => \N__5500\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_2_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5522\,
            in2 => \N__4468\,
            in3 => \N__5322\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5666\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6033\,
            in2 => \_gnd_net_\,
            in3 => \N__5910\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5459\,
            in2 => \N__4438\,
            in3 => \N__6165\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5055\,
            in2 => \N__4435\,
            in3 => \N__5006\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6152\,
            in1 => \N__4560\,
            in2 => \_gnd_net_\,
            in3 => \N__5292\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000010"
        )
    port map (
            in0 => \N__4432\,
            in1 => \N__6027\,
            in2 => \N__6172\,
            in3 => \N__4976\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000101"
        )
    port map (
            in0 => \N__6026\,
            in1 => \N__5494\,
            in2 => \N__6266\,
            in3 => \N__5246\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOMFN2_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001000000010"
        )
    port map (
            in0 => \N__4552\,
            in1 => \N__6151\,
            in2 => \N__5467\,
            in3 => \N__5175\,
            lcout => \U712_CHIP_RAM.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6028\,
            in1 => \N__5909\,
            in2 => \_gnd_net_\,
            in3 => \N__5291\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5462\,
            in1 => \N__6150\,
            in2 => \_gnd_net_\,
            in3 => \N__5381\,
            lcout => \U712_CHIP_RAM.N_58\,
            ltout => \U712_CHIP_RAM.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__6025\,
            in1 => \_gnd_net_\,
            in2 => \N__4564\,
            in3 => \N__5908\,
            lcout => \U712_CHIP_RAM.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4561\,
            in1 => \N__6153\,
            in2 => \N__5293\,
            in3 => \N__5461\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__5323\,
            in1 => \N__5851\,
            in2 => \_gnd_net_\,
            in3 => \N__4543\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9256\,
            ce => 'H',
            sr => \N__9026\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI0U9V_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__4542\,
            in1 => \N__5895\,
            in2 => \N__4855\,
            in3 => \N__6235\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4541\,
            in2 => \_gnd_net_\,
            in3 => \N__4854\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER46\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0U9V_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5896\,
            in2 => \N__4531\,
            in3 => \N__6236\,
            lcout => \U712_CHIP_RAM.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101100"
        )
    port map (
            in0 => \N__4787\,
            in1 => \N__7313\,
            in2 => \N__4807\,
            in3 => \N__4940\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__4939\,
            in1 => \N__4892\,
            in2 => \N__4915\,
            in3 => \N__4954\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000110000"
        )
    port map (
            in0 => \N__4788\,
            in1 => \N__4913\,
            in2 => \N__4894\,
            in3 => \N__4803\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4873\,
            in1 => \N__8415\,
            in2 => \N__5611\,
            in3 => \N__4867\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__4789\,
            in1 => \N__4843\,
            in2 => \N__4831\,
            in3 => \N__4802\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4691\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9265\,
            ce => 'H',
            sr => \N__9007\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4776\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9265\,
            ce => 'H',
            sr => \N__9007\
        );

    \U712_REG_SM.REGENn_1_ess_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4744\,
            in1 => \N__4725\,
            in2 => \N__4693\,
            in3 => \N__4651\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9267\,
            ce => \N__4588\,
            sr => \N__9003\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5757\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7938\,
            in1 => \N__6594\,
            in2 => \N__7066\,
            in3 => \N__5707\,
            lcout => \U712_CHIP_RAM.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5137\,
            in1 => \N__5122\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \U712_CHIP_RAM.REFRESH6lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9091\,
            in1 => \N__5082\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__9093\,
            in2 => \N__5071\,
            in3 => \N__5022\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__5067\,
            in2 => \_gnd_net_\,
            in3 => \N__5037\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5054\,
            in1 => \N__5036\,
            in2 => \N__5023\,
            in3 => \N__5005\,
            lcout => \U712_CHIP_RAM.N_54\,
            ltout => \U712_CHIP_RAM.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4987\,
            in3 => \N__5453\,
            lcout => \U712_CHIP_RAM.N_59\,
            ltout => \U712_CHIP_RAM.N_59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__6023\,
            in1 => \N__6162\,
            in2 => \N__4957\,
            in3 => \N__5904\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISSMN4_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7153\,
            in1 => \N__5563\,
            in2 => \N__5263\,
            in3 => \N__6274\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__5260\,
            in1 => \N__6024\,
            in2 => \N__5254\,
            in3 => \N__5211\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9036\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL41I5_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__6195\,
            in1 => \N__6092\,
            in2 => \_gnd_net_\,
            in3 => \N__5495\,
            lcout => \U712_CHIP_RAM.N_74\,
            ltout => \U712_CHIP_RAM.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6031\,
            in2 => \N__5200\,
            in3 => \N__5197\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL41I5_0_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__7151\,
            in2 => \N__5394\,
            in3 => \N__5410\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4U4DE_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__6100\,
            in1 => \N__5349\,
            in2 => \N__5191\,
            in3 => \N__5188\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE2282_3_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__7150\,
            in2 => \N__5182\,
            in3 => \N__6154\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a3_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5385\,
            in2 => \N__5161\,
            in3 => \N__6029\,
            lcout => \U712_CHIP_RAM.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIV8F93_3_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5455\,
            in1 => \N__7152\,
            in2 => \N__5393\,
            in3 => \N__6155\,
            lcout => \U712_CHIP_RAM.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010100"
        )
    port map (
            in0 => \N__5356\,
            in1 => \N__5350\,
            in2 => \N__5332\,
            in3 => \N__6032\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9245\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3EN62_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__6269\,
            in2 => \_gnd_net_\,
            in3 => \N__5569\,
            lcout => \U712_CHIP_RAM.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27CG_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5556\,
            in2 => \_gnd_net_\,
            in3 => \N__6267\,
            lcout => \U712_CHIP_RAM.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_SYNC_RNI17BM1_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5817\,
            in1 => \N__5274\,
            in2 => \N__5673\,
            in3 => \N__5610\,
            lcout => \U712_CHIP_RAM.N_55\,
            ltout => \U712_CHIP_RAM.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3EN62_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5558\,
            in1 => \_gnd_net_\,
            in2 => \N__5536\,
            in3 => \N__6268\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIN5LK4_3_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6163\,
            in1 => \N__5493\,
            in2 => \N__5466\,
            in3 => \N__5409\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKJ6F7_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__9087\,
            in1 => \N__6037\,
            in2 => \N__5398\,
            in3 => \N__5395\,
            lcout => \U712_CHIP_RAM.N_61\,
            ltout => \U712_CHIP_RAM.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRDCDD_0_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5348\,
            in2 => \N__5335\,
            in3 => \N__5321\,
            lcout => \U712_CHIP_RAM.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5816\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9257\,
            ce => 'H',
            sr => \N__9008\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9257\,
            ce => 'H',
            sr => \N__9008\
        );

    \TACKn_obuft_RNO_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_517_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5758\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REF_SYNC_1_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7939\,
            lcout => \U712_CHIP_RAM.REF_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9228\,
            ce => 'H',
            sr => \N__9041\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7065\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9228\,
            ce => 'H',
            sr => \N__9041\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8113\,
            in1 => \N__8222\,
            in2 => \N__8792\,
            in3 => \N__8641\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__7285\,
            in1 => \N__5689\,
            in2 => \_gnd_net_\,
            in3 => \N__5656\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9235\,
            ce => 'H',
            sr => \N__9027\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6196\,
            in2 => \_gnd_net_\,
            in3 => \N__6094\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__6492\,
            in1 => \N__6078\,
            in2 => \N__5614\,
            in3 => \N__8221\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__6020\,
            in1 => \N__5911\,
            in2 => \_gnd_net_\,
            in3 => \N__6270\,
            lcout => \U712_CHIP_RAM.N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6076\,
            in2 => \_gnd_net_\,
            in3 => \N__8135\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__6079\,
            in1 => \N__6493\,
            in2 => \N__8648\,
            in3 => \N__6178\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7156\,
            in1 => \N__6021\,
            in2 => \N__5919\,
            in3 => \N__6170\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6022\,
            in1 => \N__6093\,
            in2 => \N__5938\,
            in3 => \N__5915\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__6478\,
            in1 => \N__6077\,
            in2 => \N__6064\,
            in3 => \N__8757\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6713\,
            in2 => \_gnd_net_\,
            in3 => \N__7297\,
            lcout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__5950\,
            in2 => \N__5937\,
            in3 => \N__5920\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7154\,
            in2 => \N__5842\,
            in3 => \N__6491\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7155\,
            in1 => \N__6403\,
            in2 => \N__6469\,
            in3 => \N__6444\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9086\,
            in1 => \_gnd_net_\,
            in2 => \N__6448\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__6445\,
            in1 => \N__7141\,
            in2 => \_gnd_net_\,
            in3 => \N__6413\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9251\,
            ce => \N__6367\,
            sr => \N__9004\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__6961\,
            in1 => \N__7228\,
            in2 => \N__8449\,
            in3 => \N__6355\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6640\,
            in1 => \N__8247\,
            in2 => \_gnd_net_\,
            in3 => \N__8140\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9227\,
            ce => \N__8023\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6547\,
            in1 => \N__8248\,
            in2 => \_gnd_net_\,
            in3 => \N__8141\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9227\,
            ce => \N__8023\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7393\,
            in1 => \N__8454\,
            in2 => \N__8811\,
            in3 => \N__7858\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8455\,
            in1 => \N__6679\,
            in2 => \N__6664\,
            in3 => \N__6661\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__6634\,
            in1 => \N__8459\,
            in2 => \N__6619\,
            in3 => \N__6541\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__7055\,
            in1 => \N__9089\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => \U712_CHIP_RAM.N_50_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__6583\,
            in1 => \N__6568\,
            in2 => \N__8461\,
            in3 => \N__7447\,
            lcout => \U712_CHIP_RAM.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6535\,
            in1 => \N__8379\,
            in2 => \N__8816\,
            in3 => \N__7627\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7618\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9230\,
            ce => \N__7505\,
            sr => \N__9013\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__7663\,
            in1 => \N__8733\,
            in2 => \N__8447\,
            in3 => \N__7708\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8423\,
            in1 => \N__6529\,
            in2 => \N__6511\,
            in3 => \N__6508\,
            lcout => \U712_CHIP_RAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__8732\,
            in1 => \N__8200\,
            in2 => \N__8114\,
            in3 => \N__8631\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8420\,
            in1 => \N__7669\,
            in2 => \N__8810\,
            in3 => \N__7744\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__6997\,
            in1 => \N__6982\,
            in2 => \N__6964\,
            in3 => \N__8421\,
            lcout => \U712_CHIP_RAM.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110001"
        )
    port map (
            in0 => \N__8422\,
            in1 => \N__6957\,
            in2 => \N__6946\,
            in3 => \N__8901\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_i_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__6900\,
            in1 => \N__6866\,
            in2 => \N__7338\,
            in3 => \N__7298\,
            lcout => \DRDDIR_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8777\,
            in1 => \N__7516\,
            in2 => \N__8448\,
            in3 => \N__7657\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__6781\,
            in2 => \N__6766\,
            in3 => \N__6763\,
            lcout => \U712_CHIP_RAM.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__6745\,
            in1 => \N__8263\,
            in2 => \N__8809\,
            in3 => \N__8139\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9243\,
            ce => \N__8021\,
            sr => \N__9001\
        );

    \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6720\,
            in2 => \_gnd_net_\,
            in3 => \N__7300\,
            lcout => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\,
            ltout => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__7227\,
            in1 => \N__8431\,
            in2 => \N__6682\,
            in3 => \N__7372\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7299\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__7162\,
            in2 => \_gnd_net_\,
            in3 => \N__7173\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8894\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7214\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9260\,
            ce => 'H',
            sr => \N__8997\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7174\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9260\,
            ce => 'H',
            sr => \N__8997\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7108\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7963\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9229\,
            ce => 'H',
            sr => \N__9042\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8146\,
            in1 => \N__7042\,
            in2 => \_gnd_net_\,
            in3 => \N__8260\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__8018\,
            sr => \N__9037\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8259\,
            in1 => \N__8813\,
            in2 => \N__8158\,
            in3 => \N__8650\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__8018\,
            sr => \N__9037\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000101"
        )
    port map (
            in0 => \N__8812\,
            in1 => \N__7399\,
            in2 => \N__8157\,
            in3 => \N__8261\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__8018\,
            sr => \N__9037\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9090\,
            in2 => \_gnd_net_\,
            in3 => \N__7453\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7384\,
            in1 => \N__8376\,
            in2 => \N__8814\,
            in3 => \N__7783\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8793\,
            in1 => \N__7378\,
            in2 => \N__8416\,
            in3 => \N__7591\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7675\,
            in1 => \N__8377\,
            in2 => \N__8815\,
            in3 => \N__7822\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8378\,
            in1 => \N__7441\,
            in2 => \N__7423\,
            in3 => \N__7420\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7845\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9319\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7651\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7815\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => \N__7510\,
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7555\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9246\,
            ce => \N__9127\,
            sr => \N__9009\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7650\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9246\,
            ce => \N__9127\,
            sr => \N__9009\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7614\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9246\,
            ce => \N__9127\,
            sr => \N__9009\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7582\,
            in1 => \N__8262\,
            in2 => \_gnd_net_\,
            in3 => \N__8153\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9252\,
            ce => \N__8022\,
            sr => \N__9005\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7554\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9258\,
            ce => \N__7506\,
            sr => \N__9002\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7773\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9258\,
            ce => \N__7506\,
            sr => \N__9002\
        );

    \U712_CHIP_RAM.REF_SYNC_0_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7959\,
            in2 => \_gnd_net_\,
            in3 => \N__8523\,
            lcout => \U712_CHIP_RAM.REF_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9232\,
            ce => 'H',
            sr => \N__9052\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__8249\,
            in2 => \_gnd_net_\,
            in3 => \N__8142\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__7924\,
            in1 => \N__7918\,
            in2 => \N__8460\,
            in3 => \N__7903\,
            lcout => \U712_CHIP_RAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7887\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9242\,
            ce => \N__9134\,
            sr => \N__9038\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9242\,
            ce => \N__9134\,
            sr => \N__9038\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7816\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9242\,
            ce => \N__9134\,
            sr => \N__9038\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7777\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9247\,
            ce => \N__9139\,
            sr => \N__9028\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7728\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9247\,
            ce => \N__9139\,
            sr => \N__9028\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__7699\,
            in1 => \N__7684\,
            in2 => \N__8902\,
            in3 => \N__8450\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8156\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9233\,
            ce => 'H',
            sr => \N__9056\
        );

    \U712_CHIP_RAM.CASn_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8818\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9233\,
            ce => 'H',
            sr => \N__9056\
        );

    \U712_CHIP_RAM.RASn_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8266\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9236\,
            ce => 'H',
            sr => \N__9054\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9236\,
            ce => 'H',
            sr => \N__9054\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__8590\,
            in1 => \N__8264\,
            in2 => \_gnd_net_\,
            in3 => \N__8155\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => \N__8019\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__8563\,
            in1 => \N__8490\,
            in2 => \N__9286\,
            in3 => \N__8380\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => \N__8019\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__8516\,
            in1 => \N__8491\,
            in2 => \N__8482\,
            in3 => \N__8381\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => \N__8019\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8265\,
            in1 => \N__8167\,
            in2 => \_gnd_net_\,
            in3 => \N__8154\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9253\,
            ce => \N__8020\,
            sr => \N__9039\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9259\,
            ce => \N__9135\,
            sr => \N__9029\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 21 2024 14:06:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    A : in std_logic_vector(31 downto 1);
    RnW : in std_logic;
    CIACS1n : out std_logic;
    TT1 : in std_logic;
    TICK50 : out std_logic;
    RAMSPACEn : out std_logic;
    TT0 : in std_logic;
    TICK60 : out std_logic;
    LBENn : in std_logic;
    CLKCIA : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    BUFENn : out std_logic;
    TSn : in std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2373\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_CIA.g0Z0Z_11\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_CIA.g0Z0Z_8\ : std_logic;
signal \A_c_21\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_30\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U409_CIA.g0Z0Z_2\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_CIA.g0Z0Z_10_cascade_\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un10_ROMENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un6_ROMENZ0\ : std_logic;
signal \OVL_c\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.RESETn_c_i\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ROMEN_0\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_97\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \U409_TICK.TICK603_11_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_353_i\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4692\,
            RESETB => \N__4977\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6077\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6079\,
            DIN => \N__6078\,
            DOUT => \N__6077\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6079\,
            PADOUT => \N__6078\,
            PADIN => \N__6077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6067\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6069\,
            DIN => \N__6068\,
            DOUT => \N__6067\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6069\,
            PADOUT => \N__6068\,
            PADIN => \N__6067\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6058\,
            DIN => \N__6057\,
            DOUT => \N__6056\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6058\,
            PADOUT => \N__6057\,
            PADIN => \N__6056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4275\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6049\,
            DIN => \N__6048\,
            DOUT => \N__6047\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6049\,
            PADOUT => \N__6048\,
            PADIN => \N__6047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6040\,
            DIN => \N__6039\,
            DOUT => \N__6038\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6040\,
            PADOUT => \N__6039\,
            PADIN => \N__6038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6031\,
            DIN => \N__6030\,
            DOUT => \N__6029\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6031\,
            PADOUT => \N__6030\,
            PADIN => \N__6029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6022\,
            DIN => \N__6021\,
            DOUT => \N__6020\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6022\,
            PADOUT => \N__6021\,
            PADIN => \N__6020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2916\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6013\,
            DIN => \N__6012\,
            DOUT => \N__6011\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6013\,
            PADOUT => \N__6012\,
            PADIN => \N__6011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3072\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6004\,
            DIN => \N__6003\,
            DOUT => \N__6002\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6004\,
            PADOUT => \N__6003\,
            PADIN => \N__6002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5995\,
            DIN => \N__5994\,
            DOUT => \N__5993\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5995\,
            PADOUT => \N__5994\,
            PADIN => \N__5993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5986\,
            DIN => \N__5985\,
            DOUT => \N__5984\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5986\,
            PADOUT => \N__5985\,
            PADIN => \N__5984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3048\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5977\,
            DIN => \N__5976\,
            DOUT => \N__5975\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__5977\,
            PADOUT => \N__5976\,
            PADIN => \N__5975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5610\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__3597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5968\,
            DIN => \N__5967\,
            DOUT => \N__5966\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5968\,
            PADOUT => \N__5967\,
            PADIN => \N__5966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5959\,
            DIN => \N__5958\,
            DOUT => \N__5957\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5959\,
            PADOUT => \N__5958\,
            PADIN => \N__5957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5950\,
            DIN => \N__5949\,
            DOUT => \N__5948\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5950\,
            PADOUT => \N__5949\,
            PADIN => \N__5948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5941\,
            DIN => \N__5940\,
            DOUT => \N__5939\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5941\,
            PADOUT => \N__5940\,
            PADIN => \N__5939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5586\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5932\,
            DIN => \N__5931\,
            DOUT => \N__5930\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5932\,
            PADOUT => \N__5931\,
            PADIN => \N__5930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3162\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5923\,
            DIN => \N__5922\,
            DOUT => \N__5921\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5923\,
            PADOUT => \N__5922\,
            PADIN => \N__5921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5914\,
            DIN => \N__5913\,
            DOUT => \N__5912\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5914\,
            PADOUT => \N__5913\,
            PADIN => \N__5912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5905\,
            DIN => \N__5904\,
            DOUT => \N__5903\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5905\,
            PADOUT => \N__5904\,
            PADIN => \N__5903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5896\,
            DIN => \N__5895\,
            DOUT => \N__5894\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5896\,
            PADOUT => \N__5895\,
            PADIN => \N__5894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5887\,
            DIN => \N__5886\,
            DOUT => \N__5885\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5887\,
            PADOUT => \N__5886\,
            PADIN => \N__5885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5878\,
            DIN => \N__5877\,
            DOUT => \N__5876\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5878\,
            PADOUT => \N__5877\,
            PADIN => \N__5876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5869\,
            DIN => \N__5868\,
            DOUT => \N__5867\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5869\,
            PADOUT => \N__5868\,
            PADIN => \N__5867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5860\,
            DIN => \N__5859\,
            DOUT => \N__5858\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5860\,
            PADOUT => \N__5859\,
            PADIN => \N__5858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5851\,
            DIN => \N__5850\,
            DOUT => \N__5849\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5851\,
            PADOUT => \N__5850\,
            PADIN => \N__5849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5842\,
            DIN => \N__5841\,
            DOUT => \N__5840\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5842\,
            PADOUT => \N__5841\,
            PADIN => \N__5840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2880\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5833\,
            DIN => \N__5832\,
            DOUT => \N__5831\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5833\,
            PADOUT => \N__5832\,
            PADIN => \N__5831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4350\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5824\,
            DIN => \N__5823\,
            DOUT => \N__5822\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5824\,
            PADOUT => \N__5823\,
            PADIN => \N__5822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5815\,
            DIN => \N__5814\,
            DOUT => \N__5813\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5815\,
            PADOUT => \N__5814\,
            PADIN => \N__5813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5806\,
            DIN => \N__5805\,
            DOUT => \N__5804\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5806\,
            PADOUT => \N__5805\,
            PADIN => \N__5804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5797\,
            DIN => \N__5796\,
            DOUT => \N__5795\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5797\,
            PADOUT => \N__5796\,
            PADIN => \N__5795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5788\,
            DIN => \N__5787\,
            DOUT => \N__5786\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5788\,
            PADOUT => \N__5787\,
            PADIN => \N__5786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5779\,
            DIN => \N__5778\,
            DOUT => \N__5777\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5779\,
            PADOUT => \N__5778\,
            PADIN => \N__5777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4209\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__5770\,
            DIN => \N__5769\,
            DOUT => \N__5768\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5770\,
            PADOUT => \N__5769\,
            PADIN => \N__5768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__5751\,
            I => \N__5746\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5740\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5740\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5737\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5734\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__5740\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5734\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5724\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5718\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__5715\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__5712\,
            I => \N__5702\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5699\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5696\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5689\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5689\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5689\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5682\
        );

    \I__1313\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5682\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5682\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5699\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5696\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5689\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5682\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5664\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5657\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5657\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5657\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5650\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5650\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5650\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5664\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5657\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__5650\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1297\ : ClkMux
    port map (
            O => \N__5643\,
            I => \N__5631\
        );

    \I__1296\ : ClkMux
    port map (
            O => \N__5642\,
            I => \N__5631\
        );

    \I__1295\ : ClkMux
    port map (
            O => \N__5641\,
            I => \N__5631\
        );

    \I__1294\ : ClkMux
    port map (
            O => \N__5640\,
            I => \N__5631\
        );

    \I__1293\ : GlobalMux
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__1292\ : gio2CtrlBuf
    port map (
            O => \N__5628\,
            I => \CLK28_IN_c_g\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5622\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__5619\,
            I => \N__5616\
        );

    \I__1288\ : Sp12to4
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__5613\,
            I => \TACK_EN_i\
        );

    \I__1286\ : IoInMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__1284\ : IoSpan4Mux
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__1283\ : Span4Mux_s1_v
    port map (
            O => \N__5601\,
            I => \N__5598\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__5598\,
            I => \N__5595\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__5595\,
            I => \N__5592\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__5589\,
            I => \N_353_i\
        );

    \I__1278\ : IoInMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5580\
        );

    \I__1276\ : Span4Mux_s1_v
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__1275\ : Sp12to4
    port map (
            O => \N__5577\,
            I => \N__5573\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5570\
        );

    \I__1273\ : Span12Mux_h
    port map (
            O => \N__5573\,
            I => \N__5567\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5564\
        );

    \I__1271\ : Span12Mux_v
    port map (
            O => \N__5567\,
            I => \N__5559\
        );

    \I__1270\ : Span12Mux_h
    port map (
            O => \N__5564\,
            I => \N__5559\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__5559\,
            I => \BUFENn_c\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1266\ : Span12Mux_h
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1265\ : Span12Mux_v
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__1264\ : Odrv12
    port map (
            O => \N__5544\,
            I => \TACKn_in\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5538\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5534\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5530\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__5534\,
            I => \N__5526\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \N__5517\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5508\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5505\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__5526\,
            I => \N__5501\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5492\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5492\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5492\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5492\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5489\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5486\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5479\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5479\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5479\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5476\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5469\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5469\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5469\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__5508\,
            I => \N__5463\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5505\,
            I => \N__5463\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5460\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__5501\,
            I => \N__5444\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5492\,
            I => \N__5444\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5489\,
            I => \N__5444\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5486\,
            I => \N__5444\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5444\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5476\,
            I => \N__5444\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5469\,
            I => \N__5444\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5441\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5463\,
            I => \N__5436\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5460\,
            I => \N__5436\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5432\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__5444\,
            I => \N__5429\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__5441\,
            I => \N__5426\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__5436\,
            I => \N__5423\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5420\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5432\,
            I => \N__5417\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__5429\,
            I => \N__5414\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5411\
        );

    \I__1221\ : Span4Mux_h
    port map (
            O => \N__5423\,
            I => \N__5408\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5405\
        );

    \I__1219\ : Span4Mux_h
    port map (
            O => \N__5417\,
            I => \N__5402\
        );

    \I__1218\ : Sp12to4
    port map (
            O => \N__5414\,
            I => \N__5397\
        );

    \I__1217\ : Sp12to4
    port map (
            O => \N__5411\,
            I => \N__5397\
        );

    \I__1216\ : Sp12to4
    port map (
            O => \N__5408\,
            I => \N__5392\
        );

    \I__1215\ : Span12Mux_h
    port map (
            O => \N__5405\,
            I => \N__5392\
        );

    \I__1214\ : Span4Mux_h
    port map (
            O => \N__5402\,
            I => \N__5389\
        );

    \I__1213\ : Span12Mux_h
    port map (
            O => \N__5397\,
            I => \N__5386\
        );

    \I__1212\ : Span12Mux_v
    port map (
            O => \N__5392\,
            I => \N__5383\
        );

    \I__1211\ : Sp12to4
    port map (
            O => \N__5389\,
            I => \N__5380\
        );

    \I__1210\ : Span12Mux_v
    port map (
            O => \N__5386\,
            I => \N__5375\
        );

    \I__1209\ : Span12Mux_h
    port map (
            O => \N__5383\,
            I => \N__5375\
        );

    \I__1208\ : Span12Mux_v
    port map (
            O => \N__5380\,
            I => \N__5372\
        );

    \I__1207\ : Odrv12
    port map (
            O => \N__5375\,
            I => \RESETn_c\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__5372\,
            I => \RESETn_c\
        );

    \I__1205\ : SRMux
    port map (
            O => \N__5367\,
            I => \N__5362\
        );

    \I__1204\ : SRMux
    port map (
            O => \N__5366\,
            I => \N__5359\
        );

    \I__1203\ : SRMux
    port map (
            O => \N__5365\,
            I => \N__5356\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5362\,
            I => \N__5353\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5350\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5347\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__5353\,
            I => \N__5344\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__5350\,
            I => \N__5341\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__5347\,
            I => \N__5338\
        );

    \I__1196\ : Sp12to4
    port map (
            O => \N__5344\,
            I => \N__5335\
        );

    \I__1195\ : Span4Mux_h
    port map (
            O => \N__5341\,
            I => \N__5332\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__5338\,
            I => \N__5329\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__5335\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5332\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__5329\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5322\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5315\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5312\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5315\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5312\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1185\ : ClkMux
    port map (
            O => \N__5307\,
            I => \N__5280\
        );

    \I__1184\ : ClkMux
    port map (
            O => \N__5306\,
            I => \N__5280\
        );

    \I__1183\ : ClkMux
    port map (
            O => \N__5305\,
            I => \N__5280\
        );

    \I__1182\ : ClkMux
    port map (
            O => \N__5304\,
            I => \N__5280\
        );

    \I__1181\ : ClkMux
    port map (
            O => \N__5303\,
            I => \N__5280\
        );

    \I__1180\ : ClkMux
    port map (
            O => \N__5302\,
            I => \N__5280\
        );

    \I__1179\ : ClkMux
    port map (
            O => \N__5301\,
            I => \N__5280\
        );

    \I__1178\ : ClkMux
    port map (
            O => \N__5300\,
            I => \N__5280\
        );

    \I__1177\ : ClkMux
    port map (
            O => \N__5299\,
            I => \N__5280\
        );

    \I__1176\ : GlobalMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__1175\ : gio2CtrlBuf
    port map (
            O => \N__5277\,
            I => \CLK6_c_g\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5274\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5271\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5268\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5265\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5262\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5251\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5251\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5246\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5246\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5251\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5246\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5227\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5227\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5227\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5227\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5222\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5222\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5227\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5222\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5217\,
            I => \N__5213\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5208\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5203\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5203\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5200\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5203\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5200\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5186\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5183\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__5186\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5183\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5178\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5171\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5168\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5171\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5168\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5157\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5154\,
            I => \bfn_12_7_0_\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5147\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5144\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5147\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5144\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5139\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__5136\,
            I => \N__5133\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5129\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5126\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5112\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5105\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5102\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5097\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5090\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5087\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5090\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5087\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5079\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5076\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5069\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5066\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5066\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5058\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5055\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5048\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5045\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5048\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5045\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__5031\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5028\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5014\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5014\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5014\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5009\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5009\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5009\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4995\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4990\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4990\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4987\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4984\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4990\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4987\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__4984\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__1073\ : Span4Mux_s2_v
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__4965\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__4962\,
            I => \N__4958\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4952\
        );

    \I__1068\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4952\
        );

    \I__1067\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4949\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__4944\,
            I => \N__4938\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4935\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4930\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4930\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4927\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__4935\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__4930\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__4927\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4916\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4913\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4916\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__4913\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4908\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4901\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4898\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4901\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4898\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4893\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__1043\ : Span4Mux_h
    port map (
            O => \N__4881\,
            I => \N__4877\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4874\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__4877\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__4874\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4869\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4862\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4859\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4848\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4841\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4838\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4841\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4838\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4830\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4827\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4820\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4820\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4812\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4803\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4803\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4803\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__4800\,
            I => \N__4791\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4788\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4785\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4782\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4773\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4773\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4773\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4773\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4788\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4785\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4782\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4764\,
            I => \N__4757\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4754\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4747\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4747\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4747\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__996\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4735\
        );

    \I__995\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4730\
        );

    \I__994\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4730\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4730\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \N__4722\
        );

    \I__990\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4719\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__4716\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\
        );

    \I__987\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4705\
        );

    \I__986\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4705\
        );

    \I__985\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4702\
        );

    \I__984\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4699\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4705\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4702\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4699\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__980\ : IoInMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4684\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__4688\,
            I => \N__4680\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4687\,
            I => \N__4676\
        );

    \I__976\ : Span4Mux_s2_v
    port map (
            O => \N__4684\,
            I => \N__4673\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4683\,
            I => \N__4670\
        );

    \I__974\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4667\
        );

    \I__973\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4662\
        );

    \I__972\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4662\
        );

    \I__971\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4659\
        );

    \I__970\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4656\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4653\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4649\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__4659\,
            I => \N__4644\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4644\
        );

    \I__965\ : Span4Mux_v
    port map (
            O => \N__4653\,
            I => \N__4641\
        );

    \I__964\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4638\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__4649\,
            I => \N__4633\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__4644\,
            I => \N__4633\
        );

    \I__961\ : Sp12to4
    port map (
            O => \N__4641\,
            I => \N__4630\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4627\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__4633\,
            I => \N__4624\
        );

    \I__958\ : Span12Mux_h
    port map (
            O => \N__4630\,
            I => \N__4621\
        );

    \I__957\ : Sp12to4
    port map (
            O => \N__4627\,
            I => \N__4618\
        );

    \I__956\ : Span12Mux_h
    port map (
            O => \N__4624\,
            I => \N__4615\
        );

    \I__955\ : Span12Mux_v
    port map (
            O => \N__4621\,
            I => \N__4612\
        );

    \I__954\ : Span12Mux_v
    port map (
            O => \N__4618\,
            I => \N__4609\
        );

    \I__953\ : Span12Mux_v
    port map (
            O => \N__4615\,
            I => \N__4606\
        );

    \I__952\ : Odrv12
    port map (
            O => \N__4612\,
            I => \CLK40_IN_c\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__4609\,
            I => \CLK40_IN_c\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__4606\,
            I => \CLK40_IN_c\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4599\,
            I => \N__4594\
        );

    \I__948\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4591\
        );

    \I__947\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4588\
        );

    \I__946\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4585\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4591\,
            I => \N__4580\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4588\,
            I => \N__4580\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4585\,
            I => \N__4577\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__941\ : Span4Mux_v
    port map (
            O => \N__4577\,
            I => \N__4571\
        );

    \I__940\ : Sp12to4
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__939\ : Span4Mux_h
    port map (
            O => \N__4571\,
            I => \N__4565\
        );

    \I__938\ : Span12Mux_h
    port map (
            O => \N__4568\,
            I => \N__4560\
        );

    \I__937\ : Sp12to4
    port map (
            O => \N__4565\,
            I => \N__4560\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__4557\,
            I => \TSn_c\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__4554\,
            I => \N__4550\
        );

    \I__933\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4547\
        );

    \I__932\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4544\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__929\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4532\
        );

    \I__928\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4532\
        );

    \I__927\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4529\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4532\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4529\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4524\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__923\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\
        );

    \I__921\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4509\
        );

    \I__920\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4506\
        );

    \I__919\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4501\
        );

    \I__918\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4501\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4509\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4506\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4501\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__914\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4485\
        );

    \I__913\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4485\
        );

    \I__912\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4485\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4485\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__4482\,
            I => \N__4477\
        );

    \I__909\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4472\
        );

    \I__908\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4463\
        );

    \I__907\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4463\
        );

    \I__906\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4463\
        );

    \I__905\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4463\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4463\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__901\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4443\
        );

    \I__900\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4443\
        );

    \I__899\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4436\
        );

    \I__898\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4436\
        );

    \I__897\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4436\
        );

    \I__896\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4429\
        );

    \I__895\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4429\
        );

    \I__894\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4429\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4443\,
            I => \U409_TICK.TICK503_14\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4436\,
            I => \U409_TICK.TICK503_14\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4429\,
            I => \U409_TICK.TICK503_14\
        );

    \I__890\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4410\
        );

    \I__889\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4410\
        );

    \I__888\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4403\
        );

    \I__887\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4403\
        );

    \I__886\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4403\
        );

    \I__885\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4396\
        );

    \I__884\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4396\
        );

    \I__883\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4396\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4410\,
            I => \U409_TICK.TICK503_10\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4403\,
            I => \U409_TICK.TICK503_10\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4396\,
            I => \U409_TICK.TICK503_10\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4389\,
            I => \N__4384\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__4388\,
            I => \N__4379\
        );

    \I__877\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4371\
        );

    \I__876\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4371\
        );

    \I__875\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4364\
        );

    \I__874\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4364\
        );

    \I__873\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4364\
        );

    \I__872\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4357\
        );

    \I__871\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4357\
        );

    \I__870\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4357\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4371\,
            I => \U409_TICK.TICK503_9\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U409_TICK.TICK503_9\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4357\,
            I => \U409_TICK.TICK503_9\
        );

    \I__866\ : IoInMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__864\ : Span4Mux_s1_v
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__862\ : Span12Mux_h
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__861\ : Span12Mux_v
    port map (
            O => \N__4335\,
            I => \N__4331\
        );

    \I__860\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4328\
        );

    \I__859\ : Odrv12
    port map (
            O => \N__4331\,
            I => \TICK50_c\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4328\,
            I => \TICK50_c\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4323\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__855\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4313\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__4316\,
            I => \N__4309\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4313\,
            I => \N__4305\
        );

    \I__852\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4300\
        );

    \I__851\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4300\
        );

    \I__850\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4297\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4305\,
            I => \N__4292\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4300\,
            I => \N__4292\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4297\,
            I => \U409_CIA.VMAZ0\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4292\,
            I => \U409_CIA.VMAZ0\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4287\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__844\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4281\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__4278\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__841\ : IoInMux
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__839\ : Span4Mux_s1_v
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__837\ : Sp12to4
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__836\ : Span12Mux_h
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__835\ : Span12Mux_v
    port map (
            O => \N__4257\,
            I => \N__4252\
        );

    \I__834\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4249\
        );

    \I__833\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4246\
        );

    \I__832\ : Odrv12
    port map (
            O => \N__4252\,
            I => \CLKCIA_c\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4249\,
            I => \CLKCIA_c\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4246\,
            I => \CLKCIA_c\
        );

    \I__829\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4235\
        );

    \I__828\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4232\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4235\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4232\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__825\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4224\,
            I => \U409_TICK.TICK503_11\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__4221\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4212\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__819\ : IoInMux
    port map (
            O => \N__4209\,
            I => \N__4206\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__817\ : Span4Mux_s2_v
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__815\ : Span4Mux_v
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__814\ : Span4Mux_h
    port map (
            O => \N__4194\,
            I => \N__4190\
        );

    \I__813\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4187\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__4190\,
            I => \TICK60_c\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4187\,
            I => \TICK60_c\
        );

    \I__810\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4179\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__807\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__805\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4163\
        );

    \I__804\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4160\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4160\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__801\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4151\
        );

    \I__800\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4148\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4151\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4148\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__797\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4139\
        );

    \I__796\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4136\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4139\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4136\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__792\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4125\,
            I => \N__4121\
        );

    \I__790\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4121\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4118\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__787\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__786\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4109\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4106\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__4101\,
            I => \N__4096\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__4100\,
            I => \N__4092\
        );

    \I__781\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4084\
        );

    \I__780\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4084\
        );

    \I__779\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4079\
        );

    \I__778\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4079\
        );

    \I__777\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4072\
        );

    \I__776\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4072\
        );

    \I__775\ : InMux
    port map (
            O => \N__4089\,
            I => \N__4072\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4084\,
            I => \U409_TICK.TICK603_10\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4079\,
            I => \U409_TICK.TICK603_10\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4072\,
            I => \U409_TICK.TICK603_10\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__4065\,
            I => \N__4059\
        );

    \I__770\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4050\
        );

    \I__769\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4050\
        );

    \I__768\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4043\
        );

    \I__767\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4043\
        );

    \I__766\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4043\
        );

    \I__765\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4036\
        );

    \I__764\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4036\
        );

    \I__763\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4036\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4050\,
            I => \U409_TICK.TICK603_9\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4043\,
            I => \U409_TICK.TICK603_9\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4036\,
            I => \U409_TICK.TICK603_9\
        );

    \I__759\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4019\
        );

    \I__758\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4019\
        );

    \I__757\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4019\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__4026\,
            I => \N__4016\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4010\
        );

    \I__754\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4007\
        );

    \I__753\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4004\
        );

    \I__752\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4001\
        );

    \I__751\ : InMux
    port map (
            O => \N__4013\,
            I => \N__3998\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__4010\,
            I => \N__3995\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4007\,
            I => \U409_TICK.TICK603_14\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U409_TICK.TICK603_14\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4001\,
            I => \U409_TICK.TICK603_14\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3998\,
            I => \U409_TICK.TICK603_14\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__3995\,
            I => \U409_TICK.TICK603_14\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__3984\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3978\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__3975\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__3972\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__3969\,
            I => \N__3964\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__3968\,
            I => \N__3961\
        );

    \I__737\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3957\
        );

    \I__736\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3950\
        );

    \I__735\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3950\
        );

    \I__734\ : InMux
    port map (
            O => \N__3960\,
            I => \N__3950\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3957\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3950\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__731\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3939\
        );

    \I__730\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3939\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3939\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__728\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3931\
        );

    \I__727\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3928\
        );

    \I__726\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3925\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3931\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3928\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3925\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3918\,
            I => \N__3914\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3917\,
            I => \N__3909\
        );

    \I__720\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3904\
        );

    \I__719\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3904\
        );

    \I__718\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3901\
        );

    \I__717\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3898\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3904\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3898\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3888\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3888\,
            I => \N__3884\
        );

    \I__711\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3881\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__3884\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3881\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__708\ : InMux
    port map (
            O => \N__3876\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__707\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3870\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3870\,
            I => \N__3866\
        );

    \I__705\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3863\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__3866\,
            I => \N__3860\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3863\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__3860\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__701\ : InMux
    port map (
            O => \N__3855\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__700\ : InMux
    port map (
            O => \N__3852\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__699\ : InMux
    port map (
            O => \N__3849\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__698\ : InMux
    port map (
            O => \N__3846\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__697\ : InMux
    port map (
            O => \N__3843\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__695\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3833\
        );

    \I__694\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3830\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3827\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3830\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__3827\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__690\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3813\
        );

    \I__689\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3813\
        );

    \I__688\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3813\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3813\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__686\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3806\
        );

    \I__685\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3803\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3806\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3803\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__682\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3794\
        );

    \I__681\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3791\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3794\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3791\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__678\ : InMux
    port map (
            O => \N__3786\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__677\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3779\
        );

    \I__676\ : InMux
    port map (
            O => \N__3782\,
            I => \N__3776\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3779\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3776\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__673\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3768\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__671\ : InMux
    port map (
            O => \N__3765\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__670\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3758\
        );

    \I__669\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3755\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3758\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3755\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__666\ : InMux
    port map (
            O => \N__3750\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__665\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3743\
        );

    \I__664\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3740\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3743\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3740\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__661\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3732\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3732\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__659\ : InMux
    port map (
            O => \N__3729\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__658\ : InMux
    port map (
            O => \N__3726\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__3723\,
            I => \N__3720\
        );

    \I__656\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3716\
        );

    \I__655\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3713\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3716\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3713\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__652\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3705\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__650\ : InMux
    port map (
            O => \N__3702\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__649\ : InMux
    port map (
            O => \N__3699\,
            I => \bfn_10_7_0_\
        );

    \I__648\ : InMux
    port map (
            O => \N__3696\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__3693\,
            I => \U409_TICK.TICK603_11_cascade_\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__3690\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__645\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3684\,
            I => \U409_TICK.TICK603_8\
        );

    \I__643\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3677\
        );

    \I__642\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3674\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3677\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3674\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__639\ : InMux
    port map (
            O => \N__3669\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__638\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3659\
        );

    \I__637\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3656\
        );

    \I__636\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3649\
        );

    \I__635\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3649\
        );

    \I__634\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3649\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3659\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3656\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3649\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__630\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3638\
        );

    \I__629\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3635\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3638\,
            I => \U409_TRANSFER_ACK.N_97\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3635\,
            I => \U409_TRANSFER_ACK.N_97\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__3630\,
            I => \N__3626\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__3629\,
            I => \N__3623\
        );

    \I__624\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3620\
        );

    \I__623\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3615\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3620\,
            I => \N__3612\
        );

    \I__621\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3607\
        );

    \I__620\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3607\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3615\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__3612\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3607\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3600\,
            I => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\
        );

    \I__615\ : IoInMux
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__613\ : Span4Mux_s2_v
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__612\ : Span4Mux_h
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__610\ : Sp12to4
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__609\ : Span12Mux_h
    port map (
            O => \N__3579\,
            I => \N__3575\
        );

    \I__608\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3572\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__3575\,
            I => \TACK_OUTn\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3572\,
            I => \TACK_OUTn\
        );

    \I__605\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3563\
        );

    \I__604\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3560\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3563\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3560\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__601\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3546\
        );

    \I__600\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3546\
        );

    \I__599\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3546\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3546\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__3543\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\
        );

    \I__596\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3536\
        );

    \I__595\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3533\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3536\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3533\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3528\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__591\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3516\
        );

    \I__590\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3516\
        );

    \I__589\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3516\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3516\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__587\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3509\
        );

    \I__586\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3506\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3509\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3506\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__583\ : CEMux
    port map (
            O => \N__3501\,
            I => \N__3498\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3498\,
            I => \N__3495\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__3495\,
            I => \N__3492\
        );

    \I__580\ : Span4Mux_h
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__3489\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__3486\,
            I => \U409_TRANSFER_ACK.m9_bm_cascade_\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3483\,
            I => \U409_TRANSFER_ACK.N_4_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3477\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3477\,
            I => \U409_TRANSFER_ACK.m9_am\
        );

    \I__574\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3468\
        );

    \I__573\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3468\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3468\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__571\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3462\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__3459\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__568\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3450\
        );

    \I__567\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3447\
        );

    \I__566\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3442\
        );

    \I__565\ : InMux
    port map (
            O => \N__3453\,
            I => \N__3442\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3450\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3447\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3442\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__560\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3427\
        );

    \I__559\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3424\
        );

    \I__558\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3421\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3427\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3424\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3421\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__554\ : SRMux
    port map (
            O => \N__3414\,
            I => \N__3411\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__3408\,
            I => \U409_TRANSFER_ACK.RESETn_c_i\
        );

    \I__551\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3401\
        );

    \I__550\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3398\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3401\,
            I => \N__3393\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3398\,
            I => \N__3393\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__3393\,
            I => \CIA_ENABLEm\
        );

    \I__546\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3387\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3387\,
            I => \N__3383\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3386\,
            I => \N__3380\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__3383\,
            I => \N__3376\
        );

    \I__542\ : InMux
    port map (
            O => \N__3380\,
            I => \N__3373\
        );

    \I__541\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3370\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__3376\,
            I => \N__3363\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3363\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3370\,
            I => \N__3363\
        );

    \I__537\ : Span12Mux_h
    port map (
            O => \N__3363\,
            I => \N__3360\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__3360\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__535\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3353\
        );

    \I__534\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3350\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3353\,
            I => \N__3346\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3350\,
            I => \N__3343\
        );

    \I__531\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3340\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__3346\,
            I => \N__3337\
        );

    \I__529\ : Span4Mux_h
    port map (
            O => \N__3343\,
            I => \N__3332\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3340\,
            I => \N__3332\
        );

    \I__527\ : Span4Mux_v
    port map (
            O => \N__3337\,
            I => \N__3327\
        );

    \I__526\ : Span4Mux_v
    port map (
            O => \N__3332\,
            I => \N__3327\
        );

    \I__525\ : Sp12to4
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__524\ : Span12Mux_h
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__523\ : Odrv12
    port map (
            O => \N__3321\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__522\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3313\
        );

    \I__521\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3308\
        );

    \I__520\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3308\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3313\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3308\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__3303\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__3300\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\
        );

    \I__515\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3294\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__3291\,
            I => \N__3287\
        );

    \I__512\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3281\
        );

    \I__511\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3272\
        );

    \I__510\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3272\
        );

    \I__509\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3272\
        );

    \I__508\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3272\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3281\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3272\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__505\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3255\
        );

    \I__504\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3255\
        );

    \I__503\ : InMux
    port map (
            O => \N__3265\,
            I => \N__3255\
        );

    \I__502\ : InMux
    port map (
            O => \N__3264\,
            I => \N__3255\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3255\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__500\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3249\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\
        );

    \I__498\ : InMux
    port map (
            O => \N__3246\,
            I => \N__3241\
        );

    \I__497\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3238\
        );

    \I__496\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3235\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3241\,
            I => \N__3228\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3238\,
            I => \N__3228\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3235\,
            I => \N__3228\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__3228\,
            I => \N__3222\
        );

    \I__491\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3219\
        );

    \I__490\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3214\
        );

    \I__489\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3214\
        );

    \I__488\ : Sp12to4
    port map (
            O => \N__3222\,
            I => \N__3206\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3219\,
            I => \N__3206\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3214\,
            I => \N__3206\
        );

    \I__485\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3203\
        );

    \I__484\ : Span12Mux_h
    port map (
            O => \N__3206\,
            I => \N__3200\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3203\,
            I => \N__3197\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__3200\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__481\ : Odrv12
    port map (
            O => \N__3197\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__480\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3188\
        );

    \I__479\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3185\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3188\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3185\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__476\ : IoInMux
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__474\ : Span4Mux_s3_v
    port map (
            O => \N__3174\,
            I => \N__3171\
        );

    \I__473\ : Sp12to4
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__472\ : Span12Mux_h
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__471\ : Odrv12
    port map (
            O => \N__3165\,
            I => \ROMENm_i\
        );

    \I__470\ : IoInMux
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3159\,
            I => \N__3156\
        );

    \I__468\ : Span4Mux_s1_v
    port map (
            O => \N__3156\,
            I => \N__3153\
        );

    \I__467\ : Sp12to4
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__466\ : Span12Mux_h
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__465\ : Span12Mux_v
    port map (
            O => \N__3147\,
            I => \N__3144\
        );

    \I__464\ : Odrv12
    port map (
            O => \N__3144\,
            I => \PORTSIZE_0_i\
        );

    \I__463\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3131\
        );

    \I__462\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3131\
        );

    \I__461\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3131\
        );

    \I__460\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3126\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3131\,
            I => \N__3123\
        );

    \I__458\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3120\
        );

    \I__457\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3117\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3126\,
            I => \N__3114\
        );

    \I__455\ : Span4Mux_v
    port map (
            O => \N__3123\,
            I => \N__3111\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3120\,
            I => \N__3106\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3117\,
            I => \N__3106\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__3114\,
            I => \N__3103\
        );

    \I__451\ : Span4Mux_h
    port map (
            O => \N__3111\,
            I => \N__3098\
        );

    \I__450\ : Span4Mux_v
    port map (
            O => \N__3106\,
            I => \N__3098\
        );

    \I__449\ : Span4Mux_h
    port map (
            O => \N__3103\,
            I => \N__3095\
        );

    \I__448\ : Span4Mux_h
    port map (
            O => \N__3098\,
            I => \N__3092\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__3095\,
            I => \A_c_23\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__3092\,
            I => \A_c_23\
        );

    \I__445\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3081\
        );

    \I__444\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3081\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__3075\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__3072\,
            I => \N__3069\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__438\ : IoSpan4Mux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__437\ : Span4Mux_s2_v
    port map (
            O => \N__3063\,
            I => \N__3060\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__435\ : Span12Mux_v
    port map (
            O => \N__3057\,
            I => \N__3054\
        );

    \I__434\ : Span12Mux_h
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__3051\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__430\ : IoSpan4Mux
    port map (
            O => \N__3042\,
            I => \N__3039\
        );

    \I__429\ : Span4Mux_s2_v
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__428\ : Sp12to4
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__427\ : Span12Mux_v
    port map (
            O => \N__3033\,
            I => \N__3030\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__3030\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__425\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__3021\,
            I => \U409_ADDRESS_DECODE.un10_ROMENZ0\
        );

    \I__422\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3012\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\
        );

    \I__419\ : InMux
    port map (
            O => \N__3009\,
            I => \N__3004\
        );

    \I__418\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3001\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__3007\,
            I => \N__2998\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3004\,
            I => \N__2993\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3001\,
            I => \N__2993\
        );

    \I__414\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2990\
        );

    \I__413\ : Span4Mux_v
    port map (
            O => \N__2993\,
            I => \N__2985\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2990\,
            I => \N__2985\
        );

    \I__411\ : Span4Mux_h
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__2982\,
            I => \U409_ADDRESS_DECODE.un6_ROMENZ0\
        );

    \I__409\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2975\
        );

    \I__408\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2972\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2975\,
            I => \N__2966\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2966\
        );

    \I__405\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2963\
        );

    \I__404\ : Span4Mux_v
    port map (
            O => \N__2966\,
            I => \N__2960\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N__2957\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__2960\,
            I => \N__2954\
        );

    \I__401\ : Span12Mux_h
    port map (
            O => \N__2957\,
            I => \N__2951\
        );

    \I__400\ : Span12Mux_h
    port map (
            O => \N__2954\,
            I => \N__2948\
        );

    \I__399\ : Span12Mux_v
    port map (
            O => \N__2951\,
            I => \N__2945\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__2948\,
            I => \N__2942\
        );

    \I__397\ : Span12Mux_h
    port map (
            O => \N__2945\,
            I => \N__2939\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__2942\,
            I => \OVL_c\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__2939\,
            I => \OVL_c\
        );

    \I__394\ : InMux
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__391\ : Sp12to4
    port map (
            O => \N__2925\,
            I => \N__2922\
        );

    \I__390\ : Span12Mux_h
    port map (
            O => \N__2922\,
            I => \N__2919\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__2919\,
            I => \A_c_13\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__2916\,
            I => \N__2913\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2913\,
            I => \N__2910\
        );

    \I__386\ : IoSpan4Mux
    port map (
            O => \N__2910\,
            I => \N__2907\
        );

    \I__385\ : IoSpan4Mux
    port map (
            O => \N__2907\,
            I => \N__2904\
        );

    \I__384\ : Span4Mux_s3_h
    port map (
            O => \N__2904\,
            I => \N__2901\
        );

    \I__383\ : Sp12to4
    port map (
            O => \N__2901\,
            I => \N__2898\
        );

    \I__382\ : Span12Mux_s11_h
    port map (
            O => \N__2898\,
            I => \N__2895\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__2895\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__380\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2889\,
            I => \N__2886\
        );

    \I__378\ : Span12Mux_h
    port map (
            O => \N__2886\,
            I => \N__2883\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__2883\,
            I => \A_c_12\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__374\ : Span4Mux_s3_h
    port map (
            O => \N__2874\,
            I => \N__2871\
        );

    \I__373\ : Span4Mux_v
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__371\ : Sp12to4
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__370\ : Span12Mux_h
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__369\ : Odrv12
    port map (
            O => \N__2859\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__368\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2850\
        );

    \I__367\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2850\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__365\ : Span4Mux_h
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__364\ : Span4Mux_v
    port map (
            O => \N__2844\,
            I => \N__2841\
        );

    \I__363\ : Odrv4
    port map (
            O => \N__2841\,
            I => \A_c_29\
        );

    \I__362\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2832\
        );

    \I__361\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2832\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__359\ : Span4Mux_v
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__358\ : Span4Mux_h
    port map (
            O => \N__2826\,
            I => \N__2823\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__2823\,
            I => \A_c_30\
        );

    \I__356\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2817\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\
        );

    \I__354\ : InMux
    port map (
            O => \N__2814\,
            I => \N__2810\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2813\,
            I => \N__2807\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2810\,
            I => \N__2804\
        );

    \I__351\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2801\
        );

    \I__350\ : Span4Mux_v
    port map (
            O => \N__2804\,
            I => \N__2798\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2801\,
            I => \N__2795\
        );

    \I__348\ : Span4Mux_v
    port map (
            O => \N__2798\,
            I => \N__2790\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__2795\,
            I => \N__2790\
        );

    \I__346\ : Sp12to4
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__345\ : Odrv12
    port map (
            O => \N__2787\,
            I => \A_c_25\
        );

    \I__344\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2781\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__342\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2772\
        );

    \I__341\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2772\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__338\ : Sp12to4
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__337\ : Odrv12
    port map (
            O => \N__2763\,
            I => \A_c_27\
        );

    \I__336\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2754\
        );

    \I__335\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2754\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2754\,
            I => \N__2751\
        );

    \I__333\ : Span4Mux_v
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__331\ : Sp12to4
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__330\ : Odrv12
    port map (
            O => \N__2742\,
            I => \A_c_26\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__328\ : InMux
    port map (
            O => \N__2736\,
            I => \N__2730\
        );

    \I__327\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2730\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__325\ : Span4Mux_h
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__324\ : Span4Mux_v
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__323\ : Odrv4
    port map (
            O => \N__2721\,
            I => \A_c_24\
        );

    \I__322\ : InMux
    port map (
            O => \N__2718\,
            I => \N__2712\
        );

    \I__321\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2712\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__2709\,
            I => \N__2706\
        );

    \I__318\ : Sp12to4
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__2703\,
            I => \A_c_31\
        );

    \I__316\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2697\,
            I => \U409_CIA.g0Z0Z_2\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2694\,
            I => \N__2690\
        );

    \I__313\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2685\
        );

    \I__312\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2685\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__2682\,
            I => \N__2679\
        );

    \I__309\ : Span4Mux_v
    port map (
            O => \N__2679\,
            I => \N__2676\
        );

    \I__308\ : Sp12to4
    port map (
            O => \N__2676\,
            I => \N__2673\
        );

    \I__307\ : Odrv12
    port map (
            O => \N__2673\,
            I => \A_c_28\
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2670\,
            I => \U409_CIA.g0Z0Z_10_cascade_\
        );

    \I__305\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2661\
        );

    \I__304\ : InMux
    port map (
            O => \N__2666\,
            I => \N__2656\
        );

    \I__303\ : InMux
    port map (
            O => \N__2665\,
            I => \N__2656\
        );

    \I__302\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2653\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2661\,
            I => \N__2645\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2656\,
            I => \N__2645\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2653\,
            I => \N__2645\
        );

    \I__298\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2642\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__2645\,
            I => \N__2637\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2642\,
            I => \N__2637\
        );

    \I__295\ : Sp12to4
    port map (
            O => \N__2637\,
            I => \N__2634\
        );

    \I__294\ : Span12Mux_v
    port map (
            O => \N__2634\,
            I => \N__2631\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2631\,
            I => \A_c_22\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__291\ : InMux
    port map (
            O => \N__2625\,
            I => \N__2622\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2622\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\
        );

    \I__289\ : InMux
    port map (
            O => \N__2619\,
            I => \N__2616\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2616\,
            I => \N__2611\
        );

    \I__287\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2606\
        );

    \I__286\ : InMux
    port map (
            O => \N__2614\,
            I => \N__2606\
        );

    \I__285\ : Span4Mux_v
    port map (
            O => \N__2611\,
            I => \N__2603\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2606\,
            I => \N__2600\
        );

    \I__283\ : Sp12to4
    port map (
            O => \N__2603\,
            I => \N__2597\
        );

    \I__282\ : Span4Mux_h
    port map (
            O => \N__2600\,
            I => \N__2594\
        );

    \I__281\ : Span12Mux_h
    port map (
            O => \N__2597\,
            I => \N__2589\
        );

    \I__280\ : Sp12to4
    port map (
            O => \N__2594\,
            I => \N__2589\
        );

    \I__279\ : Span12Mux_v
    port map (
            O => \N__2589\,
            I => \N__2586\
        );

    \I__278\ : Odrv12
    port map (
            O => \N__2586\,
            I => \A_c_19\
        );

    \I__277\ : InMux
    port map (
            O => \N__2583\,
            I => \N__2580\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2580\,
            I => \N__2577\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2577\,
            I => \N__2574\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2574\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2571\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_\
        );

    \I__272\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2562\
        );

    \I__271\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2562\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2562\,
            I => \N__2559\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2559\,
            I => \N__2556\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__2556\,
            I => \N__2553\
        );

    \I__267\ : Span4Mux_v
    port map (
            O => \N__2553\,
            I => \N__2550\
        );

    \I__266\ : Sp12to4
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__265\ : Odrv12
    port map (
            O => \N__2547\,
            I => \A_c_18\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2544\,
            I => \N__2540\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2543\,
            I => \N__2537\
        );

    \I__262\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2532\
        );

    \I__261\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2532\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2532\,
            I => \N__2529\
        );

    \I__259\ : Span4Mux_h
    port map (
            O => \N__2529\,
            I => \N__2526\
        );

    \I__258\ : Sp12to4
    port map (
            O => \N__2526\,
            I => \N__2523\
        );

    \I__257\ : Span12Mux_v
    port map (
            O => \N__2523\,
            I => \N__2520\
        );

    \I__256\ : Odrv12
    port map (
            O => \N__2520\,
            I => \A_c_16\
        );

    \I__255\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2514\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2514\,
            I => \U409_CIA.g0Z0Z_11\
        );

    \I__253\ : CascadeMux
    port map (
            O => \N__2511\,
            I => \N__2508\
        );

    \I__252\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2504\
        );

    \I__251\ : InMux
    port map (
            O => \N__2507\,
            I => \N__2501\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2504\,
            I => \N__2498\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2501\,
            I => \N__2495\
        );

    \I__248\ : Span12Mux_s5_h
    port map (
            O => \N__2498\,
            I => \N__2490\
        );

    \I__247\ : Sp12to4
    port map (
            O => \N__2495\,
            I => \N__2490\
        );

    \I__246\ : Span12Mux_v
    port map (
            O => \N__2490\,
            I => \N__2487\
        );

    \I__245\ : Odrv12
    port map (
            O => \N__2487\,
            I => \A_c_17\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__2484\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\
        );

    \I__243\ : InMux
    port map (
            O => \N__2481\,
            I => \N__2475\
        );

    \I__242\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2475\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2475\,
            I => \N__2472\
        );

    \I__240\ : Odrv4
    port map (
            O => \N__2472\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__239\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2466\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2466\,
            I => \N__2462\
        );

    \I__237\ : CascadeMux
    port map (
            O => \N__2465\,
            I => \N__2459\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__2462\,
            I => \N__2455\
        );

    \I__235\ : InMux
    port map (
            O => \N__2459\,
            I => \N__2450\
        );

    \I__234\ : InMux
    port map (
            O => \N__2458\,
            I => \N__2450\
        );

    \I__233\ : Sp12to4
    port map (
            O => \N__2455\,
            I => \N__2445\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2450\,
            I => \N__2445\
        );

    \I__231\ : Odrv12
    port map (
            O => \N__2445\,
            I => \A_c_20\
        );

    \I__230\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2439\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2439\,
            I => \N__2436\
        );

    \I__228\ : Odrv4
    port map (
            O => \N__2436\,
            I => \U409_CIA.g0Z0Z_8\
        );

    \I__227\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2423\
        );

    \I__226\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2423\
        );

    \I__225\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2423\
        );

    \I__224\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2420\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2423\,
            I => \N__2415\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2420\,
            I => \N__2415\
        );

    \I__221\ : Span4Mux_v
    port map (
            O => \N__2415\,
            I => \N__2412\
        );

    \I__220\ : Span4Mux_h
    port map (
            O => \N__2412\,
            I => \N__2409\
        );

    \I__219\ : Odrv4
    port map (
            O => \N__2409\,
            I => \A_c_21\
        );

    \I__218\ : ClkMux
    port map (
            O => \N__2406\,
            I => \N__2373\
        );

    \I__217\ : ClkMux
    port map (
            O => \N__2405\,
            I => \N__2373\
        );

    \I__216\ : ClkMux
    port map (
            O => \N__2404\,
            I => \N__2373\
        );

    \I__215\ : ClkMux
    port map (
            O => \N__2403\,
            I => \N__2373\
        );

    \I__214\ : ClkMux
    port map (
            O => \N__2402\,
            I => \N__2373\
        );

    \I__213\ : ClkMux
    port map (
            O => \N__2401\,
            I => \N__2373\
        );

    \I__212\ : ClkMux
    port map (
            O => \N__2400\,
            I => \N__2373\
        );

    \I__211\ : ClkMux
    port map (
            O => \N__2399\,
            I => \N__2373\
        );

    \I__210\ : ClkMux
    port map (
            O => \N__2398\,
            I => \N__2373\
        );

    \I__209\ : ClkMux
    port map (
            O => \N__2397\,
            I => \N__2373\
        );

    \I__208\ : ClkMux
    port map (
            O => \N__2396\,
            I => \N__2373\
        );

    \I__207\ : GlobalMux
    port map (
            O => \N__2373\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            I => \N__2403\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2399\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2402\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2397\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2405\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            I => \N__2404\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2401\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__2398\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2396\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__2406\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2400\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2615\,
            in1 => \N__2814\,
            in2 => \N__2544\,
            in3 => \N__2568\,
            lcout => \U409_CIA.g0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2614\,
            in1 => \N__2567\,
            in2 => \N__2543\,
            in3 => \N__2507\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2517\,
            in1 => \N__2469\,
            in2 => \N__2511\,
            in3 => \N__2442\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2431\,
            in2 => \_gnd_net_\,
            in3 => \N__2458\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3213\,
            in1 => \N__2480\,
            in2 => \N__2484\,
            in3 => \N__2665\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2432\,
            in1 => \N__2481\,
            in2 => \N__2465\,
            in3 => \N__2666\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5541\,
            in1 => \N__3130\,
            in2 => \_gnd_net_\,
            in3 => \N__2433\,
            lcout => \U409_CIA.g0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un6_ROMEN_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2664\,
            in1 => \N__3129\,
            in2 => \_gnd_net_\,
            in3 => \N__2430\,
            lcout => \U409_ADDRESS_DECODE.un6_ROMENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__2820\,
            in1 => \N__2855\,
            in2 => \N__2694\,
            in3 => \N__2784\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2838\,
            lcout => \U409_CIA.g0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2717\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2759\,
            in1 => \N__2777\,
            in2 => \N__2813\,
            in3 => \N__2735\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2778\,
            in1 => \N__2760\,
            in2 => \N__2739\,
            in3 => \N__2718\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2700\,
            in1 => \N__2693\,
            in2 => \N__2670\,
            in3 => \N__2652\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3138\,
            in1 => \N__2667\,
            in2 => \N__2628\,
            in3 => \N__2619\,
            lcout => \U409_ADDRESS_DECODE.un10_ROMENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3140\,
            in1 => \N__3225\,
            in2 => \_gnd_net_\,
            in3 => \N__3086\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0\,
            ltout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__2583\,
            in1 => \N__3139\,
            in2 => \N__2571\,
            in3 => \N__5537\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3141\,
            in1 => \N__3226\,
            in2 => \_gnd_net_\,
            in3 => \N__3087\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__2971\,
            in1 => \N__3245\,
            in2 => \_gnd_net_\,
            in3 => \N__3009\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__3008\,
            in1 => \N__3027\,
            in2 => \_gnd_net_\,
            in3 => \N__2978\,
            lcout => \U409_ADDRESS_DECODE_un1_ROMEN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__3018\,
            in1 => \N__3227\,
            in2 => \N__3007\,
            in3 => \N__2979\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__2934\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3405\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__3404\,
            in1 => \N__2892\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__3356\,
            in1 => \N__3390\,
            in2 => \N__4320\,
            in3 => \N__3318\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__3414\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__3317\,
            in1 => \N__4312\,
            in2 => \N__3386\,
            in3 => \N__3357\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__3379\,
            in1 => \N__3349\,
            in2 => \N__4316\,
            in3 => \N__3316\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__3266\,
            in1 => \N__5522\,
            in2 => \N__3291\,
            in3 => \N__3252\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__3192\,
            in2 => \N__4599\,
            in3 => \N__3246\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100110011001"
        )
    port map (
            in0 => \N__3265\,
            in1 => \N__3290\,
            in2 => \N__3303\,
            in3 => \N__4679\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__5525\,
            in1 => \N__3285\,
            in2 => \N__3300\,
            in3 => \N__3540\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__3286\,
            in2 => \_gnd_net_\,
            in3 => \N__3267\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3297\,
            in1 => \N__3284\,
            in2 => \N__4687\,
            in3 => \N__3264\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__3244\,
            in1 => \N__3191\,
            in2 => \_gnd_net_\,
            in3 => \N__5529\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__3431\,
            in1 => \N__3455\,
            in2 => \N__3629\,
            in3 => \N__3642\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__5435\,
            in1 => \N__3666\,
            in2 => \N__3486\,
            in3 => \N__3480\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5513\,
            in2 => \_gnd_net_\,
            in3 => \N__3822\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3473\,
            in2 => \_gnd_net_\,
            in3 => \N__3820\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => \U409_TRANSFER_ACK.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__3618\,
            in1 => \N__3430\,
            in2 => \N__3483\,
            in3 => \N__3453\,
            lcout => \U409_TRANSFER_ACK.m9_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3662\,
            in1 => \N__3474\,
            in2 => \N__4683\,
            in3 => \N__3821\,
            lcout => \U409_TRANSFER_ACK.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110011"
        )
    port map (
            in0 => \N__3456\,
            in1 => \N__3465\,
            in2 => \N__3435\,
            in3 => \N__3663\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__3664\,
            in1 => \N__5512\,
            in2 => \N__3459\,
            in3 => \N__3619\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3454\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001000"
        )
    port map (
            in0 => \N__3665\,
            in1 => \N__3641\,
            in2 => \N__3630\,
            in3 => \N__3567\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5514\,
            in1 => \_gnd_net_\,
            in2 => \N__3600\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3525\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011101100"
        )
    port map (
            in0 => \N__3555\,
            in1 => \N__3578\,
            in2 => \N__5533\,
            in3 => \N__3513\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__3554\,
            in1 => \N__5520\,
            in2 => \_gnd_net_\,
            in3 => \N__3524\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3809\,
            in2 => \_gnd_net_\,
            in3 => \N__3566\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__3553\,
            in1 => \N__3523\,
            in2 => \N__3543\,
            in3 => \N__3539\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3528\,
            in3 => \N__5515\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5521\,
            in2 => \_gnd_net_\,
            in3 => \N__3512\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__3501\,
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__4090\,
            in1 => \N__3735\,
            in2 => \N__4026\,
            in3 => \N__4062\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4013\,
            in1 => \N__4091\,
            in2 => \N__4065\,
            in3 => \N__3708\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3873\,
            in1 => \N__3681\,
            in2 => \N__3840\,
            in3 => \N__3935\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3687\,
            in1 => \N__3891\,
            in2 => \N__3693\,
            in3 => \N__3798\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4089\,
            in1 => \N__4058\,
            in2 => \N__3690\,
            in3 => \N__3771\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__3762\,
            in1 => \N__3783\,
            in2 => \_gnd_net_\,
            in3 => \N__3912\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3747\,
            in1 => \N__4167\,
            in2 => \N__3723\,
            in3 => \N__4239\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3934\,
            in2 => \N__3917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3680\,
            in2 => \_gnd_net_\,
            in3 => \N__3669\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__5304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3797\,
            in2 => \_gnd_net_\,
            in3 => \N__3786\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__5304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3782\,
            in2 => \_gnd_net_\,
            in3 => \N__3765\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3761\,
            in2 => \_gnd_net_\,
            in3 => \N__3750\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__5304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3746\,
            in2 => \_gnd_net_\,
            in3 => \N__3729\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4124\,
            in2 => \_gnd_net_\,
            in3 => \N__3726\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__5304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3719\,
            in2 => \_gnd_net_\,
            in3 => \N__3702\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4166\,
            in2 => \_gnd_net_\,
            in3 => \N__3699\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4142\,
            in2 => \_gnd_net_\,
            in3 => \N__3696\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3887\,
            in2 => \_gnd_net_\,
            in3 => \N__3876\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3869\,
            in2 => \_gnd_net_\,
            in3 => \N__3855\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4154\,
            in2 => \_gnd_net_\,
            in3 => \N__3852\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4238\,
            in2 => \_gnd_net_\,
            in3 => \N__3849\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4112\,
            in2 => \_gnd_net_\,
            in3 => \N__3846\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3836\,
            in2 => \_gnd_net_\,
            in3 => \N__3843\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5468\,
            in2 => \_gnd_net_\,
            in3 => \N__4256\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__4597\,
            in2 => \N__4688\,
            in3 => \N__4797\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5367\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__3810\,
            in1 => \N__4538\,
            in2 => \_gnd_net_\,
            in3 => \N__4553\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5367\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4798\,
            in1 => \N__3967\,
            in2 => \_gnd_net_\,
            in3 => \N__4764\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5367\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4761\,
            in1 => \N__4514\,
            in2 => \N__3968\,
            in3 => \N__4795\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4762\,
            in1 => \_gnd_net_\,
            in2 => \N__3969\,
            in3 => \N__4796\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4710\,
            in1 => \N__4513\,
            in2 => \N__4800\,
            in3 => \N__4738\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \N__5022\,
            in2 => \N__3975\,
            in3 => \N__3944\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5021\,
            in1 => \N__4512\,
            in2 => \N__5004\,
            in3 => \N__4739\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4711\,
            in1 => \N__4794\,
            in2 => \N__3972\,
            in3 => \N__3945\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4760\,
            in2 => \_gnd_net_\,
            in3 => \N__3960\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3913\,
            in2 => \_gnd_net_\,
            in3 => \N__3936\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4063\,
            in2 => \N__3918\,
            in3 => \N__4014\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__4015\,
            in1 => \N__4064\,
            in2 => \N__4100\,
            in3 => \N__4193\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4421\,
            in1 => \N__4454\,
            in2 => \N__4389\,
            in3 => \N__4854\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__4833\,
            in1 => \N__4422\,
            in2 => \N__4458\,
            in3 => \N__4387\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__4943\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5193\,
            in1 => \N__4920\,
            in2 => \N__4962\,
            in3 => \N__5318\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4027\,
            in1 => \N__4057\,
            in2 => \N__4101\,
            in3 => \N__4182\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4056\,
            in1 => \N__4029\,
            in2 => \N__4176\,
            in3 => \N__4099\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4155\,
            in1 => \N__4143\,
            in2 => \N__4131\,
            in3 => \N__4113\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4055\,
            in1 => \N__4028\,
            in2 => \N__3984\,
            in3 => \N__3981\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4866\,
            in1 => \N__4905\,
            in2 => \_gnd_net_\,
            in3 => \N__4941\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__5109\,
            in2 => \N__4221\,
            in3 => \N__5151\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4415\,
            in1 => \N__4378\,
            in2 => \N__4218\,
            in3 => \N__5061\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4377\,
            in1 => \N__4452\,
            in2 => \N__5040\,
            in3 => \N__4417\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5073\,
            in1 => \N__4824\,
            in2 => \N__4890\,
            in3 => \N__5052\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4376\,
            in1 => \N__4451\,
            in2 => \N__4215\,
            in3 => \N__5082\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5094\,
            in1 => \N__4845\,
            in2 => \N__5136\,
            in3 => \N__5175\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4942\,
            in1 => \N__4416\,
            in2 => \N__4212\,
            in3 => \N__4453\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4418\,
            in1 => \N__4449\,
            in2 => \N__5121\,
            in3 => \N__4382\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4419\,
            in1 => \N__4383\,
            in2 => \N__5163\,
            in3 => \N__4450\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__4448\,
            in1 => \N__4420\,
            in2 => \N__4388\,
            in3 => \N__4334\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5259\,
            in1 => \N__5216\,
            in2 => \N__5751\,
            in3 => \N__5673\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5711\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__5708\,
            in2 => \_gnd_net_\,
            in3 => \N__5239\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__4308\,
            in1 => \N__5672\,
            in2 => \N__4323\,
            in3 => \N__4809\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5670\,
            in1 => \N__5707\,
            in2 => \_gnd_net_\,
            in3 => \N__5238\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4255\,
            in2 => \N__4287\,
            in3 => \N__4808\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__4284\,
            in1 => \N__5709\,
            in2 => \N__4278\,
            in3 => \N__5241\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5745\,
            in1 => \N__5211\,
            in2 => \_gnd_net_\,
            in3 => \N__5258\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4799\,
            in1 => \N__4763\,
            in2 => \_gnd_net_\,
            in3 => \N__4481\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5366\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4740\,
            in1 => \N__4713\,
            in2 => \N__4725\,
            in3 => \N__4480\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5365\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4492\,
            in1 => \N__4999\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4712\,
            in2 => \N__4716\,
            in3 => \N__4476\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5365\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__4652\,
            in1 => \N__4598\,
            in2 => \N__4554\,
            in3 => \N__4537\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5024\,
            in1 => \_gnd_net_\,
            in2 => \N__4524\,
            in3 => \N__4493\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5365\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4521\,
            in1 => \N__4515\,
            in2 => \_gnd_net_\,
            in3 => \N__4475\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5365\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__4494\,
            in1 => \N__5000\,
            in2 => \N__4482\,
            in3 => \N__5025\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__5365\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4957\,
            in2 => \N__4944\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4919\,
            in2 => \_gnd_net_\,
            in3 => \N__4908\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__5300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4904\,
            in2 => \_gnd_net_\,
            in3 => \N__4893\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__5300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4880\,
            in2 => \_gnd_net_\,
            in3 => \N__4869\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__5300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4865\,
            in2 => \_gnd_net_\,
            in3 => \N__4848\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4844\,
            in2 => \_gnd_net_\,
            in3 => \N__4827\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4823\,
            in2 => \_gnd_net_\,
            in3 => \N__4812\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__5300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5189\,
            in2 => \_gnd_net_\,
            in3 => \N__5178\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__5300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5174\,
            in2 => \_gnd_net_\,
            in3 => \N__5154\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5150\,
            in2 => \_gnd_net_\,
            in3 => \N__5139\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__5303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5132\,
            in2 => \_gnd_net_\,
            in3 => \N__5112\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5108\,
            in2 => \_gnd_net_\,
            in3 => \N__5097\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__5303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5093\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5072\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5051\,
            in2 => \_gnd_net_\,
            in3 => \N__5028\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5319\,
            in2 => \_gnd_net_\,
            in3 => \N__5322\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5710\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5642\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5236\,
            in2 => \N__5712\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5256\,
            in2 => \_gnd_net_\,
            in3 => \N__5274\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__5640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__5271\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5212\,
            in2 => \_gnd_net_\,
            in3 => \N__5268\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__5640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5750\,
            in2 => \_gnd_net_\,
            in3 => \N__5265\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__5669\,
            in1 => \N__5727\,
            in2 => \N__5262\,
            in3 => \N__5705\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5257\,
            in1 => \N__5237\,
            in2 => \N__5217\,
            in3 => \N__5749\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011001100110"
        )
    port map (
            in0 => \N__5668\,
            in1 => \N__5721\,
            in2 => \N__5715\,
            in3 => \N__5706\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5625\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_353_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5576\,
            in1 => \N__5556\,
            in2 => \_gnd_net_\,
            in3 => \N__5459\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 30 2025 12:31:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    SIZ,
    DRA,
    A,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [1:0] SIZ;
    input [9:0] DRA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12142;
    wire N__12141;
    wire N__12140;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12088;
    wire N__12087;
    wire N__12086;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12070;
    wire N__12069;
    wire N__12068;
    wire N__12061;
    wire N__12060;
    wire N__12059;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12034;
    wire N__12033;
    wire N__12032;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12016;
    wire N__12015;
    wire N__12014;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11971;
    wire N__11970;
    wire N__11969;
    wire N__11962;
    wire N__11961;
    wire N__11960;
    wire N__11953;
    wire N__11952;
    wire N__11951;
    wire N__11944;
    wire N__11943;
    wire N__11942;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11917;
    wire N__11916;
    wire N__11915;
    wire N__11908;
    wire N__11907;
    wire N__11906;
    wire N__11899;
    wire N__11898;
    wire N__11897;
    wire N__11890;
    wire N__11889;
    wire N__11888;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11863;
    wire N__11862;
    wire N__11861;
    wire N__11854;
    wire N__11853;
    wire N__11852;
    wire N__11845;
    wire N__11844;
    wire N__11843;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11827;
    wire N__11826;
    wire N__11825;
    wire N__11818;
    wire N__11817;
    wire N__11816;
    wire N__11809;
    wire N__11808;
    wire N__11807;
    wire N__11800;
    wire N__11799;
    wire N__11798;
    wire N__11791;
    wire N__11790;
    wire N__11789;
    wire N__11782;
    wire N__11781;
    wire N__11780;
    wire N__11773;
    wire N__11772;
    wire N__11771;
    wire N__11764;
    wire N__11763;
    wire N__11762;
    wire N__11755;
    wire N__11754;
    wire N__11753;
    wire N__11746;
    wire N__11745;
    wire N__11744;
    wire N__11737;
    wire N__11736;
    wire N__11735;
    wire N__11728;
    wire N__11727;
    wire N__11726;
    wire N__11719;
    wire N__11718;
    wire N__11717;
    wire N__11710;
    wire N__11709;
    wire N__11708;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11692;
    wire N__11691;
    wire N__11690;
    wire N__11683;
    wire N__11682;
    wire N__11681;
    wire N__11674;
    wire N__11673;
    wire N__11672;
    wire N__11665;
    wire N__11664;
    wire N__11663;
    wire N__11656;
    wire N__11655;
    wire N__11654;
    wire N__11647;
    wire N__11646;
    wire N__11645;
    wire N__11638;
    wire N__11637;
    wire N__11636;
    wire N__11629;
    wire N__11628;
    wire N__11627;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11557;
    wire N__11556;
    wire N__11555;
    wire N__11548;
    wire N__11547;
    wire N__11546;
    wire N__11539;
    wire N__11538;
    wire N__11537;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11521;
    wire N__11520;
    wire N__11519;
    wire N__11512;
    wire N__11511;
    wire N__11510;
    wire N__11503;
    wire N__11502;
    wire N__11501;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11485;
    wire N__11484;
    wire N__11483;
    wire N__11476;
    wire N__11475;
    wire N__11474;
    wire N__11467;
    wire N__11466;
    wire N__11465;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11440;
    wire N__11439;
    wire N__11438;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11422;
    wire N__11421;
    wire N__11420;
    wire N__11413;
    wire N__11412;
    wire N__11411;
    wire N__11404;
    wire N__11403;
    wire N__11402;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11386;
    wire N__11385;
    wire N__11384;
    wire N__11377;
    wire N__11376;
    wire N__11375;
    wire N__11368;
    wire N__11367;
    wire N__11366;
    wire N__11349;
    wire N__11346;
    wire N__11345;
    wire N__11342;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11299;
    wire N__11296;
    wire N__11291;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11267;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11211;
    wire N__11210;
    wire N__11209;
    wire N__11206;
    wire N__11205;
    wire N__11202;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11180;
    wire N__11177;
    wire N__11172;
    wire N__11169;
    wire N__11164;
    wire N__11161;
    wire N__11156;
    wire N__11151;
    wire N__11148;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11137;
    wire N__11136;
    wire N__11133;
    wire N__11132;
    wire N__11129;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11101;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11095;
    wire N__11094;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11075;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11023;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11000;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10929;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10923;
    wire N__10920;
    wire N__10915;
    wire N__10912;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10851;
    wire N__10850;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10827;
    wire N__10826;
    wire N__10825;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10799;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10762;
    wire N__10755;
    wire N__10752;
    wire N__10747;
    wire N__10744;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10679;
    wire N__10678;
    wire N__10677;
    wire N__10676;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10659;
    wire N__10658;
    wire N__10569;
    wire N__10566;
    wire N__10565;
    wire N__10562;
    wire N__10561;
    wire N__10560;
    wire N__10557;
    wire N__10556;
    wire N__10555;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10547;
    wire N__10544;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10464;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10456;
    wire N__10455;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10419;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10362;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10326;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10315;
    wire N__10312;
    wire N__10311;
    wire N__10310;
    wire N__10309;
    wire N__10308;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10300;
    wire N__10299;
    wire N__10298;
    wire N__10297;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10289;
    wire N__10288;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10236;
    wire N__10227;
    wire N__10222;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10187;
    wire N__10180;
    wire N__10175;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10149;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10093;
    wire N__10092;
    wire N__10091;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10067;
    wire N__10066;
    wire N__10065;
    wire N__10064;
    wire N__10063;
    wire N__10062;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10058;
    wire N__10057;
    wire N__10056;
    wire N__10055;
    wire N__10054;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10016;
    wire N__10015;
    wire N__10014;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9994;
    wire N__9993;
    wire N__9992;
    wire N__9991;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9986;
    wire N__9985;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9975;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9744;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9678;
    wire N__9673;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9643;
    wire N__9642;
    wire N__9641;
    wire N__9638;
    wire N__9633;
    wire N__9632;
    wire N__9629;
    wire N__9624;
    wire N__9621;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9582;
    wire N__9579;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9563;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9557;
    wire N__9552;
    wire N__9547;
    wire N__9546;
    wire N__9543;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9529;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9466;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9442;
    wire N__9439;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9384;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9374;
    wire N__9371;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9343;
    wire N__9342;
    wire N__9337;
    wire N__9334;
    wire N__9333;
    wire N__9332;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9320;
    wire N__9317;
    wire N__9310;
    wire N__9305;
    wire N__9300;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9280;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9212;
    wire N__9209;
    wire N__9208;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9015;
    wire N__9012;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8900;
    wire N__8899;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8885;
    wire N__8882;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8842;
    wire N__8837;
    wire N__8836;
    wire N__8831;
    wire N__8830;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8824;
    wire N__8823;
    wire N__8822;
    wire N__8821;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8810;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8792;
    wire N__8789;
    wire N__8788;
    wire N__8787;
    wire N__8784;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8754;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8727;
    wire N__8718;
    wire N__8709;
    wire N__8704;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8639;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8618;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8591;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8528;
    wire N__8525;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8486;
    wire N__8483;
    wire N__8482;
    wire N__8481;
    wire N__8480;
    wire N__8479;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8465;
    wire N__8460;
    wire N__8451;
    wire N__8448;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8436;
    wire N__8435;
    wire N__8434;
    wire N__8431;
    wire N__8426;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8409;
    wire N__8404;
    wire N__8401;
    wire N__8400;
    wire N__8399;
    wire N__8398;
    wire N__8397;
    wire N__8396;
    wire N__8395;
    wire N__8394;
    wire N__8389;
    wire N__8386;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8368;
    wire N__8365;
    wire N__8352;
    wire N__8351;
    wire N__8348;
    wire N__8347;
    wire N__8346;
    wire N__8343;
    wire N__8342;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8327;
    wire N__8324;
    wire N__8317;
    wire N__8310;
    wire N__8309;
    wire N__8308;
    wire N__8307;
    wire N__8306;
    wire N__8305;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8300;
    wire N__8297;
    wire N__8296;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8277;
    wire N__8276;
    wire N__8273;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8250;
    wire N__8247;
    wire N__8242;
    wire N__8239;
    wire N__8232;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8216;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8208;
    wire N__8203;
    wire N__8202;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8191;
    wire N__8190;
    wire N__8189;
    wire N__8188;
    wire N__8187;
    wire N__8186;
    wire N__8181;
    wire N__8176;
    wire N__8173;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8161;
    wire N__8156;
    wire N__8153;
    wire N__8148;
    wire N__8141;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8129;
    wire N__8128;
    wire N__8127;
    wire N__8126;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8115;
    wire N__8104;
    wire N__8101;
    wire N__8096;
    wire N__8095;
    wire N__8092;
    wire N__8085;
    wire N__8078;
    wire N__8075;
    wire N__8074;
    wire N__8073;
    wire N__8072;
    wire N__8071;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8049;
    wire N__8044;
    wire N__8037;
    wire N__8030;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8001;
    wire N__8000;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7952;
    wire N__7949;
    wire N__7948;
    wire N__7945;
    wire N__7940;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7651;
    wire N__7648;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7630;
    wire N__7627;
    wire N__7614;
    wire N__7613;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7598;
    wire N__7595;
    wire N__7594;
    wire N__7593;
    wire N__7592;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7578;
    wire N__7575;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7455;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7386;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7378;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7353;
    wire N__7352;
    wire N__7349;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7322;
    wire N__7321;
    wire N__7318;
    wire N__7313;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7260;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7208;
    wire N__7205;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7185;
    wire N__7182;
    wire N__7181;
    wire N__7180;
    wire N__7179;
    wire N__7176;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7159;
    wire N__7158;
    wire N__7157;
    wire N__7156;
    wire N__7155;
    wire N__7154;
    wire N__7153;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7145;
    wire N__7144;
    wire N__7139;
    wire N__7134;
    wire N__7133;
    wire N__7130;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7065;
    wire N__7064;
    wire N__7061;
    wire N__7060;
    wire N__7059;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7051;
    wire N__7050;
    wire N__7049;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7040;
    wire N__7039;
    wire N__7034;
    wire N__7031;
    wire N__7026;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7022;
    wire N__7021;
    wire N__7020;
    wire N__7019;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6990;
    wire N__6985;
    wire N__6976;
    wire N__6971;
    wire N__6948;
    wire N__6947;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6941;
    wire N__6938;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6926;
    wire N__6923;
    wire N__6922;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6901;
    wire N__6888;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6869;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6855;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6824;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6788;
    wire N__6787;
    wire N__6786;
    wire N__6783;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6768;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6752;
    wire N__6749;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6730;
    wire N__6725;
    wire N__6724;
    wire N__6719;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6699;
    wire N__6698;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6681;
    wire N__6680;
    wire N__6679;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6666;
    wire N__6663;
    wire N__6662;
    wire N__6661;
    wire N__6660;
    wire N__6659;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6629;
    wire N__6624;
    wire N__6615;
    wire N__6600;
    wire N__6599;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6591;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6583;
    wire N__6576;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6565;
    wire N__6564;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6552;
    wire N__6547;
    wire N__6542;
    wire N__6539;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6490;
    wire N__6487;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6476;
    wire N__6471;
    wire N__6470;
    wire N__6465;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6431;
    wire N__6428;
    wire N__6423;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6368;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6356;
    wire N__6355;
    wire N__6352;
    wire N__6347;
    wire N__6344;
    wire N__6343;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6332;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6298;
    wire N__6295;
    wire N__6290;
    wire N__6287;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6252;
    wire N__6249;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6236;
    wire N__6235;
    wire N__6234;
    wire N__6233;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6199;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6166;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6143;
    wire N__6142;
    wire N__6141;
    wire N__6140;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6123;
    wire N__6120;
    wire N__6115;
    wire N__6110;
    wire N__6103;
    wire N__6098;
    wire N__6095;
    wire N__6090;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6048;
    wire N__6047;
    wire N__6042;
    wire N__6041;
    wire N__6038;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5885;
    wire N__5884;
    wire N__5883;
    wire N__5882;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5853;
    wire N__5846;
    wire N__5843;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5747;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5717;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5664;
    wire N__5661;
    wire N__5660;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5627;
    wire N__5624;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5613;
    wire N__5606;
    wire N__5603;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5579;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5538;
    wire N__5535;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5502;
    wire N__5499;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5487;
    wire N__5484;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5472;
    wire N__5471;
    wire N__5470;
    wire N__5469;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5465;
    wire N__5464;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5379;
    wire N__5376;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5364;
    wire N__5361;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5349;
    wire N__5346;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5331;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5316;
    wire N__5313;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5301;
    wire N__5298;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5264;
    wire N__5261;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5236;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5220;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5161;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5141;
    wire N__5136;
    wire N__5133;
    wire N__5124;
    wire N__5121;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5096;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5010;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4769;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4745;
    wire N__4744;
    wire N__4741;
    wire N__4736;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4699;
    wire N__4694;
    wire N__4691;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4674;
    wire N__4671;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4403;
    wire N__4402;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire N_861_i;
    wire DBRn_c;
    wire DBRn_c_i;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire VBENn_c;
    wire A_c_14;
    wire A_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0 ;
    wire DBDIR_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CHIP_RAM.DBENn_8_0 ;
    wire \U712_CHIP_RAM.N_341 ;
    wire \U712_CHIP_RAM.N_341_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ;
    wire A_c_20;
    wire TACK_EN_i_ess;
    wire TACK_OUTn;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.N_387_cascade_ ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_186_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_387 ;
    wire \U712_CHIP_RAM.N_385_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ;
    wire \U712_CHIP_RAM.N_223 ;
    wire \U712_CHIP_RAM.N_335_cascade_ ;
    wire \U712_CHIP_RAM.N_342_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_6_0_a2_2 ;
    wire \U712_CHIP_RAM.CLK_EN_6_0_a2_1 ;
    wire \U712_CHIP_RAM.CLK_EN_6_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ;
    wire \U712_CHIP_RAM.N_385 ;
    wire \U712_CHIP_RAM.N_338_cascade_ ;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire \U712_CHIP_RAM.N_239_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_208 ;
    wire \U712_CYCLE_TERM.N_217_i_0_en_0 ;
    wire ASn_c;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire RAMENn_c;
    wire \U712_REG_SM.N_270_cascade_ ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.N_289 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_3 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_ ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_4 ;
    wire \U712_CHIP_RAM.N_186 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_306 ;
    wire \U712_CHIP_RAM.N_333_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ;
    wire \U712_CHIP_RAM.N_239 ;
    wire \U712_CHIP_RAM.N_269 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire bfn_10_12_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_46 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CYCLE_TERM.N_217_i_0_en ;
    wire \U712_REG_SM.START_RST_0_sqmuxa ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire \U712_REG_SM.N_285_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ;
    wire \U712_REG_SM.N_222 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_284_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_10_15_0_;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.N_134 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire N_116_i;
    wire \U712_CHIP_RAM.N_207_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_ ;
    wire \U712_CHIP_RAM.N_333 ;
    wire \U712_CHIP_RAM.N_310_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ;
    wire DMA_CYCLEm;
    wire DBENn_c;
    wire \U712_CHIP_RAM.N_334 ;
    wire \U712_CHIP_RAM.N_297 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0 ;
    wire \U712_CHIP_RAM.N_202 ;
    wire \U712_CHIP_RAM.N_184_cascade_ ;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_392_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0 ;
    wire \U712_REG_SM.N_196 ;
    wire \U712_REG_SM.N_383 ;
    wire \U712_REG_SM.N_383_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_321_cascade_ ;
    wire CPU_TACKm;
    wire N_156_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0 ;
    wire N_126_i;
    wire \U712_BYTE_ENABLE.N_315 ;
    wire \U712_BYTE_ENABLE.N_319 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire \U712_REG_SM.un1_STATE_COUNT_4_i_i_0 ;
    wire \U712_REG_SM.N_26 ;
    wire \U712_REG_SM.N_274 ;
    wire DMA_LATCH_EN_c;
    wire CONSTANT_ONE_NET;
    wire A_c_15;
    wire A_c_8;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.N_207 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_262 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0 ;
    wire \U712_CHIP_RAM.N_237 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0 ;
    wire \U712_CHIP_RAM.N_335 ;
    wire \U712_CHIP_RAM.N_261 ;
    wire \U712_CHIP_RAM.N_180 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_386 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_338 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2 ;
    wire \U712_CHIP_RAM.N_342 ;
    wire \U712_CHIP_RAM.N_293_cascade_ ;
    wire \U712_CHIP_RAM.N_294 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_235_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_REG_SM.N_281 ;
    wire \U712_REG_SM.N_235 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_REG_SM.N_212 ;
    wire \U712_REG_SM.REG_TACK_RNOZ0Z_0 ;
    wire REG_TACK;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_220_cascade_ ;
    wire N_151_i;
    wire \U712_BYTE_ENABLE.N_314 ;
    wire \U712_BYTE_ENABLE.UUBE ;
    wire RESETn_c_i;
    wire WEn_c;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire A_c_16;
    wire A_c_18;
    wire \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire A_c_6;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_236_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_273 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire A_c_19;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire CMA_c_9;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire UMBEn_c;
    wire U712_BYTE_ENABLE_UUBE_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire U712_BYTE_ENABLE_un1_UDSn_i;
    wire LLBEn_c;
    wire DS_ENm;
    wire N_119;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire N_220_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire RAS0n_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire DRA_c_6;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_3;
    wire AGNUS_REV_c;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire RnW_c;
    wire CASUn_c;
    wire CASLn_c;
    wire WRITE_CYCLEm;
    wire N_238;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4113),
            .RESETB(N__5976),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12169),
            .DIN(N__12168),
            .DOUT(N__12167),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12169),
            .PADOUT(N__12168),
            .PADIN(N__12167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5586),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12160),
            .DIN(N__12159),
            .DOUT(N__12158),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12160),
            .PADOUT(N__12159),
            .PADIN(N__12158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12151),
            .DIN(N__12150),
            .DOUT(N__12149),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12151),
            .PADOUT(N__12150),
            .PADIN(N__12149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9246),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12142),
            .DIN(N__12141),
            .DOUT(N__12140),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12142),
            .PADOUT(N__12141),
            .PADIN(N__12140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12133),
            .DIN(N__12132),
            .DOUT(N__12131),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12133),
            .PADOUT(N__12132),
            .PADIN(N__12131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12124),
            .DIN(N__12123),
            .DOUT(N__12122),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12124),
            .PADOUT(N__12123),
            .PADIN(N__12122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12115),
            .DIN(N__12114),
            .DOUT(N__12113),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12115),
            .PADOUT(N__12114),
            .PADIN(N__12113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12106),
            .DIN(N__12105),
            .DOUT(N__12104),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12106),
            .PADOUT(N__12105),
            .PADIN(N__12104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12097),
            .DIN(N__12096),
            .DOUT(N__12095),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12097),
            .PADOUT(N__12096),
            .PADIN(N__12095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12088),
            .DIN(N__12087),
            .DOUT(N__12086),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12088),
            .PADOUT(N__12087),
            .PADIN(N__12086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12079),
            .DIN(N__12078),
            .DOUT(N__12077),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12079),
            .PADOUT(N__12078),
            .PADIN(N__12077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8979),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12070),
            .DIN(N__12069),
            .DOUT(N__12068),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12070),
            .PADOUT(N__12069),
            .PADIN(N__12068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12061),
            .DIN(N__12060),
            .DOUT(N__12059),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12061),
            .PADOUT(N__12060),
            .PADIN(N__12059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12052),
            .DIN(N__12051),
            .DOUT(N__12050),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12052),
            .PADOUT(N__12051),
            .PADIN(N__12050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12043),
            .DIN(N__12042),
            .DOUT(N__12041),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12043),
            .PADOUT(N__12042),
            .PADIN(N__12041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12034),
            .DIN(N__12033),
            .DOUT(N__12032),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12034),
            .PADOUT(N__12033),
            .PADIN(N__12032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12025),
            .DIN(N__12024),
            .DOUT(N__12023),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12025),
            .PADOUT(N__12024),
            .PADIN(N__12023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12016),
            .DIN(N__12015),
            .DOUT(N__12014),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12016),
            .PADOUT(N__12015),
            .PADIN(N__12014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12007),
            .DIN(N__12006),
            .DOUT(N__12005),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12007),
            .PADOUT(N__12006),
            .PADIN(N__12005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11998),
            .DIN(N__11997),
            .DOUT(N__11996),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11998),
            .PADOUT(N__11997),
            .PADIN(N__11996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11049),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11989),
            .DIN(N__11988),
            .DOUT(N__11987),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11989),
            .PADOUT(N__11988),
            .PADIN(N__11987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11980),
            .DIN(N__11979),
            .DOUT(N__11978),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11980),
            .PADOUT(N__11979),
            .PADIN(N__11978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9003),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11971),
            .DIN(N__11970),
            .DOUT(N__11969),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11971),
            .PADOUT(N__11970),
            .PADIN(N__11969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11962),
            .DIN(N__11961),
            .DOUT(N__11960),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11962),
            .PADOUT(N__11961),
            .PADIN(N__11960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9774),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11953),
            .DIN(N__11952),
            .DOUT(N__11951),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11953),
            .PADOUT(N__11952),
            .PADIN(N__11951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11944),
            .DIN(N__11943),
            .DOUT(N__11942),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11944),
            .PADOUT(N__11943),
            .PADIN(N__11942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11935),
            .DIN(N__11934),
            .DOUT(N__11933),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11935),
            .PADOUT(N__11934),
            .PADIN(N__11933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11926),
            .DIN(N__11925),
            .DOUT(N__11924),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11926),
            .PADOUT(N__11925),
            .PADIN(N__11924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11917),
            .DIN(N__11916),
            .DOUT(N__11915),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11917),
            .PADOUT(N__11916),
            .PADIN(N__11915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11908),
            .DIN(N__11907),
            .DOUT(N__11906),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11908),
            .PADOUT(N__11907),
            .PADIN(N__11906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5997),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11899),
            .DIN(N__11898),
            .DOUT(N__11897),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11899),
            .PADOUT(N__11898),
            .PADIN(N__11897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11890),
            .DIN(N__11889),
            .DOUT(N__11888),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11890),
            .PADOUT(N__11889),
            .PADIN(N__11888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11881),
            .DIN(N__11880),
            .DOUT(N__11879),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11881),
            .PADOUT(N__11880),
            .PADIN(N__11879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11872),
            .DIN(N__11871),
            .DOUT(N__11870),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11872),
            .PADOUT(N__11871),
            .PADIN(N__11870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11863),
            .DIN(N__11862),
            .DOUT(N__11861),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11863),
            .PADOUT(N__11862),
            .PADIN(N__11861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11854),
            .DIN(N__11853),
            .DOUT(N__11852),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11854),
            .PADOUT(N__11853),
            .PADIN(N__11852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7698),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11845),
            .DIN(N__11844),
            .DOUT(N__11843),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11845),
            .PADOUT(N__11844),
            .PADIN(N__11843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4986),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11836),
            .DIN(N__11835),
            .DOUT(N__11834),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11836),
            .PADOUT(N__11835),
            .PADIN(N__11834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11827),
            .DIN(N__11826),
            .DOUT(N__11825),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11827),
            .PADOUT(N__11826),
            .PADIN(N__11825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4722),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11818),
            .DIN(N__11817),
            .DOUT(N__11816),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11818),
            .PADOUT(N__11817),
            .PADIN(N__11816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11809),
            .DIN(N__11808),
            .DOUT(N__11807),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11809),
            .PADOUT(N__11808),
            .PADIN(N__11807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11800),
            .DIN(N__11799),
            .DOUT(N__11798),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11800),
            .PADOUT(N__11799),
            .PADIN(N__11798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11791),
            .DIN(N__11790),
            .DOUT(N__11789),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11791),
            .PADOUT(N__11790),
            .PADIN(N__11789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11782),
            .DIN(N__11781),
            .DOUT(N__11780),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11782),
            .PADOUT(N__11781),
            .PADIN(N__11780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11773),
            .DIN(N__11772),
            .DOUT(N__11771),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11773),
            .PADOUT(N__11772),
            .PADIN(N__11771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7566),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11764),
            .DIN(N__11763),
            .DOUT(N__11762),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11764),
            .PADOUT(N__11763),
            .PADIN(N__11762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11755),
            .DIN(N__11754),
            .DOUT(N__11753),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11755),
            .PADOUT(N__11754),
            .PADIN(N__11753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8569),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11746),
            .DIN(N__11745),
            .DOUT(N__11744),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11746),
            .PADOUT(N__11745),
            .PADIN(N__11744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8952),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11737),
            .DIN(N__11736),
            .DOUT(N__11735),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11737),
            .PADOUT(N__11736),
            .PADIN(N__11735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11728),
            .DIN(N__11727),
            .DOUT(N__11726),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11728),
            .PADOUT(N__11727),
            .PADIN(N__11726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5805),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11719),
            .DIN(N__11718),
            .DOUT(N__11717),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11719),
            .PADOUT(N__11718),
            .PADIN(N__11717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7935),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11710),
            .DIN(N__11709),
            .DOUT(N__11708),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11710),
            .PADOUT(N__11709),
            .PADIN(N__11708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4718),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11701),
            .DIN(N__11700),
            .DOUT(N__11699),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11701),
            .PADOUT(N__11700),
            .PADIN(N__11699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11692),
            .DIN(N__11691),
            .DOUT(N__11690),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11692),
            .PADOUT(N__11691),
            .PADIN(N__11690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11683),
            .DIN(N__11682),
            .DOUT(N__11681),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11683),
            .PADOUT(N__11682),
            .PADIN(N__11681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7239),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11674),
            .DIN(N__11673),
            .DOUT(N__11672),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11674),
            .PADOUT(N__11673),
            .PADIN(N__11672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7713),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11665),
            .DIN(N__11664),
            .DOUT(N__11663),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11665),
            .PADOUT(N__11664),
            .PADIN(N__11663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4209),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11656),
            .DIN(N__11655),
            .DOUT(N__11654),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11656),
            .PADOUT(N__11655),
            .PADIN(N__11654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11647),
            .DIN(N__11646),
            .DOUT(N__11645),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11647),
            .PADOUT(N__11646),
            .PADIN(N__11645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11638),
            .DIN(N__11637),
            .DOUT(N__11636),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11638),
            .PADOUT(N__11637),
            .PADIN(N__11636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11629),
            .DIN(N__11628),
            .DOUT(N__11627),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11629),
            .PADOUT(N__11628),
            .PADIN(N__11627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11620),
            .DIN(N__11619),
            .DOUT(N__11618),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11620),
            .PADOUT(N__11619),
            .PADIN(N__11618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11611),
            .DIN(N__11610),
            .DOUT(N__11609),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11611),
            .PADOUT(N__11610),
            .PADIN(N__11609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11602),
            .DIN(N__11601),
            .DOUT(N__11600),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11602),
            .PADOUT(N__11601),
            .PADIN(N__11600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11593),
            .DIN(N__11592),
            .DOUT(N__11591),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11593),
            .PADOUT(N__11592),
            .PADIN(N__11591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11584),
            .DIN(N__11583),
            .DOUT(N__11582),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11584),
            .PADOUT(N__11583),
            .PADIN(N__11582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5427),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11575),
            .DIN(N__11574),
            .DOUT(N__11573),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11575),
            .PADOUT(N__11574),
            .PADIN(N__11573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4158),
            .DIN0(),
            .DOUT0(N__4488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11566),
            .DIN(N__11565),
            .DOUT(N__11564),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11566),
            .PADOUT(N__11565),
            .PADIN(N__11564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7794),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11557),
            .DIN(N__11556),
            .DOUT(N__11555),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11557),
            .PADOUT(N__11556),
            .PADIN(N__11555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11548),
            .DIN(N__11547),
            .DOUT(N__11546),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11548),
            .PADOUT(N__11547),
            .PADIN(N__11546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11539),
            .DIN(N__11538),
            .DOUT(N__11537),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11539),
            .PADOUT(N__11538),
            .PADIN(N__11537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11530),
            .DIN(N__11529),
            .DOUT(N__11528),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11530),
            .PADOUT(N__11529),
            .PADIN(N__11528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11521),
            .DIN(N__11520),
            .DOUT(N__11519),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11521),
            .PADOUT(N__11520),
            .PADIN(N__11519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11512),
            .DIN(N__11511),
            .DOUT(N__11510),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11512),
            .PADOUT(N__11511),
            .PADIN(N__11510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11503),
            .DIN(N__11502),
            .DOUT(N__11501),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11503),
            .PADOUT(N__11502),
            .PADIN(N__11501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11494),
            .DIN(N__11493),
            .DOUT(N__11492),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11494),
            .PADOUT(N__11493),
            .PADIN(N__11492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4449),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11485),
            .DIN(N__11484),
            .DOUT(N__11483),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11485),
            .PADOUT(N__11484),
            .PADIN(N__11483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9792),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11476),
            .DIN(N__11475),
            .DOUT(N__11474),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11476),
            .PADOUT(N__11475),
            .PADIN(N__11474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8517),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11467),
            .DIN(N__11466),
            .DOUT(N__11465),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11467),
            .PADOUT(N__11466),
            .PADIN(N__11465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11458),
            .DIN(N__11457),
            .DOUT(N__11456),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11458),
            .PADOUT(N__11457),
            .PADIN(N__11456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11449),
            .DIN(N__11448),
            .DOUT(N__11447),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11449),
            .PADOUT(N__11448),
            .PADIN(N__11447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11440),
            .DIN(N__11439),
            .DOUT(N__11438),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11440),
            .PADOUT(N__11439),
            .PADIN(N__11438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9087),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11431),
            .DIN(N__11430),
            .DOUT(N__11429),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11431),
            .PADOUT(N__11430),
            .PADIN(N__11429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11422),
            .DIN(N__11421),
            .DOUT(N__11420),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11422),
            .PADOUT(N__11421),
            .PADIN(N__11420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11413),
            .DIN(N__11412),
            .DOUT(N__11411),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11413),
            .PADOUT(N__11412),
            .PADIN(N__11411),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4242),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11404),
            .DIN(N__11403),
            .DOUT(N__11402),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11404),
            .PADOUT(N__11403),
            .PADIN(N__11402),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9732),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11395),
            .DIN(N__11394),
            .DOUT(N__11393),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11395),
            .PADOUT(N__11394),
            .PADIN(N__11393),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8571),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11386),
            .DIN(N__11385),
            .DOUT(N__11384),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11386),
            .PADOUT(N__11385),
            .PADIN(N__11384),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11377),
            .DIN(N__11376),
            .DOUT(N__11375),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11377),
            .PADOUT(N__11376),
            .PADIN(N__11375),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8570),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11368),
            .DIN(N__11367),
            .DOUT(N__11366),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11368),
            .PADOUT(N__11367),
            .PADIN(N__11366),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4173),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2773 (
            .O(N__11349),
            .I(N__11346));
    LocalMux I__2772 (
            .O(N__11346),
            .I(N__11342));
    InMux I__2771 (
            .O(N__11345),
            .I(N__11338));
    Span4Mux_v I__2770 (
            .O(N__11342),
            .I(N__11335));
    InMux I__2769 (
            .O(N__11341),
            .I(N__11331));
    LocalMux I__2768 (
            .O(N__11338),
            .I(N__11328));
    Span4Mux_v I__2767 (
            .O(N__11335),
            .I(N__11325));
    InMux I__2766 (
            .O(N__11334),
            .I(N__11322));
    LocalMux I__2765 (
            .O(N__11331),
            .I(N__11319));
    Span12Mux_h I__2764 (
            .O(N__11328),
            .I(N__11316));
    Sp12to4 I__2763 (
            .O(N__11325),
            .I(N__11313));
    LocalMux I__2762 (
            .O(N__11322),
            .I(N__11310));
    Span12Mux_h I__2761 (
            .O(N__11319),
            .I(N__11307));
    Span12Mux_h I__2760 (
            .O(N__11316),
            .I(N__11304));
    Span12Mux_h I__2759 (
            .O(N__11313),
            .I(N__11299));
    Span12Mux_v I__2758 (
            .O(N__11310),
            .I(N__11299));
    Span12Mux_v I__2757 (
            .O(N__11307),
            .I(N__11296));
    Span12Mux_v I__2756 (
            .O(N__11304),
            .I(N__11291));
    Span12Mux_h I__2755 (
            .O(N__11299),
            .I(N__11291));
    Odrv12 I__2754 (
            .O(N__11296),
            .I(RnW_c));
    Odrv12 I__2753 (
            .O(N__11291),
            .I(RnW_c));
    InMux I__2752 (
            .O(N__11286),
            .I(N__11283));
    LocalMux I__2751 (
            .O(N__11283),
            .I(N__11280));
    Span4Mux_v I__2750 (
            .O(N__11280),
            .I(N__11276));
    InMux I__2749 (
            .O(N__11279),
            .I(N__11273));
    Span4Mux_v I__2748 (
            .O(N__11276),
            .I(N__11267));
    LocalMux I__2747 (
            .O(N__11273),
            .I(N__11267));
    InMux I__2746 (
            .O(N__11272),
            .I(N__11263));
    Span4Mux_h I__2745 (
            .O(N__11267),
            .I(N__11260));
    InMux I__2744 (
            .O(N__11266),
            .I(N__11257));
    LocalMux I__2743 (
            .O(N__11263),
            .I(N__11254));
    Span4Mux_v I__2742 (
            .O(N__11260),
            .I(N__11249));
    LocalMux I__2741 (
            .O(N__11257),
            .I(N__11249));
    Sp12to4 I__2740 (
            .O(N__11254),
            .I(N__11244));
    Span4Mux_v I__2739 (
            .O(N__11249),
            .I(N__11241));
    InMux I__2738 (
            .O(N__11248),
            .I(N__11236));
    InMux I__2737 (
            .O(N__11247),
            .I(N__11236));
    Span12Mux_v I__2736 (
            .O(N__11244),
            .I(N__11233));
    Sp12to4 I__2735 (
            .O(N__11241),
            .I(N__11230));
    LocalMux I__2734 (
            .O(N__11236),
            .I(N__11227));
    Span12Mux_h I__2733 (
            .O(N__11233),
            .I(N__11224));
    Span12Mux_h I__2732 (
            .O(N__11230),
            .I(N__11221));
    Span4Mux_v I__2731 (
            .O(N__11227),
            .I(N__11218));
    Odrv12 I__2730 (
            .O(N__11224),
            .I(CASUn_c));
    Odrv12 I__2729 (
            .O(N__11221),
            .I(CASUn_c));
    Odrv4 I__2728 (
            .O(N__11218),
            .I(CASUn_c));
    CascadeMux I__2727 (
            .O(N__11211),
            .I(N__11206));
    InMux I__2726 (
            .O(N__11210),
            .I(N__11202));
    InMux I__2725 (
            .O(N__11209),
            .I(N__11197));
    InMux I__2724 (
            .O(N__11206),
            .I(N__11197));
    InMux I__2723 (
            .O(N__11205),
            .I(N__11194));
    LocalMux I__2722 (
            .O(N__11202),
            .I(N__11191));
    LocalMux I__2721 (
            .O(N__11197),
            .I(N__11187));
    LocalMux I__2720 (
            .O(N__11194),
            .I(N__11184));
    Span4Mux_v I__2719 (
            .O(N__11191),
            .I(N__11181));
    CascadeMux I__2718 (
            .O(N__11190),
            .I(N__11177));
    Sp12to4 I__2717 (
            .O(N__11187),
            .I(N__11172));
    Sp12to4 I__2716 (
            .O(N__11184),
            .I(N__11172));
    Sp12to4 I__2715 (
            .O(N__11181),
            .I(N__11169));
    InMux I__2714 (
            .O(N__11180),
            .I(N__11164));
    InMux I__2713 (
            .O(N__11177),
            .I(N__11164));
    Span12Mux_v I__2712 (
            .O(N__11172),
            .I(N__11161));
    Span12Mux_h I__2711 (
            .O(N__11169),
            .I(N__11156));
    LocalMux I__2710 (
            .O(N__11164),
            .I(N__11156));
    Span12Mux_h I__2709 (
            .O(N__11161),
            .I(N__11151));
    Span12Mux_v I__2708 (
            .O(N__11156),
            .I(N__11151));
    Odrv12 I__2707 (
            .O(N__11151),
            .I(CASLn_c));
    InMux I__2706 (
            .O(N__11148),
            .I(N__11144));
    InMux I__2705 (
            .O(N__11147),
            .I(N__11141));
    LocalMux I__2704 (
            .O(N__11144),
            .I(N__11138));
    LocalMux I__2703 (
            .O(N__11141),
            .I(N__11133));
    Span4Mux_v I__2702 (
            .O(N__11138),
            .I(N__11129));
    InMux I__2701 (
            .O(N__11137),
            .I(N__11124));
    InMux I__2700 (
            .O(N__11136),
            .I(N__11124));
    Span4Mux_h I__2699 (
            .O(N__11133),
            .I(N__11120));
    InMux I__2698 (
            .O(N__11132),
            .I(N__11117));
    Span4Mux_v I__2697 (
            .O(N__11129),
            .I(N__11112));
    LocalMux I__2696 (
            .O(N__11124),
            .I(N__11112));
    InMux I__2695 (
            .O(N__11123),
            .I(N__11109));
    Sp12to4 I__2694 (
            .O(N__11120),
            .I(N__11106));
    LocalMux I__2693 (
            .O(N__11117),
            .I(N__11101));
    Span4Mux_v I__2692 (
            .O(N__11112),
            .I(N__11101));
    LocalMux I__2691 (
            .O(N__11109),
            .I(N__11097));
    Span12Mux_v I__2690 (
            .O(N__11106),
            .I(N__11089));
    Sp12to4 I__2689 (
            .O(N__11101),
            .I(N__11089));
    InMux I__2688 (
            .O(N__11100),
            .I(N__11086));
    Span4Mux_v I__2687 (
            .O(N__11097),
            .I(N__11083));
    InMux I__2686 (
            .O(N__11096),
            .I(N__11080));
    InMux I__2685 (
            .O(N__11095),
            .I(N__11075));
    InMux I__2684 (
            .O(N__11094),
            .I(N__11075));
    Odrv12 I__2683 (
            .O(N__11089),
            .I(WRITE_CYCLEm));
    LocalMux I__2682 (
            .O(N__11086),
            .I(WRITE_CYCLEm));
    Odrv4 I__2681 (
            .O(N__11083),
            .I(WRITE_CYCLEm));
    LocalMux I__2680 (
            .O(N__11080),
            .I(WRITE_CYCLEm));
    LocalMux I__2679 (
            .O(N__11075),
            .I(WRITE_CYCLEm));
    IoInMux I__2678 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__2677 (
            .O(N__11061),
            .I(N__11058));
    Span4Mux_s3_h I__2676 (
            .O(N__11058),
            .I(N__11055));
    Span4Mux_v I__2675 (
            .O(N__11055),
            .I(N__11052));
    Odrv4 I__2674 (
            .O(N__11052),
            .I(N_238));
    IoInMux I__2673 (
            .O(N__11049),
            .I(N__11046));
    LocalMux I__2672 (
            .O(N__11046),
            .I(N__11043));
    IoSpan4Mux I__2671 (
            .O(N__11043),
            .I(N__11040));
    Span4Mux_s3_v I__2670 (
            .O(N__11040),
            .I(N__11037));
    Sp12to4 I__2669 (
            .O(N__11037),
            .I(N__11034));
    Span12Mux_v I__2668 (
            .O(N__11034),
            .I(N__11031));
    Odrv12 I__2667 (
            .O(N__11031),
            .I(CMA_c_0));
    InMux I__2666 (
            .O(N__11028),
            .I(N__11024));
    InMux I__2665 (
            .O(N__11027),
            .I(N__11019));
    LocalMux I__2664 (
            .O(N__11024),
            .I(N__11016));
    InMux I__2663 (
            .O(N__11023),
            .I(N__11013));
    InMux I__2662 (
            .O(N__11022),
            .I(N__11010));
    LocalMux I__2661 (
            .O(N__11019),
            .I(N__11007));
    Span4Mux_v I__2660 (
            .O(N__11016),
            .I(N__11000));
    LocalMux I__2659 (
            .O(N__11013),
            .I(N__11000));
    LocalMux I__2658 (
            .O(N__11010),
            .I(N__11000));
    Span4Mux_h I__2657 (
            .O(N__11007),
            .I(N__10995));
    Span4Mux_h I__2656 (
            .O(N__11000),
            .I(N__10995));
    Sp12to4 I__2655 (
            .O(N__10995),
            .I(N__10992));
    Span12Mux_v I__2654 (
            .O(N__10992),
            .I(N__10989));
    Odrv12 I__2653 (
            .O(N__10989),
            .I(DRA_c_1));
    InMux I__2652 (
            .O(N__10986),
            .I(N__10983));
    LocalMux I__2651 (
            .O(N__10983),
            .I(N__10979));
    InMux I__2650 (
            .O(N__10982),
            .I(N__10976));
    Sp12to4 I__2649 (
            .O(N__10979),
            .I(N__10971));
    LocalMux I__2648 (
            .O(N__10976),
            .I(N__10971));
    Span12Mux_v I__2647 (
            .O(N__10971),
            .I(N__10968));
    Span12Mux_h I__2646 (
            .O(N__10968),
            .I(N__10965));
    Odrv12 I__2645 (
            .O(N__10965),
            .I(DRA_c_0));
    InMux I__2644 (
            .O(N__10962),
            .I(N__10959));
    LocalMux I__2643 (
            .O(N__10959),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2642 (
            .O(N__10956),
            .I(N__10953));
    LocalMux I__2641 (
            .O(N__10953),
            .I(N__10949));
    InMux I__2640 (
            .O(N__10952),
            .I(N__10946));
    Span4Mux_h I__2639 (
            .O(N__10949),
            .I(N__10943));
    LocalMux I__2638 (
            .O(N__10946),
            .I(N__10940));
    Span4Mux_h I__2637 (
            .O(N__10943),
            .I(N__10937));
    Span12Mux_v I__2636 (
            .O(N__10940),
            .I(N__10934));
    Odrv4 I__2635 (
            .O(N__10937),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    Odrv12 I__2634 (
            .O(N__10934),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2633 (
            .O(N__10929),
            .I(N__10926));
    LocalMux I__2632 (
            .O(N__10926),
            .I(N__10920));
    InMux I__2631 (
            .O(N__10925),
            .I(N__10915));
    InMux I__2630 (
            .O(N__10924),
            .I(N__10915));
    InMux I__2629 (
            .O(N__10923),
            .I(N__10912));
    Span4Mux_h I__2628 (
            .O(N__10920),
            .I(N__10907));
    LocalMux I__2627 (
            .O(N__10915),
            .I(N__10907));
    LocalMux I__2626 (
            .O(N__10912),
            .I(N__10904));
    Span4Mux_v I__2625 (
            .O(N__10907),
            .I(N__10901));
    Span12Mux_v I__2624 (
            .O(N__10904),
            .I(N__10898));
    Sp12to4 I__2623 (
            .O(N__10901),
            .I(N__10895));
    Span12Mux_h I__2622 (
            .O(N__10898),
            .I(N__10892));
    Odrv12 I__2621 (
            .O(N__10895),
            .I(DRA_c_5));
    Odrv12 I__2620 (
            .O(N__10892),
            .I(DRA_c_5));
    InMux I__2619 (
            .O(N__10887),
            .I(N__10884));
    LocalMux I__2618 (
            .O(N__10884),
            .I(N__10881));
    Odrv4 I__2617 (
            .O(N__10881),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2616 (
            .O(N__10878),
            .I(N__10873));
    InMux I__2615 (
            .O(N__10877),
            .I(N__10870));
    InMux I__2614 (
            .O(N__10876),
            .I(N__10867));
    LocalMux I__2613 (
            .O(N__10873),
            .I(N__10862));
    LocalMux I__2612 (
            .O(N__10870),
            .I(N__10859));
    LocalMux I__2611 (
            .O(N__10867),
            .I(N__10856));
    InMux I__2610 (
            .O(N__10866),
            .I(N__10851));
    InMux I__2609 (
            .O(N__10865),
            .I(N__10851));
    Span4Mux_h I__2608 (
            .O(N__10862),
            .I(N__10845));
    Span4Mux_h I__2607 (
            .O(N__10859),
            .I(N__10845));
    Span4Mux_h I__2606 (
            .O(N__10856),
            .I(N__10842));
    LocalMux I__2605 (
            .O(N__10851),
            .I(N__10839));
    InMux I__2604 (
            .O(N__10850),
            .I(N__10836));
    Odrv4 I__2603 (
            .O(N__10845),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    Odrv4 I__2602 (
            .O(N__10842),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    Odrv12 I__2601 (
            .O(N__10839),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__2600 (
            .O(N__10836),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    CascadeMux I__2599 (
            .O(N__10827),
            .I(N__10822));
    CascadeMux I__2598 (
            .O(N__10826),
            .I(N__10816));
    CascadeMux I__2597 (
            .O(N__10825),
            .I(N__10813));
    InMux I__2596 (
            .O(N__10822),
            .I(N__10810));
    CascadeMux I__2595 (
            .O(N__10821),
            .I(N__10807));
    CascadeMux I__2594 (
            .O(N__10820),
            .I(N__10804));
    CascadeMux I__2593 (
            .O(N__10819),
            .I(N__10799));
    InMux I__2592 (
            .O(N__10816),
            .I(N__10795));
    InMux I__2591 (
            .O(N__10813),
            .I(N__10792));
    LocalMux I__2590 (
            .O(N__10810),
            .I(N__10789));
    InMux I__2589 (
            .O(N__10807),
            .I(N__10784));
    InMux I__2588 (
            .O(N__10804),
            .I(N__10784));
    InMux I__2587 (
            .O(N__10803),
            .I(N__10781));
    InMux I__2586 (
            .O(N__10802),
            .I(N__10778));
    InMux I__2585 (
            .O(N__10799),
            .I(N__10775));
    CascadeMux I__2584 (
            .O(N__10798),
            .I(N__10772));
    LocalMux I__2583 (
            .O(N__10795),
            .I(N__10769));
    LocalMux I__2582 (
            .O(N__10792),
            .I(N__10762));
    Span4Mux_h I__2581 (
            .O(N__10789),
            .I(N__10762));
    LocalMux I__2580 (
            .O(N__10784),
            .I(N__10762));
    LocalMux I__2579 (
            .O(N__10781),
            .I(N__10755));
    LocalMux I__2578 (
            .O(N__10778),
            .I(N__10755));
    LocalMux I__2577 (
            .O(N__10775),
            .I(N__10755));
    InMux I__2576 (
            .O(N__10772),
            .I(N__10752));
    Span4Mux_v I__2575 (
            .O(N__10769),
            .I(N__10747));
    Span4Mux_v I__2574 (
            .O(N__10762),
            .I(N__10747));
    Span4Mux_h I__2573 (
            .O(N__10755),
            .I(N__10744));
    LocalMux I__2572 (
            .O(N__10752),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2571 (
            .O(N__10747),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2570 (
            .O(N__10744),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__2569 (
            .O(N__10737),
            .I(N__10734));
    LocalMux I__2568 (
            .O(N__10734),
            .I(N__10731));
    Odrv4 I__2567 (
            .O(N__10731),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__2566 (
            .O(N__10728),
            .I(N__10725));
    LocalMux I__2565 (
            .O(N__10725),
            .I(N__10722));
    Span4Mux_s0_h I__2564 (
            .O(N__10722),
            .I(N__10719));
    Sp12to4 I__2563 (
            .O(N__10719),
            .I(N__10716));
    Span12Mux_s6_v I__2562 (
            .O(N__10716),
            .I(N__10713));
    Span12Mux_h I__2561 (
            .O(N__10713),
            .I(N__10710));
    Odrv12 I__2560 (
            .O(N__10710),
            .I(CMA_c_3));
    InMux I__2559 (
            .O(N__10707),
            .I(N__10704));
    LocalMux I__2558 (
            .O(N__10704),
            .I(N__10663));
    ClkMux I__2557 (
            .O(N__10703),
            .I(N__10569));
    ClkMux I__2556 (
            .O(N__10702),
            .I(N__10569));
    ClkMux I__2555 (
            .O(N__10701),
            .I(N__10569));
    ClkMux I__2554 (
            .O(N__10700),
            .I(N__10569));
    ClkMux I__2553 (
            .O(N__10699),
            .I(N__10569));
    ClkMux I__2552 (
            .O(N__10698),
            .I(N__10569));
    ClkMux I__2551 (
            .O(N__10697),
            .I(N__10569));
    ClkMux I__2550 (
            .O(N__10696),
            .I(N__10569));
    ClkMux I__2549 (
            .O(N__10695),
            .I(N__10569));
    ClkMux I__2548 (
            .O(N__10694),
            .I(N__10569));
    ClkMux I__2547 (
            .O(N__10693),
            .I(N__10569));
    ClkMux I__2546 (
            .O(N__10692),
            .I(N__10569));
    ClkMux I__2545 (
            .O(N__10691),
            .I(N__10569));
    ClkMux I__2544 (
            .O(N__10690),
            .I(N__10569));
    ClkMux I__2543 (
            .O(N__10689),
            .I(N__10569));
    ClkMux I__2542 (
            .O(N__10688),
            .I(N__10569));
    ClkMux I__2541 (
            .O(N__10687),
            .I(N__10569));
    ClkMux I__2540 (
            .O(N__10686),
            .I(N__10569));
    ClkMux I__2539 (
            .O(N__10685),
            .I(N__10569));
    ClkMux I__2538 (
            .O(N__10684),
            .I(N__10569));
    ClkMux I__2537 (
            .O(N__10683),
            .I(N__10569));
    ClkMux I__2536 (
            .O(N__10682),
            .I(N__10569));
    ClkMux I__2535 (
            .O(N__10681),
            .I(N__10569));
    ClkMux I__2534 (
            .O(N__10680),
            .I(N__10569));
    ClkMux I__2533 (
            .O(N__10679),
            .I(N__10569));
    ClkMux I__2532 (
            .O(N__10678),
            .I(N__10569));
    ClkMux I__2531 (
            .O(N__10677),
            .I(N__10569));
    ClkMux I__2530 (
            .O(N__10676),
            .I(N__10569));
    ClkMux I__2529 (
            .O(N__10675),
            .I(N__10569));
    ClkMux I__2528 (
            .O(N__10674),
            .I(N__10569));
    ClkMux I__2527 (
            .O(N__10673),
            .I(N__10569));
    ClkMux I__2526 (
            .O(N__10672),
            .I(N__10569));
    ClkMux I__2525 (
            .O(N__10671),
            .I(N__10569));
    ClkMux I__2524 (
            .O(N__10670),
            .I(N__10569));
    ClkMux I__2523 (
            .O(N__10669),
            .I(N__10569));
    ClkMux I__2522 (
            .O(N__10668),
            .I(N__10569));
    ClkMux I__2521 (
            .O(N__10667),
            .I(N__10569));
    ClkMux I__2520 (
            .O(N__10666),
            .I(N__10569));
    Glb2LocalMux I__2519 (
            .O(N__10663),
            .I(N__10569));
    ClkMux I__2518 (
            .O(N__10662),
            .I(N__10569));
    ClkMux I__2517 (
            .O(N__10661),
            .I(N__10569));
    ClkMux I__2516 (
            .O(N__10660),
            .I(N__10569));
    ClkMux I__2515 (
            .O(N__10659),
            .I(N__10569));
    ClkMux I__2514 (
            .O(N__10658),
            .I(N__10569));
    GlobalMux I__2513 (
            .O(N__10569),
            .I(CLK80_PLL));
    CEMux I__2512 (
            .O(N__10566),
            .I(N__10562));
    CEMux I__2511 (
            .O(N__10565),
            .I(N__10557));
    LocalMux I__2510 (
            .O(N__10562),
            .I(N__10551));
    CEMux I__2509 (
            .O(N__10561),
            .I(N__10548));
    CEMux I__2508 (
            .O(N__10560),
            .I(N__10544));
    LocalMux I__2507 (
            .O(N__10557),
            .I(N__10540));
    CEMux I__2506 (
            .O(N__10556),
            .I(N__10537));
    CEMux I__2505 (
            .O(N__10555),
            .I(N__10534));
    CEMux I__2504 (
            .O(N__10554),
            .I(N__10531));
    Span4Mux_v I__2503 (
            .O(N__10551),
            .I(N__10526));
    LocalMux I__2502 (
            .O(N__10548),
            .I(N__10526));
    CEMux I__2501 (
            .O(N__10547),
            .I(N__10523));
    LocalMux I__2500 (
            .O(N__10544),
            .I(N__10520));
    CEMux I__2499 (
            .O(N__10543),
            .I(N__10517));
    Span4Mux_h I__2498 (
            .O(N__10540),
            .I(N__10512));
    LocalMux I__2497 (
            .O(N__10537),
            .I(N__10512));
    LocalMux I__2496 (
            .O(N__10534),
            .I(N__10509));
    LocalMux I__2495 (
            .O(N__10531),
            .I(N__10506));
    Span4Mux_v I__2494 (
            .O(N__10526),
            .I(N__10503));
    LocalMux I__2493 (
            .O(N__10523),
            .I(N__10500));
    Span4Mux_h I__2492 (
            .O(N__10520),
            .I(N__10495));
    LocalMux I__2491 (
            .O(N__10517),
            .I(N__10495));
    Span4Mux_h I__2490 (
            .O(N__10512),
            .I(N__10492));
    Span4Mux_v I__2489 (
            .O(N__10509),
            .I(N__10489));
    Span4Mux_h I__2488 (
            .O(N__10506),
            .I(N__10486));
    Span4Mux_h I__2487 (
            .O(N__10503),
            .I(N__10483));
    Span4Mux_h I__2486 (
            .O(N__10500),
            .I(N__10480));
    Span4Mux_v I__2485 (
            .O(N__10495),
            .I(N__10477));
    Odrv4 I__2484 (
            .O(N__10492),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2483 (
            .O(N__10489),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2482 (
            .O(N__10486),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2481 (
            .O(N__10483),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2480 (
            .O(N__10480),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2479 (
            .O(N__10477),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2478 (
            .O(N__10464),
            .I(N__10460));
    InMux I__2477 (
            .O(N__10463),
            .I(N__10457));
    LocalMux I__2476 (
            .O(N__10460),
            .I(N__10450));
    LocalMux I__2475 (
            .O(N__10457),
            .I(N__10450));
    InMux I__2474 (
            .O(N__10456),
            .I(N__10447));
    InMux I__2473 (
            .O(N__10455),
            .I(N__10444));
    Span4Mux_v I__2472 (
            .O(N__10450),
            .I(N__10441));
    LocalMux I__2471 (
            .O(N__10447),
            .I(N__10436));
    LocalMux I__2470 (
            .O(N__10444),
            .I(N__10436));
    Sp12to4 I__2469 (
            .O(N__10441),
            .I(N__10433));
    Span4Mux_v I__2468 (
            .O(N__10436),
            .I(N__10430));
    Span12Mux_h I__2467 (
            .O(N__10433),
            .I(N__10427));
    Sp12to4 I__2466 (
            .O(N__10430),
            .I(N__10424));
    Odrv12 I__2465 (
            .O(N__10427),
            .I(DRA_c_6));
    Odrv12 I__2464 (
            .O(N__10424),
            .I(DRA_c_6));
    InMux I__2463 (
            .O(N__10419),
            .I(N__10414));
    InMux I__2462 (
            .O(N__10418),
            .I(N__10410));
    InMux I__2461 (
            .O(N__10417),
            .I(N__10407));
    LocalMux I__2460 (
            .O(N__10414),
            .I(N__10404));
    InMux I__2459 (
            .O(N__10413),
            .I(N__10401));
    LocalMux I__2458 (
            .O(N__10410),
            .I(N__10396));
    LocalMux I__2457 (
            .O(N__10407),
            .I(N__10396));
    Span12Mux_v I__2456 (
            .O(N__10404),
            .I(N__10391));
    LocalMux I__2455 (
            .O(N__10401),
            .I(N__10391));
    Span12Mux_h I__2454 (
            .O(N__10396),
            .I(N__10388));
    Span12Mux_h I__2453 (
            .O(N__10391),
            .I(N__10385));
    Odrv12 I__2452 (
            .O(N__10388),
            .I(DRA_c_7));
    Odrv12 I__2451 (
            .O(N__10385),
            .I(DRA_c_7));
    InMux I__2450 (
            .O(N__10380),
            .I(N__10377));
    LocalMux I__2449 (
            .O(N__10377),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2448 (
            .O(N__10374),
            .I(N__10369));
    InMux I__2447 (
            .O(N__10373),
            .I(N__10366));
    InMux I__2446 (
            .O(N__10372),
            .I(N__10363));
    LocalMux I__2445 (
            .O(N__10369),
            .I(N__10357));
    LocalMux I__2444 (
            .O(N__10366),
            .I(N__10357));
    LocalMux I__2443 (
            .O(N__10363),
            .I(N__10354));
    InMux I__2442 (
            .O(N__10362),
            .I(N__10351));
    Span4Mux_v I__2441 (
            .O(N__10357),
            .I(N__10348));
    Span4Mux_h I__2440 (
            .O(N__10354),
            .I(N__10343));
    LocalMux I__2439 (
            .O(N__10351),
            .I(N__10343));
    Sp12to4 I__2438 (
            .O(N__10348),
            .I(N__10340));
    Span4Mux_v I__2437 (
            .O(N__10343),
            .I(N__10337));
    Span12Mux_h I__2436 (
            .O(N__10340),
            .I(N__10334));
    Sp12to4 I__2435 (
            .O(N__10337),
            .I(N__10331));
    Odrv12 I__2434 (
            .O(N__10334),
            .I(DRA_c_3));
    Odrv12 I__2433 (
            .O(N__10331),
            .I(DRA_c_3));
    InMux I__2432 (
            .O(N__10326),
            .I(N__10322));
    InMux I__2431 (
            .O(N__10325),
            .I(N__10319));
    LocalMux I__2430 (
            .O(N__10322),
            .I(N__10316));
    LocalMux I__2429 (
            .O(N__10319),
            .I(N__10312));
    Span4Mux_v I__2428 (
            .O(N__10316),
            .I(N__10304));
    InMux I__2427 (
            .O(N__10315),
            .I(N__10301));
    Span4Mux_v I__2426 (
            .O(N__10312),
            .I(N__10293));
    InMux I__2425 (
            .O(N__10311),
            .I(N__10290));
    InMux I__2424 (
            .O(N__10310),
            .I(N__10284));
    InMux I__2423 (
            .O(N__10309),
            .I(N__10281));
    InMux I__2422 (
            .O(N__10308),
            .I(N__10278));
    InMux I__2421 (
            .O(N__10307),
            .I(N__10275));
    Span4Mux_h I__2420 (
            .O(N__10304),
            .I(N__10270));
    LocalMux I__2419 (
            .O(N__10301),
            .I(N__10270));
    InMux I__2418 (
            .O(N__10300),
            .I(N__10267));
    InMux I__2417 (
            .O(N__10299),
            .I(N__10264));
    InMux I__2416 (
            .O(N__10298),
            .I(N__10261));
    InMux I__2415 (
            .O(N__10297),
            .I(N__10258));
    InMux I__2414 (
            .O(N__10296),
            .I(N__10255));
    Span4Mux_h I__2413 (
            .O(N__10293),
            .I(N__10247));
    LocalMux I__2412 (
            .O(N__10290),
            .I(N__10244));
    InMux I__2411 (
            .O(N__10289),
            .I(N__10241));
    InMux I__2410 (
            .O(N__10288),
            .I(N__10236));
    InMux I__2409 (
            .O(N__10287),
            .I(N__10236));
    LocalMux I__2408 (
            .O(N__10284),
            .I(N__10227));
    LocalMux I__2407 (
            .O(N__10281),
            .I(N__10227));
    LocalMux I__2406 (
            .O(N__10278),
            .I(N__10227));
    LocalMux I__2405 (
            .O(N__10275),
            .I(N__10227));
    Span4Mux_v I__2404 (
            .O(N__10270),
            .I(N__10222));
    LocalMux I__2403 (
            .O(N__10267),
            .I(N__10222));
    LocalMux I__2402 (
            .O(N__10264),
            .I(N__10215));
    LocalMux I__2401 (
            .O(N__10261),
            .I(N__10215));
    LocalMux I__2400 (
            .O(N__10258),
            .I(N__10215));
    LocalMux I__2399 (
            .O(N__10255),
            .I(N__10212));
    InMux I__2398 (
            .O(N__10254),
            .I(N__10209));
    InMux I__2397 (
            .O(N__10253),
            .I(N__10204));
    InMux I__2396 (
            .O(N__10252),
            .I(N__10204));
    InMux I__2395 (
            .O(N__10251),
            .I(N__10201));
    InMux I__2394 (
            .O(N__10250),
            .I(N__10198));
    Span4Mux_h I__2393 (
            .O(N__10247),
            .I(N__10187));
    Span4Mux_v I__2392 (
            .O(N__10244),
            .I(N__10187));
    LocalMux I__2391 (
            .O(N__10241),
            .I(N__10187));
    LocalMux I__2390 (
            .O(N__10236),
            .I(N__10187));
    Span4Mux_v I__2389 (
            .O(N__10227),
            .I(N__10187));
    Span4Mux_h I__2388 (
            .O(N__10222),
            .I(N__10180));
    Span4Mux_v I__2387 (
            .O(N__10215),
            .I(N__10180));
    Span4Mux_v I__2386 (
            .O(N__10212),
            .I(N__10180));
    LocalMux I__2385 (
            .O(N__10209),
            .I(N__10175));
    LocalMux I__2384 (
            .O(N__10204),
            .I(N__10175));
    LocalMux I__2383 (
            .O(N__10201),
            .I(N__10166));
    LocalMux I__2382 (
            .O(N__10198),
            .I(N__10166));
    Sp12to4 I__2381 (
            .O(N__10187),
            .I(N__10166));
    Sp12to4 I__2380 (
            .O(N__10180),
            .I(N__10166));
    Span12Mux_v I__2379 (
            .O(N__10175),
            .I(N__10163));
    Span12Mux_h I__2378 (
            .O(N__10166),
            .I(N__10160));
    Span12Mux_h I__2377 (
            .O(N__10163),
            .I(N__10157));
    Span12Mux_v I__2376 (
            .O(N__10160),
            .I(N__10154));
    Odrv12 I__2375 (
            .O(N__10157),
            .I(AGNUS_REV_c));
    Odrv12 I__2374 (
            .O(N__10154),
            .I(AGNUS_REV_c));
    InMux I__2373 (
            .O(N__10149),
            .I(N__10143));
    InMux I__2372 (
            .O(N__10148),
            .I(N__10140));
    InMux I__2371 (
            .O(N__10147),
            .I(N__10137));
    InMux I__2370 (
            .O(N__10146),
            .I(N__10134));
    LocalMux I__2369 (
            .O(N__10143),
            .I(N__10129));
    LocalMux I__2368 (
            .O(N__10140),
            .I(N__10129));
    LocalMux I__2367 (
            .O(N__10137),
            .I(N__10126));
    LocalMux I__2366 (
            .O(N__10134),
            .I(N__10123));
    Span4Mux_v I__2365 (
            .O(N__10129),
            .I(N__10120));
    Span4Mux_v I__2364 (
            .O(N__10126),
            .I(N__10117));
    Span12Mux_v I__2363 (
            .O(N__10123),
            .I(N__10110));
    Sp12to4 I__2362 (
            .O(N__10120),
            .I(N__10110));
    Sp12to4 I__2361 (
            .O(N__10117),
            .I(N__10110));
    Span12Mux_h I__2360 (
            .O(N__10110),
            .I(N__10107));
    Odrv12 I__2359 (
            .O(N__10107),
            .I(DRA_c_4));
    InMux I__2358 (
            .O(N__10104),
            .I(N__10101));
    LocalMux I__2357 (
            .O(N__10101),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    ClkMux I__2356 (
            .O(N__10098),
            .I(N__10074));
    ClkMux I__2355 (
            .O(N__10097),
            .I(N__10074));
    ClkMux I__2354 (
            .O(N__10096),
            .I(N__10074));
    ClkMux I__2353 (
            .O(N__10095),
            .I(N__10074));
    ClkMux I__2352 (
            .O(N__10094),
            .I(N__10074));
    ClkMux I__2351 (
            .O(N__10093),
            .I(N__10074));
    ClkMux I__2350 (
            .O(N__10092),
            .I(N__10074));
    ClkMux I__2349 (
            .O(N__10091),
            .I(N__10074));
    GlobalMux I__2348 (
            .O(N__10074),
            .I(N__10071));
    gio2CtrlBuf I__2347 (
            .O(N__10071),
            .I(C3_c_g));
    CEMux I__2346 (
            .O(N__10068),
            .I(N__10023));
    CEMux I__2345 (
            .O(N__10067),
            .I(N__10023));
    CEMux I__2344 (
            .O(N__10066),
            .I(N__10023));
    CEMux I__2343 (
            .O(N__10065),
            .I(N__10023));
    CEMux I__2342 (
            .O(N__10064),
            .I(N__10023));
    CEMux I__2341 (
            .O(N__10063),
            .I(N__10023));
    CEMux I__2340 (
            .O(N__10062),
            .I(N__10023));
    CEMux I__2339 (
            .O(N__10061),
            .I(N__10023));
    CEMux I__2338 (
            .O(N__10060),
            .I(N__10023));
    CEMux I__2337 (
            .O(N__10059),
            .I(N__10023));
    CEMux I__2336 (
            .O(N__10058),
            .I(N__10023));
    CEMux I__2335 (
            .O(N__10057),
            .I(N__10023));
    CEMux I__2334 (
            .O(N__10056),
            .I(N__10023));
    CEMux I__2333 (
            .O(N__10055),
            .I(N__10023));
    CEMux I__2332 (
            .O(N__10054),
            .I(N__10023));
    GlobalMux I__2331 (
            .O(N__10023),
            .I(N__10020));
    gio2CtrlBuf I__2330 (
            .O(N__10020),
            .I(DBRn_c_i_0_g));
    InMux I__2329 (
            .O(N__10017),
            .I(N__10010));
    InMux I__2328 (
            .O(N__10016),
            .I(N__10007));
    InMux I__2327 (
            .O(N__10015),
            .I(N__10004));
    InMux I__2326 (
            .O(N__10014),
            .I(N__10001));
    InMux I__2325 (
            .O(N__10013),
            .I(N__9998));
    LocalMux I__2324 (
            .O(N__10010),
            .I(N__9995));
    LocalMux I__2323 (
            .O(N__10007),
            .I(N__9975));
    LocalMux I__2322 (
            .O(N__10004),
            .I(N__9962));
    LocalMux I__2321 (
            .O(N__10001),
            .I(N__9955));
    LocalMux I__2320 (
            .O(N__9998),
            .I(N__9947));
    Glb2LocalMux I__2319 (
            .O(N__9995),
            .I(N__9849));
    SRMux I__2318 (
            .O(N__9994),
            .I(N__9849));
    SRMux I__2317 (
            .O(N__9993),
            .I(N__9849));
    SRMux I__2316 (
            .O(N__9992),
            .I(N__9849));
    SRMux I__2315 (
            .O(N__9991),
            .I(N__9849));
    SRMux I__2314 (
            .O(N__9990),
            .I(N__9849));
    SRMux I__2313 (
            .O(N__9989),
            .I(N__9849));
    SRMux I__2312 (
            .O(N__9988),
            .I(N__9849));
    SRMux I__2311 (
            .O(N__9987),
            .I(N__9849));
    SRMux I__2310 (
            .O(N__9986),
            .I(N__9849));
    SRMux I__2309 (
            .O(N__9985),
            .I(N__9849));
    SRMux I__2308 (
            .O(N__9984),
            .I(N__9849));
    SRMux I__2307 (
            .O(N__9983),
            .I(N__9849));
    SRMux I__2306 (
            .O(N__9982),
            .I(N__9849));
    SRMux I__2305 (
            .O(N__9981),
            .I(N__9849));
    SRMux I__2304 (
            .O(N__9980),
            .I(N__9849));
    SRMux I__2303 (
            .O(N__9979),
            .I(N__9849));
    SRMux I__2302 (
            .O(N__9978),
            .I(N__9849));
    Glb2LocalMux I__2301 (
            .O(N__9975),
            .I(N__9849));
    SRMux I__2300 (
            .O(N__9974),
            .I(N__9849));
    SRMux I__2299 (
            .O(N__9973),
            .I(N__9849));
    SRMux I__2298 (
            .O(N__9972),
            .I(N__9849));
    SRMux I__2297 (
            .O(N__9971),
            .I(N__9849));
    SRMux I__2296 (
            .O(N__9970),
            .I(N__9849));
    SRMux I__2295 (
            .O(N__9969),
            .I(N__9849));
    SRMux I__2294 (
            .O(N__9968),
            .I(N__9849));
    SRMux I__2293 (
            .O(N__9967),
            .I(N__9849));
    SRMux I__2292 (
            .O(N__9966),
            .I(N__9849));
    SRMux I__2291 (
            .O(N__9965),
            .I(N__9849));
    Glb2LocalMux I__2290 (
            .O(N__9962),
            .I(N__9849));
    SRMux I__2289 (
            .O(N__9961),
            .I(N__9849));
    SRMux I__2288 (
            .O(N__9960),
            .I(N__9849));
    SRMux I__2287 (
            .O(N__9959),
            .I(N__9849));
    SRMux I__2286 (
            .O(N__9958),
            .I(N__9849));
    Glb2LocalMux I__2285 (
            .O(N__9955),
            .I(N__9849));
    SRMux I__2284 (
            .O(N__9954),
            .I(N__9849));
    SRMux I__2283 (
            .O(N__9953),
            .I(N__9849));
    SRMux I__2282 (
            .O(N__9952),
            .I(N__9849));
    SRMux I__2281 (
            .O(N__9951),
            .I(N__9849));
    SRMux I__2280 (
            .O(N__9950),
            .I(N__9849));
    Glb2LocalMux I__2279 (
            .O(N__9947),
            .I(N__9849));
    SRMux I__2278 (
            .O(N__9946),
            .I(N__9849));
    SRMux I__2277 (
            .O(N__9945),
            .I(N__9849));
    SRMux I__2276 (
            .O(N__9944),
            .I(N__9849));
    SRMux I__2275 (
            .O(N__9943),
            .I(N__9849));
    SRMux I__2274 (
            .O(N__9942),
            .I(N__9849));
    GlobalMux I__2273 (
            .O(N__9849),
            .I(N__9846));
    gio2CtrlBuf I__2272 (
            .O(N__9846),
            .I(RESETn_c_i_g));
    InMux I__2271 (
            .O(N__9843),
            .I(N__9839));
    InMux I__2270 (
            .O(N__9842),
            .I(N__9836));
    LocalMux I__2269 (
            .O(N__9839),
            .I(N__9833));
    LocalMux I__2268 (
            .O(N__9836),
            .I(N__9830));
    Span12Mux_v I__2267 (
            .O(N__9833),
            .I(N__9826));
    Span4Mux_h I__2266 (
            .O(N__9830),
            .I(N__9823));
    CascadeMux I__2265 (
            .O(N__9829),
            .I(N__9820));
    Span12Mux_h I__2264 (
            .O(N__9826),
            .I(N__9817));
    Span4Mux_v I__2263 (
            .O(N__9823),
            .I(N__9814));
    InMux I__2262 (
            .O(N__9820),
            .I(N__9811));
    Odrv12 I__2261 (
            .O(N__9817),
            .I(REG_CYCLEm));
    Odrv4 I__2260 (
            .O(N__9814),
            .I(REG_CYCLEm));
    LocalMux I__2259 (
            .O(N__9811),
            .I(REG_CYCLEm));
    IoInMux I__2258 (
            .O(N__9804),
            .I(N__9801));
    LocalMux I__2257 (
            .O(N__9801),
            .I(N__9798));
    Span12Mux_s6_v I__2256 (
            .O(N__9798),
            .I(N__9795));
    Odrv12 I__2255 (
            .O(N__9795),
            .I(DRDENn_c));
    IoInMux I__2254 (
            .O(N__9792),
            .I(N__9789));
    LocalMux I__2253 (
            .O(N__9789),
            .I(N__9786));
    Span4Mux_s3_v I__2252 (
            .O(N__9786),
            .I(N__9783));
    Span4Mux_h I__2251 (
            .O(N__9783),
            .I(N__9780));
    Span4Mux_v I__2250 (
            .O(N__9780),
            .I(N__9777));
    Odrv4 I__2249 (
            .O(N__9777),
            .I(U712_BYTE_ENABLE_un1_UDSn_i));
    IoInMux I__2248 (
            .O(N__9774),
            .I(N__9771));
    LocalMux I__2247 (
            .O(N__9771),
            .I(N__9768));
    Span4Mux_s0_v I__2246 (
            .O(N__9768),
            .I(N__9765));
    Span4Mux_v I__2245 (
            .O(N__9765),
            .I(N__9762));
    Odrv4 I__2244 (
            .O(N__9762),
            .I(LLBEn_c));
    CascadeMux I__2243 (
            .O(N__9759),
            .I(N__9756));
    InMux I__2242 (
            .O(N__9756),
            .I(N__9752));
    InMux I__2241 (
            .O(N__9755),
            .I(N__9749));
    LocalMux I__2240 (
            .O(N__9752),
            .I(N__9744));
    LocalMux I__2239 (
            .O(N__9749),
            .I(N__9744));
    Span4Mux_v I__2238 (
            .O(N__9744),
            .I(N__9740));
    InMux I__2237 (
            .O(N__9743),
            .I(N__9737));
    Odrv4 I__2236 (
            .O(N__9740),
            .I(DS_ENm));
    LocalMux I__2235 (
            .O(N__9737),
            .I(DS_ENm));
    IoInMux I__2234 (
            .O(N__9732),
            .I(N__9729));
    LocalMux I__2233 (
            .O(N__9729),
            .I(N__9726));
    Span4Mux_s3_v I__2232 (
            .O(N__9726),
            .I(N__9723));
    Span4Mux_h I__2231 (
            .O(N__9723),
            .I(N__9720));
    Span4Mux_h I__2230 (
            .O(N__9720),
            .I(N__9717));
    Odrv4 I__2229 (
            .O(N__9717),
            .I(N_119));
    InMux I__2228 (
            .O(N__9714),
            .I(N__9709));
    InMux I__2227 (
            .O(N__9713),
            .I(N__9706));
    InMux I__2226 (
            .O(N__9712),
            .I(N__9703));
    LocalMux I__2225 (
            .O(N__9709),
            .I(N__9691));
    LocalMux I__2224 (
            .O(N__9706),
            .I(N__9691));
    LocalMux I__2223 (
            .O(N__9703),
            .I(N__9691));
    InMux I__2222 (
            .O(N__9702),
            .I(N__9688));
    InMux I__2221 (
            .O(N__9701),
            .I(N__9683));
    InMux I__2220 (
            .O(N__9700),
            .I(N__9683));
    InMux I__2219 (
            .O(N__9699),
            .I(N__9678));
    InMux I__2218 (
            .O(N__9698),
            .I(N__9678));
    Span4Mux_h I__2217 (
            .O(N__9691),
            .I(N__9673));
    LocalMux I__2216 (
            .O(N__9688),
            .I(N__9673));
    LocalMux I__2215 (
            .O(N__9683),
            .I(N__9668));
    LocalMux I__2214 (
            .O(N__9678),
            .I(N__9668));
    Span4Mux_v I__2213 (
            .O(N__9673),
            .I(N__9665));
    Span4Mux_v I__2212 (
            .O(N__9668),
            .I(N__9662));
    Sp12to4 I__2211 (
            .O(N__9665),
            .I(N__9657));
    Sp12to4 I__2210 (
            .O(N__9662),
            .I(N__9657));
    Span12Mux_h I__2209 (
            .O(N__9657),
            .I(N__9654));
    Odrv12 I__2208 (
            .O(N__9654),
            .I(A_c_1));
    CascadeMux I__2207 (
            .O(N__9651),
            .I(N__9643));
    CascadeMux I__2206 (
            .O(N__9650),
            .I(N__9638));
    InMux I__2205 (
            .O(N__9649),
            .I(N__9633));
    InMux I__2204 (
            .O(N__9648),
            .I(N__9633));
    InMux I__2203 (
            .O(N__9647),
            .I(N__9629));
    InMux I__2202 (
            .O(N__9646),
            .I(N__9624));
    InMux I__2201 (
            .O(N__9643),
            .I(N__9624));
    InMux I__2200 (
            .O(N__9642),
            .I(N__9621));
    InMux I__2199 (
            .O(N__9641),
            .I(N__9616));
    InMux I__2198 (
            .O(N__9638),
            .I(N__9616));
    LocalMux I__2197 (
            .O(N__9633),
            .I(N__9613));
    InMux I__2196 (
            .O(N__9632),
            .I(N__9610));
    LocalMux I__2195 (
            .O(N__9629),
            .I(N__9603));
    LocalMux I__2194 (
            .O(N__9624),
            .I(N__9603));
    LocalMux I__2193 (
            .O(N__9621),
            .I(N__9603));
    LocalMux I__2192 (
            .O(N__9616),
            .I(N__9600));
    Span4Mux_h I__2191 (
            .O(N__9613),
            .I(N__9597));
    LocalMux I__2190 (
            .O(N__9610),
            .I(N__9594));
    Span4Mux_v I__2189 (
            .O(N__9603),
            .I(N__9590));
    Span4Mux_v I__2188 (
            .O(N__9600),
            .I(N__9587));
    Span4Mux_v I__2187 (
            .O(N__9597),
            .I(N__9582));
    Span4Mux_v I__2186 (
            .O(N__9594),
            .I(N__9582));
    InMux I__2185 (
            .O(N__9593),
            .I(N__9579));
    Sp12to4 I__2184 (
            .O(N__9590),
            .I(N__9570));
    Sp12to4 I__2183 (
            .O(N__9587),
            .I(N__9570));
    Sp12to4 I__2182 (
            .O(N__9582),
            .I(N__9570));
    LocalMux I__2181 (
            .O(N__9579),
            .I(N__9570));
    Span12Mux_h I__2180 (
            .O(N__9570),
            .I(N__9567));
    Odrv12 I__2179 (
            .O(N__9567),
            .I(A_c_0));
    CascadeMux I__2178 (
            .O(N__9564),
            .I(N__9560));
    InMux I__2177 (
            .O(N__9563),
            .I(N__9552));
    InMux I__2176 (
            .O(N__9560),
            .I(N__9552));
    InMux I__2175 (
            .O(N__9559),
            .I(N__9547));
    InMux I__2174 (
            .O(N__9558),
            .I(N__9547));
    CascadeMux I__2173 (
            .O(N__9557),
            .I(N__9543));
    LocalMux I__2172 (
            .O(N__9552),
            .I(N__9539));
    LocalMux I__2171 (
            .O(N__9547),
            .I(N__9536));
    InMux I__2170 (
            .O(N__9546),
            .I(N__9529));
    InMux I__2169 (
            .O(N__9543),
            .I(N__9529));
    InMux I__2168 (
            .O(N__9542),
            .I(N__9529));
    Span4Mux_v I__2167 (
            .O(N__9539),
            .I(N__9525));
    Span4Mux_v I__2166 (
            .O(N__9536),
            .I(N__9522));
    LocalMux I__2165 (
            .O(N__9529),
            .I(N__9519));
    CascadeMux I__2164 (
            .O(N__9528),
            .I(N__9516));
    Span4Mux_v I__2163 (
            .O(N__9525),
            .I(N__9513));
    Span4Mux_v I__2162 (
            .O(N__9522),
            .I(N__9508));
    Span4Mux_h I__2161 (
            .O(N__9519),
            .I(N__9508));
    InMux I__2160 (
            .O(N__9516),
            .I(N__9505));
    Span4Mux_v I__2159 (
            .O(N__9513),
            .I(N__9502));
    Span4Mux_v I__2158 (
            .O(N__9508),
            .I(N__9499));
    LocalMux I__2157 (
            .O(N__9505),
            .I(N__9496));
    Sp12to4 I__2156 (
            .O(N__9502),
            .I(N__9489));
    Sp12to4 I__2155 (
            .O(N__9499),
            .I(N__9489));
    Span12Mux_v I__2154 (
            .O(N__9496),
            .I(N__9489));
    Span12Mux_h I__2153 (
            .O(N__9489),
            .I(N__9486));
    Odrv12 I__2152 (
            .O(N__9486),
            .I(SIZ_c_1));
    InMux I__2151 (
            .O(N__9483),
            .I(N__9476));
    InMux I__2150 (
            .O(N__9482),
            .I(N__9473));
    InMux I__2149 (
            .O(N__9481),
            .I(N__9466));
    InMux I__2148 (
            .O(N__9480),
            .I(N__9466));
    InMux I__2147 (
            .O(N__9479),
            .I(N__9466));
    LocalMux I__2146 (
            .O(N__9476),
            .I(N__9462));
    LocalMux I__2145 (
            .O(N__9473),
            .I(N__9459));
    LocalMux I__2144 (
            .O(N__9466),
            .I(N__9456));
    InMux I__2143 (
            .O(N__9465),
            .I(N__9453));
    Span4Mux_v I__2142 (
            .O(N__9462),
            .I(N__9450));
    Span4Mux_v I__2141 (
            .O(N__9459),
            .I(N__9447));
    Span4Mux_h I__2140 (
            .O(N__9456),
            .I(N__9442));
    LocalMux I__2139 (
            .O(N__9453),
            .I(N__9442));
    Span4Mux_v I__2138 (
            .O(N__9450),
            .I(N__9439));
    Span4Mux_v I__2137 (
            .O(N__9447),
            .I(N__9434));
    Span4Mux_h I__2136 (
            .O(N__9442),
            .I(N__9434));
    Span4Mux_v I__2135 (
            .O(N__9439),
            .I(N__9431));
    Span4Mux_v I__2134 (
            .O(N__9434),
            .I(N__9428));
    Span4Mux_h I__2133 (
            .O(N__9431),
            .I(N__9425));
    Span4Mux_h I__2132 (
            .O(N__9428),
            .I(N__9422));
    Sp12to4 I__2131 (
            .O(N__9425),
            .I(N__9417));
    Sp12to4 I__2130 (
            .O(N__9422),
            .I(N__9417));
    Odrv12 I__2129 (
            .O(N__9417),
            .I(SIZ_c_0));
    IoInMux I__2128 (
            .O(N__9414),
            .I(N__9411));
    LocalMux I__2127 (
            .O(N__9411),
            .I(N__9408));
    Span4Mux_s3_v I__2126 (
            .O(N__9408),
            .I(N__9405));
    Odrv4 I__2125 (
            .O(N__9405),
            .I(N_220_i));
    CascadeMux I__2124 (
            .O(N__9402),
            .I(N__9393));
    InMux I__2123 (
            .O(N__9401),
            .I(N__9389));
    InMux I__2122 (
            .O(N__9400),
            .I(N__9384));
    InMux I__2121 (
            .O(N__9399),
            .I(N__9384));
    InMux I__2120 (
            .O(N__9398),
            .I(N__9381));
    InMux I__2119 (
            .O(N__9397),
            .I(N__9374));
    InMux I__2118 (
            .O(N__9396),
            .I(N__9374));
    InMux I__2117 (
            .O(N__9393),
            .I(N__9371));
    InMux I__2116 (
            .O(N__9392),
            .I(N__9367));
    LocalMux I__2115 (
            .O(N__9389),
            .I(N__9364));
    LocalMux I__2114 (
            .O(N__9384),
            .I(N__9353));
    LocalMux I__2113 (
            .O(N__9381),
            .I(N__9350));
    CascadeMux I__2112 (
            .O(N__9380),
            .I(N__9347));
    CascadeMux I__2111 (
            .O(N__9379),
            .I(N__9344));
    LocalMux I__2110 (
            .O(N__9374),
            .I(N__9337));
    LocalMux I__2109 (
            .O(N__9371),
            .I(N__9337));
    InMux I__2108 (
            .O(N__9370),
            .I(N__9334));
    LocalMux I__2107 (
            .O(N__9367),
            .I(N__9327));
    Span4Mux_v I__2106 (
            .O(N__9364),
            .I(N__9327));
    InMux I__2105 (
            .O(N__9363),
            .I(N__9324));
    InMux I__2104 (
            .O(N__9362),
            .I(N__9321));
    InMux I__2103 (
            .O(N__9361),
            .I(N__9317));
    InMux I__2102 (
            .O(N__9360),
            .I(N__9310));
    InMux I__2101 (
            .O(N__9359),
            .I(N__9310));
    InMux I__2100 (
            .O(N__9358),
            .I(N__9310));
    InMux I__2099 (
            .O(N__9357),
            .I(N__9305));
    InMux I__2098 (
            .O(N__9356),
            .I(N__9305));
    Span4Mux_v I__2097 (
            .O(N__9353),
            .I(N__9300));
    Span4Mux_v I__2096 (
            .O(N__9350),
            .I(N__9300));
    InMux I__2095 (
            .O(N__9347),
            .I(N__9291));
    InMux I__2094 (
            .O(N__9344),
            .I(N__9291));
    InMux I__2093 (
            .O(N__9343),
            .I(N__9291));
    InMux I__2092 (
            .O(N__9342),
            .I(N__9291));
    Span4Mux_v I__2091 (
            .O(N__9337),
            .I(N__9288));
    LocalMux I__2090 (
            .O(N__9334),
            .I(N__9285));
    InMux I__2089 (
            .O(N__9333),
            .I(N__9280));
    InMux I__2088 (
            .O(N__9332),
            .I(N__9280));
    Span4Mux_h I__2087 (
            .O(N__9327),
            .I(N__9273));
    LocalMux I__2086 (
            .O(N__9324),
            .I(N__9273));
    LocalMux I__2085 (
            .O(N__9321),
            .I(N__9273));
    InMux I__2084 (
            .O(N__9320),
            .I(N__9270));
    LocalMux I__2083 (
            .O(N__9317),
            .I(N__9267));
    LocalMux I__2082 (
            .O(N__9310),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2081 (
            .O(N__9305),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2080 (
            .O(N__9300),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2079 (
            .O(N__9291),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2078 (
            .O(N__9288),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2077 (
            .O(N__9285),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2076 (
            .O(N__9280),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2075 (
            .O(N__9273),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2074 (
            .O(N__9270),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2073 (
            .O(N__9267),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__2072 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__2071 (
            .O(N__9243),
            .I(N__9240));
    Span4Mux_s2_v I__2070 (
            .O(N__9240),
            .I(N__9237));
    Span4Mux_v I__2069 (
            .O(N__9237),
            .I(N__9234));
    Span4Mux_v I__2068 (
            .O(N__9234),
            .I(N__9231));
    Span4Mux_h I__2067 (
            .O(N__9231),
            .I(N__9228));
    Odrv4 I__2066 (
            .O(N__9228),
            .I(CASn_c));
    InMux I__2065 (
            .O(N__9225),
            .I(N__9222));
    LocalMux I__2064 (
            .O(N__9222),
            .I(N__9219));
    Span12Mux_h I__2063 (
            .O(N__9219),
            .I(N__9216));
    Odrv12 I__2062 (
            .O(N__9216),
            .I(RAS0n_c));
    InMux I__2061 (
            .O(N__9213),
            .I(N__9209));
    InMux I__2060 (
            .O(N__9212),
            .I(N__9204));
    LocalMux I__2059 (
            .O(N__9209),
            .I(N__9201));
    InMux I__2058 (
            .O(N__9208),
            .I(N__9198));
    InMux I__2057 (
            .O(N__9207),
            .I(N__9195));
    LocalMux I__2056 (
            .O(N__9204),
            .I(N__9192));
    Span4Mux_h I__2055 (
            .O(N__9201),
            .I(N__9185));
    LocalMux I__2054 (
            .O(N__9198),
            .I(N__9185));
    LocalMux I__2053 (
            .O(N__9195),
            .I(N__9185));
    Span4Mux_h I__2052 (
            .O(N__9192),
            .I(N__9182));
    Span4Mux_h I__2051 (
            .O(N__9185),
            .I(N__9179));
    Sp12to4 I__2050 (
            .O(N__9182),
            .I(N__9176));
    Span4Mux_v I__2049 (
            .O(N__9179),
            .I(N__9173));
    Span12Mux_v I__2048 (
            .O(N__9176),
            .I(N__9170));
    Sp12to4 I__2047 (
            .O(N__9173),
            .I(N__9167));
    Span12Mux_h I__2046 (
            .O(N__9170),
            .I(N__9164));
    Span12Mux_v I__2045 (
            .O(N__9167),
            .I(N__9161));
    Odrv12 I__2044 (
            .O(N__9164),
            .I(DRA_c_9));
    Odrv12 I__2043 (
            .O(N__9161),
            .I(DRA_c_9));
    InMux I__2042 (
            .O(N__9156),
            .I(N__9153));
    LocalMux I__2041 (
            .O(N__9153),
            .I(N__9150));
    Span4Mux_v I__2040 (
            .O(N__9150),
            .I(N__9147));
    Odrv4 I__2039 (
            .O(N__9147),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2038 (
            .O(N__9144),
            .I(N__9141));
    LocalMux I__2037 (
            .O(N__9141),
            .I(N__9136));
    InMux I__2036 (
            .O(N__9140),
            .I(N__9133));
    InMux I__2035 (
            .O(N__9139),
            .I(N__9130));
    Span4Mux_v I__2034 (
            .O(N__9136),
            .I(N__9126));
    LocalMux I__2033 (
            .O(N__9133),
            .I(N__9123));
    LocalMux I__2032 (
            .O(N__9130),
            .I(N__9120));
    InMux I__2031 (
            .O(N__9129),
            .I(N__9117));
    Sp12to4 I__2030 (
            .O(N__9126),
            .I(N__9108));
    Span12Mux_v I__2029 (
            .O(N__9123),
            .I(N__9108));
    Span12Mux_v I__2028 (
            .O(N__9120),
            .I(N__9108));
    LocalMux I__2027 (
            .O(N__9117),
            .I(N__9108));
    Span12Mux_h I__2026 (
            .O(N__9108),
            .I(N__9105));
    Odrv12 I__2025 (
            .O(N__9105),
            .I(DRA_c_8));
    InMux I__2024 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__2023 (
            .O(N__9099),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2022 (
            .O(N__9096),
            .I(N__9093));
    LocalMux I__2021 (
            .O(N__9093),
            .I(N__9090));
    Odrv4 I__2020 (
            .O(N__9090),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__2019 (
            .O(N__9087),
            .I(N__9084));
    LocalMux I__2018 (
            .O(N__9084),
            .I(N__9081));
    Span12Mux_s5_h I__2017 (
            .O(N__9081),
            .I(N__9078));
    Span12Mux_v I__2016 (
            .O(N__9078),
            .I(N__9075));
    Odrv12 I__2015 (
            .O(N__9075),
            .I(CMA_c_6));
    InMux I__2014 (
            .O(N__9072),
            .I(N__9069));
    LocalMux I__2013 (
            .O(N__9069),
            .I(N__9066));
    Odrv12 I__2012 (
            .O(N__9066),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__2011 (
            .O(N__9063),
            .I(N__9060));
    LocalMux I__2010 (
            .O(N__9060),
            .I(N__9057));
    Span4Mux_s3_v I__2009 (
            .O(N__9057),
            .I(N__9054));
    Odrv4 I__2008 (
            .O(N__9054),
            .I(U712_BYTE_ENABLE_UUBE_i));
    CascadeMux I__2007 (
            .O(N__9051),
            .I(N__9047));
    InMux I__2006 (
            .O(N__9050),
            .I(N__9044));
    InMux I__2005 (
            .O(N__9047),
            .I(N__9041));
    LocalMux I__2004 (
            .O(N__9044),
            .I(N__9038));
    LocalMux I__2003 (
            .O(N__9041),
            .I(N__9034));
    Span4Mux_h I__2002 (
            .O(N__9038),
            .I(N__9031));
    CascadeMux I__2001 (
            .O(N__9037),
            .I(N__9026));
    Span4Mux_v I__2000 (
            .O(N__9034),
            .I(N__9023));
    Span4Mux_v I__1999 (
            .O(N__9031),
            .I(N__9020));
    InMux I__1998 (
            .O(N__9030),
            .I(N__9015));
    InMux I__1997 (
            .O(N__9029),
            .I(N__9015));
    InMux I__1996 (
            .O(N__9026),
            .I(N__9012));
    Odrv4 I__1995 (
            .O(N__9023),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1994 (
            .O(N__9020),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1993 (
            .O(N__9015),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1992 (
            .O(N__9012),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1991 (
            .O(N__9003),
            .I(N__9000));
    LocalMux I__1990 (
            .O(N__9000),
            .I(N__8997));
    Span4Mux_s3_v I__1989 (
            .O(N__8997),
            .I(N__8994));
    Span4Mux_v I__1988 (
            .O(N__8994),
            .I(N__8991));
    Span4Mux_h I__1987 (
            .O(N__8991),
            .I(N__8988));
    Odrv4 I__1986 (
            .O(N__8988),
            .I(CRCSn_c));
    InMux I__1985 (
            .O(N__8985),
            .I(N__8982));
    LocalMux I__1984 (
            .O(N__8982),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1983 (
            .O(N__8979),
            .I(N__8976));
    LocalMux I__1982 (
            .O(N__8976),
            .I(N__8973));
    IoSpan4Mux I__1981 (
            .O(N__8973),
            .I(N__8970));
    Span4Mux_s0_h I__1980 (
            .O(N__8970),
            .I(N__8967));
    Sp12to4 I__1979 (
            .O(N__8967),
            .I(N__8964));
    Span12Mux_h I__1978 (
            .O(N__8964),
            .I(N__8961));
    Odrv12 I__1977 (
            .O(N__8961),
            .I(CMA_c_7));
    InMux I__1976 (
            .O(N__8958),
            .I(N__8955));
    LocalMux I__1975 (
            .O(N__8955),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1974 (
            .O(N__8952),
            .I(N__8949));
    LocalMux I__1973 (
            .O(N__8949),
            .I(N__8946));
    Span12Mux_s5_h I__1972 (
            .O(N__8946),
            .I(N__8943));
    Span12Mux_v I__1971 (
            .O(N__8943),
            .I(N__8940));
    Odrv12 I__1970 (
            .O(N__8940),
            .I(CMA_c_4));
    InMux I__1969 (
            .O(N__8937),
            .I(N__8934));
    LocalMux I__1968 (
            .O(N__8934),
            .I(N__8931));
    Span4Mux_h I__1967 (
            .O(N__8931),
            .I(N__8928));
    Span4Mux_h I__1966 (
            .O(N__8928),
            .I(N__8925));
    Odrv4 I__1965 (
            .O(N__8925),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1964 (
            .O(N__8922),
            .I(N__8919));
    LocalMux I__1963 (
            .O(N__8919),
            .I(N__8916));
    Odrv12 I__1962 (
            .O(N__8916),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1961 (
            .O(N__8913),
            .I(N__8910));
    LocalMux I__1960 (
            .O(N__8910),
            .I(N__8907));
    Span4Mux_h I__1959 (
            .O(N__8907),
            .I(N__8904));
    Odrv4 I__1958 (
            .O(N__8904),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1957 (
            .O(N__8901),
            .I(N__8894));
    InMux I__1956 (
            .O(N__8900),
            .I(N__8894));
    InMux I__1955 (
            .O(N__8899),
            .I(N__8891));
    LocalMux I__1954 (
            .O(N__8894),
            .I(N__8885));
    LocalMux I__1953 (
            .O(N__8891),
            .I(N__8885));
    InMux I__1952 (
            .O(N__8890),
            .I(N__8882));
    Span4Mux_v I__1951 (
            .O(N__8885),
            .I(N__8877));
    LocalMux I__1950 (
            .O(N__8882),
            .I(N__8877));
    Span4Mux_h I__1949 (
            .O(N__8877),
            .I(N__8874));
    Span4Mux_v I__1948 (
            .O(N__8874),
            .I(N__8871));
    Sp12to4 I__1947 (
            .O(N__8871),
            .I(N__8868));
    Odrv12 I__1946 (
            .O(N__8868),
            .I(DRA_c_2));
    InMux I__1945 (
            .O(N__8865),
            .I(N__8862));
    LocalMux I__1944 (
            .O(N__8862),
            .I(N__8859));
    Span4Mux_h I__1943 (
            .O(N__8859),
            .I(N__8856));
    Odrv4 I__1942 (
            .O(N__8856),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__1941 (
            .O(N__8853),
            .I(N__8850));
    InMux I__1940 (
            .O(N__8850),
            .I(N__8842));
    InMux I__1939 (
            .O(N__8849),
            .I(N__8842));
    InMux I__1938 (
            .O(N__8848),
            .I(N__8837));
    InMux I__1937 (
            .O(N__8847),
            .I(N__8837));
    LocalMux I__1936 (
            .O(N__8842),
            .I(N__8831));
    LocalMux I__1935 (
            .O(N__8837),
            .I(N__8831));
    CascadeMux I__1934 (
            .O(N__8836),
            .I(N__8827));
    Span4Mux_h I__1933 (
            .O(N__8831),
            .I(N__8817));
    InMux I__1932 (
            .O(N__8830),
            .I(N__8814));
    InMux I__1931 (
            .O(N__8827),
            .I(N__8811));
    InMux I__1930 (
            .O(N__8826),
            .I(N__8806));
    InMux I__1929 (
            .O(N__8825),
            .I(N__8803));
    InMux I__1928 (
            .O(N__8824),
            .I(N__8800));
    InMux I__1927 (
            .O(N__8823),
            .I(N__8795));
    InMux I__1926 (
            .O(N__8822),
            .I(N__8795));
    InMux I__1925 (
            .O(N__8821),
            .I(N__8789));
    InMux I__1924 (
            .O(N__8820),
            .I(N__8784));
    Span4Mux_v I__1923 (
            .O(N__8817),
            .I(N__8779));
    LocalMux I__1922 (
            .O(N__8814),
            .I(N__8779));
    LocalMux I__1921 (
            .O(N__8811),
            .I(N__8770));
    InMux I__1920 (
            .O(N__8810),
            .I(N__8765));
    InMux I__1919 (
            .O(N__8809),
            .I(N__8765));
    LocalMux I__1918 (
            .O(N__8806),
            .I(N__8762));
    LocalMux I__1917 (
            .O(N__8803),
            .I(N__8759));
    LocalMux I__1916 (
            .O(N__8800),
            .I(N__8754));
    LocalMux I__1915 (
            .O(N__8795),
            .I(N__8754));
    InMux I__1914 (
            .O(N__8794),
            .I(N__8747));
    InMux I__1913 (
            .O(N__8793),
            .I(N__8747));
    InMux I__1912 (
            .O(N__8792),
            .I(N__8747));
    LocalMux I__1911 (
            .O(N__8789),
            .I(N__8744));
    InMux I__1910 (
            .O(N__8788),
            .I(N__8741));
    InMux I__1909 (
            .O(N__8787),
            .I(N__8738));
    LocalMux I__1908 (
            .O(N__8784),
            .I(N__8735));
    Span4Mux_h I__1907 (
            .O(N__8779),
            .I(N__8732));
    InMux I__1906 (
            .O(N__8778),
            .I(N__8727));
    InMux I__1905 (
            .O(N__8777),
            .I(N__8727));
    InMux I__1904 (
            .O(N__8776),
            .I(N__8718));
    InMux I__1903 (
            .O(N__8775),
            .I(N__8718));
    InMux I__1902 (
            .O(N__8774),
            .I(N__8718));
    InMux I__1901 (
            .O(N__8773),
            .I(N__8718));
    Span4Mux_v I__1900 (
            .O(N__8770),
            .I(N__8709));
    LocalMux I__1899 (
            .O(N__8765),
            .I(N__8709));
    Span4Mux_v I__1898 (
            .O(N__8762),
            .I(N__8709));
    Span4Mux_v I__1897 (
            .O(N__8759),
            .I(N__8709));
    Span12Mux_v I__1896 (
            .O(N__8754),
            .I(N__8704));
    LocalMux I__1895 (
            .O(N__8747),
            .I(N__8704));
    Odrv4 I__1894 (
            .O(N__8744),
            .I(CPU_CYCLEm));
    LocalMux I__1893 (
            .O(N__8741),
            .I(CPU_CYCLEm));
    LocalMux I__1892 (
            .O(N__8738),
            .I(CPU_CYCLEm));
    Odrv4 I__1891 (
            .O(N__8735),
            .I(CPU_CYCLEm));
    Odrv4 I__1890 (
            .O(N__8732),
            .I(CPU_CYCLEm));
    LocalMux I__1889 (
            .O(N__8727),
            .I(CPU_CYCLEm));
    LocalMux I__1888 (
            .O(N__8718),
            .I(CPU_CYCLEm));
    Odrv4 I__1887 (
            .O(N__8709),
            .I(CPU_CYCLEm));
    Odrv12 I__1886 (
            .O(N__8704),
            .I(CPU_CYCLEm));
    CascadeMux I__1885 (
            .O(N__8685),
            .I(N__8682));
    InMux I__1884 (
            .O(N__8682),
            .I(N__8679));
    LocalMux I__1883 (
            .O(N__8679),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1882 (
            .O(N__8676),
            .I(N__8673));
    LocalMux I__1881 (
            .O(N__8673),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1880 (
            .O(N__8670),
            .I(N__8667));
    LocalMux I__1879 (
            .O(N__8667),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1878 (
            .O(N__8664),
            .I(N__8661));
    LocalMux I__1877 (
            .O(N__8661),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1876 (
            .O(N__8658),
            .I(N__8655));
    LocalMux I__1875 (
            .O(N__8655),
            .I(N__8652));
    Span4Mux_v I__1874 (
            .O(N__8652),
            .I(N__8649));
    Odrv4 I__1873 (
            .O(N__8649),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1872 (
            .O(N__8646),
            .I(N__8643));
    LocalMux I__1871 (
            .O(N__8643),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1870 (
            .O(N__8640),
            .I(N__8634));
    InMux I__1869 (
            .O(N__8639),
            .I(N__8634));
    LocalMux I__1868 (
            .O(N__8634),
            .I(N__8631));
    Span4Mux_h I__1867 (
            .O(N__8631),
            .I(N__8628));
    Odrv4 I__1866 (
            .O(N__8628),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1865 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__1864 (
            .O(N__8622),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1863 (
            .O(N__8619),
            .I(N__8615));
    InMux I__1862 (
            .O(N__8618),
            .I(N__8610));
    LocalMux I__1861 (
            .O(N__8615),
            .I(N__8607));
    InMux I__1860 (
            .O(N__8614),
            .I(N__8604));
    InMux I__1859 (
            .O(N__8613),
            .I(N__8601));
    LocalMux I__1858 (
            .O(N__8610),
            .I(N__8598));
    Span4Mux_h I__1857 (
            .O(N__8607),
            .I(N__8591));
    LocalMux I__1856 (
            .O(N__8604),
            .I(N__8591));
    LocalMux I__1855 (
            .O(N__8601),
            .I(N__8591));
    Span4Mux_h I__1854 (
            .O(N__8598),
            .I(N__8586));
    Span4Mux_h I__1853 (
            .O(N__8591),
            .I(N__8586));
    Span4Mux_v I__1852 (
            .O(N__8586),
            .I(N__8583));
    Span4Mux_v I__1851 (
            .O(N__8583),
            .I(N__8580));
    Span4Mux_v I__1850 (
            .O(N__8580),
            .I(N__8577));
    Span4Mux_v I__1849 (
            .O(N__8577),
            .I(N__8574));
    Odrv4 I__1848 (
            .O(N__8574),
            .I(CLK40_PLL_i));
    IoInMux I__1847 (
            .O(N__8571),
            .I(N__8566));
    IoInMux I__1846 (
            .O(N__8570),
            .I(N__8563));
    IoInMux I__1845 (
            .O(N__8569),
            .I(N__8560));
    LocalMux I__1844 (
            .O(N__8566),
            .I(N__8557));
    LocalMux I__1843 (
            .O(N__8563),
            .I(N__8554));
    LocalMux I__1842 (
            .O(N__8560),
            .I(N__8551));
    IoSpan4Mux I__1841 (
            .O(N__8557),
            .I(N__8548));
    Span4Mux_s3_v I__1840 (
            .O(N__8554),
            .I(N__8545));
    Span4Mux_s2_h I__1839 (
            .O(N__8551),
            .I(N__8542));
    IoSpan4Mux I__1838 (
            .O(N__8548),
            .I(N__8539));
    Span4Mux_h I__1837 (
            .O(N__8545),
            .I(N__8536));
    Span4Mux_v I__1836 (
            .O(N__8542),
            .I(N__8533));
    Sp12to4 I__1835 (
            .O(N__8539),
            .I(N__8528));
    Sp12to4 I__1834 (
            .O(N__8536),
            .I(N__8528));
    Sp12to4 I__1833 (
            .O(N__8533),
            .I(N__8525));
    Span12Mux_v I__1832 (
            .O(N__8528),
            .I(N__8520));
    Span12Mux_h I__1831 (
            .O(N__8525),
            .I(N__8520));
    Odrv12 I__1830 (
            .O(N__8520),
            .I(CLK40_PLL_i_i));
    IoInMux I__1829 (
            .O(N__8517),
            .I(N__8514));
    LocalMux I__1828 (
            .O(N__8514),
            .I(N__8511));
    Span4Mux_s2_v I__1827 (
            .O(N__8511),
            .I(N__8508));
    Span4Mux_h I__1826 (
            .O(N__8508),
            .I(N__8505));
    Span4Mux_v I__1825 (
            .O(N__8505),
            .I(N__8502));
    Odrv4 I__1824 (
            .O(N__8502),
            .I(UMBEn_c));
    CascadeMux I__1823 (
            .O(N__8499),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__1822 (
            .O(N__8496),
            .I(N__8493));
    LocalMux I__1821 (
            .O(N__8493),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1820 (
            .O(N__8490),
            .I(N__8487));
    LocalMux I__1819 (
            .O(N__8487),
            .I(N__8483));
    InMux I__1818 (
            .O(N__8486),
            .I(N__8475));
    Span4Mux_h I__1817 (
            .O(N__8483),
            .I(N__8472));
    InMux I__1816 (
            .O(N__8482),
            .I(N__8465));
    InMux I__1815 (
            .O(N__8481),
            .I(N__8465));
    InMux I__1814 (
            .O(N__8480),
            .I(N__8465));
    InMux I__1813 (
            .O(N__8479),
            .I(N__8460));
    InMux I__1812 (
            .O(N__8478),
            .I(N__8460));
    LocalMux I__1811 (
            .O(N__8475),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    Odrv4 I__1810 (
            .O(N__8472),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1809 (
            .O(N__8465),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1808 (
            .O(N__8460),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__1807 (
            .O(N__8451),
            .I(N__8448));
    LocalMux I__1806 (
            .O(N__8448),
            .I(N__8444));
    InMux I__1805 (
            .O(N__8447),
            .I(N__8441));
    Span4Mux_h I__1804 (
            .O(N__8444),
            .I(N__8436));
    LocalMux I__1803 (
            .O(N__8441),
            .I(N__8436));
    Span4Mux_h I__1802 (
            .O(N__8436),
            .I(N__8431));
    InMux I__1801 (
            .O(N__8435),
            .I(N__8426));
    InMux I__1800 (
            .O(N__8434),
            .I(N__8426));
    Odrv4 I__1799 (
            .O(N__8431),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1798 (
            .O(N__8426),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__1797 (
            .O(N__8421),
            .I(\U712_REG_SM.N_236_cascade_ ));
    CascadeMux I__1796 (
            .O(N__8418),
            .I(N__8415));
    InMux I__1795 (
            .O(N__8415),
            .I(N__8409));
    InMux I__1794 (
            .O(N__8414),
            .I(N__8404));
    InMux I__1793 (
            .O(N__8413),
            .I(N__8404));
    InMux I__1792 (
            .O(N__8412),
            .I(N__8401));
    LocalMux I__1791 (
            .O(N__8409),
            .I(N__8389));
    LocalMux I__1790 (
            .O(N__8404),
            .I(N__8389));
    LocalMux I__1789 (
            .O(N__8401),
            .I(N__8386));
    InMux I__1788 (
            .O(N__8400),
            .I(N__8379));
    InMux I__1787 (
            .O(N__8399),
            .I(N__8379));
    InMux I__1786 (
            .O(N__8398),
            .I(N__8379));
    InMux I__1785 (
            .O(N__8397),
            .I(N__8376));
    InMux I__1784 (
            .O(N__8396),
            .I(N__8373));
    InMux I__1783 (
            .O(N__8395),
            .I(N__8368));
    InMux I__1782 (
            .O(N__8394),
            .I(N__8368));
    Span4Mux_h I__1781 (
            .O(N__8389),
            .I(N__8365));
    Odrv4 I__1780 (
            .O(N__8386),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1779 (
            .O(N__8379),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1778 (
            .O(N__8376),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1777 (
            .O(N__8373),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1776 (
            .O(N__8368),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1775 (
            .O(N__8365),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1774 (
            .O(N__8352),
            .I(N__8348));
    CascadeMux I__1773 (
            .O(N__8351),
            .I(N__8343));
    InMux I__1772 (
            .O(N__8348),
            .I(N__8338));
    InMux I__1771 (
            .O(N__8347),
            .I(N__8335));
    InMux I__1770 (
            .O(N__8346),
            .I(N__8332));
    InMux I__1769 (
            .O(N__8343),
            .I(N__8327));
    InMux I__1768 (
            .O(N__8342),
            .I(N__8327));
    InMux I__1767 (
            .O(N__8341),
            .I(N__8324));
    LocalMux I__1766 (
            .O(N__8338),
            .I(N__8317));
    LocalMux I__1765 (
            .O(N__8335),
            .I(N__8317));
    LocalMux I__1764 (
            .O(N__8332),
            .I(N__8317));
    LocalMux I__1763 (
            .O(N__8327),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1762 (
            .O(N__8324),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv12 I__1761 (
            .O(N__8317),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__1760 (
            .O(N__8310),
            .I(N__8297));
    InMux I__1759 (
            .O(N__8309),
            .I(N__8291));
    InMux I__1758 (
            .O(N__8308),
            .I(N__8291));
    CascadeMux I__1757 (
            .O(N__8307),
            .I(N__8288));
    CascadeMux I__1756 (
            .O(N__8306),
            .I(N__8285));
    InMux I__1755 (
            .O(N__8305),
            .I(N__8282));
    InMux I__1754 (
            .O(N__8304),
            .I(N__8277));
    InMux I__1753 (
            .O(N__8303),
            .I(N__8277));
    InMux I__1752 (
            .O(N__8302),
            .I(N__8273));
    InMux I__1751 (
            .O(N__8301),
            .I(N__8264));
    InMux I__1750 (
            .O(N__8300),
            .I(N__8264));
    InMux I__1749 (
            .O(N__8297),
            .I(N__8264));
    InMux I__1748 (
            .O(N__8296),
            .I(N__8264));
    LocalMux I__1747 (
            .O(N__8291),
            .I(N__8261));
    InMux I__1746 (
            .O(N__8288),
            .I(N__8258));
    InMux I__1745 (
            .O(N__8285),
            .I(N__8255));
    LocalMux I__1744 (
            .O(N__8282),
            .I(N__8250));
    LocalMux I__1743 (
            .O(N__8277),
            .I(N__8250));
    InMux I__1742 (
            .O(N__8276),
            .I(N__8247));
    LocalMux I__1741 (
            .O(N__8273),
            .I(N__8242));
    LocalMux I__1740 (
            .O(N__8264),
            .I(N__8242));
    Span4Mux_v I__1739 (
            .O(N__8261),
            .I(N__8239));
    LocalMux I__1738 (
            .O(N__8258),
            .I(N__8232));
    LocalMux I__1737 (
            .O(N__8255),
            .I(N__8232));
    Span4Mux_v I__1736 (
            .O(N__8250),
            .I(N__8232));
    LocalMux I__1735 (
            .O(N__8247),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1734 (
            .O(N__8242),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1733 (
            .O(N__8239),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1732 (
            .O(N__8232),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__1731 (
            .O(N__8223),
            .I(N__8220));
    LocalMux I__1730 (
            .O(N__8220),
            .I(\U712_REG_SM.N_273 ));
    InMux I__1729 (
            .O(N__8217),
            .I(N__8208));
    InMux I__1728 (
            .O(N__8216),
            .I(N__8208));
    InMux I__1727 (
            .O(N__8215),
            .I(N__8203));
    InMux I__1726 (
            .O(N__8214),
            .I(N__8203));
    CascadeMux I__1725 (
            .O(N__8213),
            .I(N__8199));
    LocalMux I__1724 (
            .O(N__8208),
            .I(N__8181));
    LocalMux I__1723 (
            .O(N__8203),
            .I(N__8181));
    InMux I__1722 (
            .O(N__8202),
            .I(N__8176));
    InMux I__1721 (
            .O(N__8199),
            .I(N__8176));
    InMux I__1720 (
            .O(N__8198),
            .I(N__8173));
    InMux I__1719 (
            .O(N__8197),
            .I(N__8168));
    InMux I__1718 (
            .O(N__8196),
            .I(N__8168));
    InMux I__1717 (
            .O(N__8195),
            .I(N__8165));
    InMux I__1716 (
            .O(N__8194),
            .I(N__8162));
    InMux I__1715 (
            .O(N__8193),
            .I(N__8156));
    InMux I__1714 (
            .O(N__8192),
            .I(N__8156));
    InMux I__1713 (
            .O(N__8191),
            .I(N__8153));
    InMux I__1712 (
            .O(N__8190),
            .I(N__8148));
    InMux I__1711 (
            .O(N__8189),
            .I(N__8148));
    InMux I__1710 (
            .O(N__8188),
            .I(N__8141));
    InMux I__1709 (
            .O(N__8187),
            .I(N__8141));
    InMux I__1708 (
            .O(N__8186),
            .I(N__8141));
    Span4Mux_v I__1707 (
            .O(N__8181),
            .I(N__8132));
    LocalMux I__1706 (
            .O(N__8176),
            .I(N__8132));
    LocalMux I__1705 (
            .O(N__8173),
            .I(N__8132));
    LocalMux I__1704 (
            .O(N__8168),
            .I(N__8132));
    LocalMux I__1703 (
            .O(N__8165),
            .I(N__8122));
    LocalMux I__1702 (
            .O(N__8162),
            .I(N__8119));
    InMux I__1701 (
            .O(N__8161),
            .I(N__8116));
    LocalMux I__1700 (
            .O(N__8156),
            .I(N__8104));
    LocalMux I__1699 (
            .O(N__8153),
            .I(N__8104));
    LocalMux I__1698 (
            .O(N__8148),
            .I(N__8104));
    LocalMux I__1697 (
            .O(N__8141),
            .I(N__8104));
    Span4Mux_v I__1696 (
            .O(N__8132),
            .I(N__8104));
    InMux I__1695 (
            .O(N__8131),
            .I(N__8101));
    InMux I__1694 (
            .O(N__8130),
            .I(N__8096));
    InMux I__1693 (
            .O(N__8129),
            .I(N__8096));
    InMux I__1692 (
            .O(N__8128),
            .I(N__8092));
    InMux I__1691 (
            .O(N__8127),
            .I(N__8085));
    InMux I__1690 (
            .O(N__8126),
            .I(N__8085));
    InMux I__1689 (
            .O(N__8125),
            .I(N__8085));
    Span4Mux_v I__1688 (
            .O(N__8122),
            .I(N__8078));
    Span4Mux_v I__1687 (
            .O(N__8119),
            .I(N__8078));
    LocalMux I__1686 (
            .O(N__8116),
            .I(N__8078));
    InMux I__1685 (
            .O(N__8115),
            .I(N__8075));
    Span4Mux_v I__1684 (
            .O(N__8104),
            .I(N__8067));
    LocalMux I__1683 (
            .O(N__8101),
            .I(N__8064));
    LocalMux I__1682 (
            .O(N__8096),
            .I(N__8061));
    InMux I__1681 (
            .O(N__8095),
            .I(N__8058));
    LocalMux I__1680 (
            .O(N__8092),
            .I(N__8049));
    LocalMux I__1679 (
            .O(N__8085),
            .I(N__8049));
    Span4Mux_h I__1678 (
            .O(N__8078),
            .I(N__8049));
    LocalMux I__1677 (
            .O(N__8075),
            .I(N__8049));
    InMux I__1676 (
            .O(N__8074),
            .I(N__8044));
    InMux I__1675 (
            .O(N__8073),
            .I(N__8044));
    InMux I__1674 (
            .O(N__8072),
            .I(N__8037));
    InMux I__1673 (
            .O(N__8071),
            .I(N__8037));
    InMux I__1672 (
            .O(N__8070),
            .I(N__8037));
    Span4Mux_h I__1671 (
            .O(N__8067),
            .I(N__8030));
    Span4Mux_v I__1670 (
            .O(N__8064),
            .I(N__8030));
    Span4Mux_v I__1669 (
            .O(N__8061),
            .I(N__8030));
    LocalMux I__1668 (
            .O(N__8058),
            .I(N__8021));
    Sp12to4 I__1667 (
            .O(N__8049),
            .I(N__8021));
    LocalMux I__1666 (
            .O(N__8044),
            .I(N__8021));
    LocalMux I__1665 (
            .O(N__8037),
            .I(N__8021));
    Span4Mux_h I__1664 (
            .O(N__8030),
            .I(N__8018));
    Span12Mux_v I__1663 (
            .O(N__8021),
            .I(N__8015));
    Span4Mux_h I__1662 (
            .O(N__8018),
            .I(N__8012));
    Span12Mux_h I__1661 (
            .O(N__8015),
            .I(N__8009));
    Span4Mux_h I__1660 (
            .O(N__8012),
            .I(N__8006));
    Odrv12 I__1659 (
            .O(N__8009),
            .I(RESETn_c));
    Odrv4 I__1658 (
            .O(N__8006),
            .I(RESETn_c));
    InMux I__1657 (
            .O(N__8001),
            .I(N__7995));
    InMux I__1656 (
            .O(N__8000),
            .I(N__7995));
    LocalMux I__1655 (
            .O(N__7995),
            .I(N__7992));
    Odrv12 I__1654 (
            .O(N__7992),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1653 (
            .O(N__7989),
            .I(N__7986));
    LocalMux I__1652 (
            .O(N__7986),
            .I(N__7983));
    Span4Mux_v I__1651 (
            .O(N__7983),
            .I(N__7980));
    Sp12to4 I__1650 (
            .O(N__7980),
            .I(N__7977));
    Span12Mux_h I__1649 (
            .O(N__7977),
            .I(N__7974));
    Span12Mux_v I__1648 (
            .O(N__7974),
            .I(N__7971));
    Odrv12 I__1647 (
            .O(N__7971),
            .I(A_c_19));
    CascadeMux I__1646 (
            .O(N__7968),
            .I(N__7965));
    InMux I__1645 (
            .O(N__7965),
            .I(N__7961));
    InMux I__1644 (
            .O(N__7964),
            .I(N__7958));
    LocalMux I__1643 (
            .O(N__7961),
            .I(N__7952));
    LocalMux I__1642 (
            .O(N__7958),
            .I(N__7952));
    CascadeMux I__1641 (
            .O(N__7957),
            .I(N__7949));
    Span4Mux_h I__1640 (
            .O(N__7952),
            .I(N__7945));
    InMux I__1639 (
            .O(N__7949),
            .I(N__7940));
    InMux I__1638 (
            .O(N__7948),
            .I(N__7940));
    Odrv4 I__1637 (
            .O(N__7945),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1636 (
            .O(N__7940),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    IoInMux I__1635 (
            .O(N__7935),
            .I(N__7932));
    LocalMux I__1634 (
            .O(N__7932),
            .I(N__7929));
    IoSpan4Mux I__1633 (
            .O(N__7929),
            .I(N__7926));
    IoSpan4Mux I__1632 (
            .O(N__7926),
            .I(N__7923));
    Span4Mux_s3_h I__1631 (
            .O(N__7923),
            .I(N__7920));
    Sp12to4 I__1630 (
            .O(N__7920),
            .I(N__7917));
    Odrv12 I__1629 (
            .O(N__7917),
            .I(CMA_c_9));
    CascadeMux I__1628 (
            .O(N__7914),
            .I(N__7911));
    InMux I__1627 (
            .O(N__7911),
            .I(N__7908));
    LocalMux I__1626 (
            .O(N__7908),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1625 (
            .O(N__7905),
            .I(N__7902));
    LocalMux I__1624 (
            .O(N__7902),
            .I(N__7899));
    Sp12to4 I__1623 (
            .O(N__7899),
            .I(N__7896));
    Span12Mux_v I__1622 (
            .O(N__7896),
            .I(N__7893));
    Span12Mux_h I__1621 (
            .O(N__7893),
            .I(N__7890));
    Odrv12 I__1620 (
            .O(N__7890),
            .I(A_c_16));
    InMux I__1619 (
            .O(N__7887),
            .I(N__7884));
    LocalMux I__1618 (
            .O(N__7884),
            .I(N__7881));
    Sp12to4 I__1617 (
            .O(N__7881),
            .I(N__7878));
    Span12Mux_v I__1616 (
            .O(N__7878),
            .I(N__7875));
    Span12Mux_h I__1615 (
            .O(N__7875),
            .I(N__7872));
    Odrv12 I__1614 (
            .O(N__7872),
            .I(A_c_18));
    CascadeMux I__1613 (
            .O(N__7869),
            .I(N__7866));
    InMux I__1612 (
            .O(N__7866),
            .I(N__7863));
    LocalMux I__1611 (
            .O(N__7863),
            .I(N__7860));
    Odrv12 I__1610 (
            .O(N__7860),
            .I(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ));
    InMux I__1609 (
            .O(N__7857),
            .I(N__7854));
    LocalMux I__1608 (
            .O(N__7854),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1607 (
            .O(N__7851),
            .I(N__7848));
    LocalMux I__1606 (
            .O(N__7848),
            .I(N__7845));
    Span4Mux_v I__1605 (
            .O(N__7845),
            .I(N__7842));
    Sp12to4 I__1604 (
            .O(N__7842),
            .I(N__7839));
    Span12Mux_h I__1603 (
            .O(N__7839),
            .I(N__7836));
    Odrv12 I__1602 (
            .O(N__7836),
            .I(A_c_6));
    InMux I__1601 (
            .O(N__7833),
            .I(N__7830));
    LocalMux I__1600 (
            .O(N__7830),
            .I(N__7827));
    Span4Mux_v I__1599 (
            .O(N__7827),
            .I(N__7824));
    Span4Mux_v I__1598 (
            .O(N__7824),
            .I(N__7821));
    Sp12to4 I__1597 (
            .O(N__7821),
            .I(N__7818));
    Span12Mux_h I__1596 (
            .O(N__7818),
            .I(N__7815));
    Odrv12 I__1595 (
            .O(N__7815),
            .I(A_c_13));
    InMux I__1594 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__1593 (
            .O(N__7809),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1592 (
            .O(N__7806),
            .I(N__7803));
    LocalMux I__1591 (
            .O(N__7803),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1590 (
            .O(N__7800),
            .I(N__7797));
    LocalMux I__1589 (
            .O(N__7797),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1588 (
            .O(N__7794),
            .I(N__7791));
    LocalMux I__1587 (
            .O(N__7791),
            .I(N__7788));
    Span12Mux_s4_v I__1586 (
            .O(N__7788),
            .I(N__7785));
    Span12Mux_v I__1585 (
            .O(N__7785),
            .I(N__7782));
    Odrv12 I__1584 (
            .O(N__7782),
            .I(CMA_c_2));
    InMux I__1583 (
            .O(N__7779),
            .I(N__7776));
    LocalMux I__1582 (
            .O(N__7776),
            .I(N__7773));
    Span4Mux_v I__1581 (
            .O(N__7773),
            .I(N__7770));
    Sp12to4 I__1580 (
            .O(N__7770),
            .I(N__7767));
    Span12Mux_h I__1579 (
            .O(N__7767),
            .I(N__7764));
    Odrv12 I__1578 (
            .O(N__7764),
            .I(A_c_5));
    InMux I__1577 (
            .O(N__7761),
            .I(N__7758));
    LocalMux I__1576 (
            .O(N__7758),
            .I(N__7755));
    Sp12to4 I__1575 (
            .O(N__7755),
            .I(N__7752));
    Span12Mux_v I__1574 (
            .O(N__7752),
            .I(N__7749));
    Span12Mux_h I__1573 (
            .O(N__7749),
            .I(N__7746));
    Odrv12 I__1572 (
            .O(N__7746),
            .I(A_c_12));
    InMux I__1571 (
            .O(N__7743),
            .I(N__7740));
    LocalMux I__1570 (
            .O(N__7740),
            .I(\U712_BYTE_ENABLE.N_314 ));
    CascadeMux I__1569 (
            .O(N__7737),
            .I(N__7734));
    InMux I__1568 (
            .O(N__7734),
            .I(N__7731));
    LocalMux I__1567 (
            .O(N__7731),
            .I(N__7728));
    Span4Mux_v I__1566 (
            .O(N__7728),
            .I(N__7725));
    Odrv4 I__1565 (
            .O(N__7725),
            .I(\U712_BYTE_ENABLE.UUBE ));
    IoInMux I__1564 (
            .O(N__7722),
            .I(N__7719));
    LocalMux I__1563 (
            .O(N__7719),
            .I(N__7716));
    Odrv12 I__1562 (
            .O(N__7716),
            .I(RESETn_c_i));
    IoInMux I__1561 (
            .O(N__7713),
            .I(N__7710));
    LocalMux I__1560 (
            .O(N__7710),
            .I(N__7707));
    Span12Mux_s3_h I__1559 (
            .O(N__7707),
            .I(N__7704));
    Span12Mux_h I__1558 (
            .O(N__7704),
            .I(N__7701));
    Odrv12 I__1557 (
            .O(N__7701),
            .I(WEn_c));
    IoInMux I__1556 (
            .O(N__7698),
            .I(N__7695));
    LocalMux I__1555 (
            .O(N__7695),
            .I(N__7692));
    Span4Mux_s2_v I__1554 (
            .O(N__7692),
            .I(N__7689));
    Span4Mux_v I__1553 (
            .O(N__7689),
            .I(N__7686));
    Sp12to4 I__1552 (
            .O(N__7686),
            .I(N__7683));
    Span12Mux_h I__1551 (
            .O(N__7683),
            .I(N__7680));
    Odrv12 I__1550 (
            .O(N__7680),
            .I(RASn_c));
    InMux I__1549 (
            .O(N__7677),
            .I(N__7673));
    InMux I__1548 (
            .O(N__7676),
            .I(N__7670));
    LocalMux I__1547 (
            .O(N__7673),
            .I(N__7667));
    LocalMux I__1546 (
            .O(N__7670),
            .I(N__7664));
    Span4Mux_h I__1545 (
            .O(N__7667),
            .I(N__7658));
    Span4Mux_h I__1544 (
            .O(N__7664),
            .I(N__7655));
    InMux I__1543 (
            .O(N__7663),
            .I(N__7652));
    CascadeMux I__1542 (
            .O(N__7662),
            .I(N__7648));
    InMux I__1541 (
            .O(N__7661),
            .I(N__7644));
    Span4Mux_v I__1540 (
            .O(N__7658),
            .I(N__7641));
    Span4Mux_v I__1539 (
            .O(N__7655),
            .I(N__7638));
    LocalMux I__1538 (
            .O(N__7652),
            .I(N__7635));
    InMux I__1537 (
            .O(N__7651),
            .I(N__7630));
    InMux I__1536 (
            .O(N__7648),
            .I(N__7630));
    InMux I__1535 (
            .O(N__7647),
            .I(N__7627));
    LocalMux I__1534 (
            .O(N__7644),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1533 (
            .O(N__7641),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1532 (
            .O(N__7638),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1531 (
            .O(N__7635),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1530 (
            .O(N__7630),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1529 (
            .O(N__7627),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1528 (
            .O(N__7614),
            .I(N__7609));
    InMux I__1527 (
            .O(N__7613),
            .I(N__7606));
    InMux I__1526 (
            .O(N__7612),
            .I(N__7603));
    LocalMux I__1525 (
            .O(N__7609),
            .I(N__7598));
    LocalMux I__1524 (
            .O(N__7606),
            .I(N__7598));
    LocalMux I__1523 (
            .O(N__7603),
            .I(N__7595));
    Span4Mux_v I__1522 (
            .O(N__7598),
            .I(N__7588));
    Span4Mux_h I__1521 (
            .O(N__7595),
            .I(N__7585));
    InMux I__1520 (
            .O(N__7594),
            .I(N__7578));
    InMux I__1519 (
            .O(N__7593),
            .I(N__7578));
    InMux I__1518 (
            .O(N__7592),
            .I(N__7578));
    InMux I__1517 (
            .O(N__7591),
            .I(N__7575));
    Odrv4 I__1516 (
            .O(N__7588),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1515 (
            .O(N__7585),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1514 (
            .O(N__7578),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1513 (
            .O(N__7575),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1512 (
            .O(N__7566),
            .I(N__7563));
    LocalMux I__1511 (
            .O(N__7563),
            .I(N__7560));
    Span4Mux_s0_v I__1510 (
            .O(N__7560),
            .I(N__7557));
    Sp12to4 I__1509 (
            .O(N__7557),
            .I(N__7554));
    Span12Mux_h I__1508 (
            .O(N__7554),
            .I(N__7551));
    Span12Mux_v I__1507 (
            .O(N__7551),
            .I(N__7548));
    Odrv12 I__1506 (
            .O(N__7548),
            .I(CMA_c_10));
    InMux I__1505 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__1504 (
            .O(N__7542),
            .I(N__7539));
    Span4Mux_v I__1503 (
            .O(N__7539),
            .I(N__7536));
    Span4Mux_v I__1502 (
            .O(N__7536),
            .I(N__7533));
    Sp12to4 I__1501 (
            .O(N__7533),
            .I(N__7530));
    Span12Mux_h I__1500 (
            .O(N__7530),
            .I(N__7527));
    Odrv12 I__1499 (
            .O(N__7527),
            .I(A_c_17));
    IoInMux I__1498 (
            .O(N__7524),
            .I(N__7521));
    LocalMux I__1497 (
            .O(N__7521),
            .I(N__7518));
    IoSpan4Mux I__1496 (
            .O(N__7518),
            .I(N__7515));
    Span4Mux_s1_h I__1495 (
            .O(N__7515),
            .I(N__7512));
    Sp12to4 I__1494 (
            .O(N__7512),
            .I(N__7509));
    Span12Mux_h I__1493 (
            .O(N__7509),
            .I(N__7506));
    Odrv12 I__1492 (
            .O(N__7506),
            .I(CMA_c_8));
    InMux I__1491 (
            .O(N__7503),
            .I(N__7500));
    LocalMux I__1490 (
            .O(N__7500),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    CascadeMux I__1489 (
            .O(N__7497),
            .I(\U712_REG_SM.N_235_cascade_ ));
    SRMux I__1488 (
            .O(N__7494),
            .I(N__7491));
    LocalMux I__1487 (
            .O(N__7491),
            .I(N__7488));
    Span4Mux_h I__1486 (
            .O(N__7488),
            .I(N__7485));
    Odrv4 I__1485 (
            .O(N__7485),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1484 (
            .O(N__7482),
            .I(N__7479));
    LocalMux I__1483 (
            .O(N__7479),
            .I(\U712_REG_SM.N_281 ));
    InMux I__1482 (
            .O(N__7476),
            .I(N__7473));
    LocalMux I__1481 (
            .O(N__7473),
            .I(\U712_REG_SM.N_235 ));
    InMux I__1480 (
            .O(N__7470),
            .I(N__7467));
    LocalMux I__1479 (
            .O(N__7467),
            .I(N__7463));
    InMux I__1478 (
            .O(N__7466),
            .I(N__7460));
    Odrv4 I__1477 (
            .O(N__7463),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1476 (
            .O(N__7460),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1475 (
            .O(N__7455),
            .I(N__7452));
    LocalMux I__1474 (
            .O(N__7452),
            .I(N__7446));
    InMux I__1473 (
            .O(N__7451),
            .I(N__7443));
    InMux I__1472 (
            .O(N__7450),
            .I(N__7440));
    InMux I__1471 (
            .O(N__7449),
            .I(N__7437));
    Odrv12 I__1470 (
            .O(N__7446),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1469 (
            .O(N__7443),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1468 (
            .O(N__7440),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1467 (
            .O(N__7437),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__1466 (
            .O(N__7428),
            .I(N__7425));
    InMux I__1465 (
            .O(N__7425),
            .I(N__7422));
    LocalMux I__1464 (
            .O(N__7422),
            .I(N__7419));
    Odrv12 I__1463 (
            .O(N__7419),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    InMux I__1462 (
            .O(N__7416),
            .I(N__7412));
    CascadeMux I__1461 (
            .O(N__7415),
            .I(N__7409));
    LocalMux I__1460 (
            .O(N__7412),
            .I(N__7405));
    InMux I__1459 (
            .O(N__7409),
            .I(N__7402));
    InMux I__1458 (
            .O(N__7408),
            .I(N__7399));
    Span4Mux_h I__1457 (
            .O(N__7405),
            .I(N__7396));
    LocalMux I__1456 (
            .O(N__7402),
            .I(N__7393));
    LocalMux I__1455 (
            .O(N__7399),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1454 (
            .O(N__7396),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1453 (
            .O(N__7393),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1452 (
            .O(N__7386),
            .I(N__7382));
    InMux I__1451 (
            .O(N__7385),
            .I(N__7379));
    LocalMux I__1450 (
            .O(N__7382),
            .I(N__7374));
    LocalMux I__1449 (
            .O(N__7379),
            .I(N__7371));
    InMux I__1448 (
            .O(N__7378),
            .I(N__7366));
    InMux I__1447 (
            .O(N__7377),
            .I(N__7366));
    Span12Mux_v I__1446 (
            .O(N__7374),
            .I(N__7363));
    Span4Mux_v I__1445 (
            .O(N__7371),
            .I(N__7360));
    LocalMux I__1444 (
            .O(N__7366),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv12 I__1443 (
            .O(N__7363),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__1442 (
            .O(N__7360),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1441 (
            .O(N__7353),
            .I(N__7349));
    InMux I__1440 (
            .O(N__7352),
            .I(N__7345));
    LocalMux I__1439 (
            .O(N__7349),
            .I(N__7342));
    InMux I__1438 (
            .O(N__7348),
            .I(N__7339));
    LocalMux I__1437 (
            .O(N__7345),
            .I(\U712_REG_SM.N_212 ));
    Odrv12 I__1436 (
            .O(N__7342),
            .I(\U712_REG_SM.N_212 ));
    LocalMux I__1435 (
            .O(N__7339),
            .I(\U712_REG_SM.N_212 ));
    InMux I__1434 (
            .O(N__7332),
            .I(N__7329));
    LocalMux I__1433 (
            .O(N__7329),
            .I(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ));
    CascadeMux I__1432 (
            .O(N__7326),
            .I(N__7323));
    InMux I__1431 (
            .O(N__7323),
            .I(N__7318));
    InMux I__1430 (
            .O(N__7322),
            .I(N__7313));
    InMux I__1429 (
            .O(N__7321),
            .I(N__7313));
    LocalMux I__1428 (
            .O(N__7318),
            .I(REG_TACK));
    LocalMux I__1427 (
            .O(N__7313),
            .I(REG_TACK));
    IoInMux I__1426 (
            .O(N__7308),
            .I(N__7305));
    LocalMux I__1425 (
            .O(N__7305),
            .I(N__7302));
    IoSpan4Mux I__1424 (
            .O(N__7302),
            .I(N__7299));
    Span4Mux_s3_h I__1423 (
            .O(N__7299),
            .I(N__7296));
    Span4Mux_v I__1422 (
            .O(N__7296),
            .I(N__7293));
    Span4Mux_v I__1421 (
            .O(N__7293),
            .I(N__7289));
    InMux I__1420 (
            .O(N__7292),
            .I(N__7286));
    Sp12to4 I__1419 (
            .O(N__7289),
            .I(N__7283));
    LocalMux I__1418 (
            .O(N__7286),
            .I(N__7280));
    Span12Mux_h I__1417 (
            .O(N__7283),
            .I(N__7275));
    Span12Mux_v I__1416 (
            .O(N__7280),
            .I(N__7275));
    Span12Mux_h I__1415 (
            .O(N__7275),
            .I(N__7272));
    Odrv12 I__1414 (
            .O(N__7272),
            .I(C3_c));
    InMux I__1413 (
            .O(N__7269),
            .I(N__7266));
    LocalMux I__1412 (
            .O(N__7266),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1411 (
            .O(N__7263),
            .I(N__7260));
    LocalMux I__1410 (
            .O(N__7260),
            .I(N__7256));
    InMux I__1409 (
            .O(N__7259),
            .I(N__7253));
    Span4Mux_v I__1408 (
            .O(N__7256),
            .I(N__7250));
    LocalMux I__1407 (
            .O(N__7253),
            .I(N__7247));
    Odrv4 I__1406 (
            .O(N__7250),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ));
    Odrv4 I__1405 (
            .O(N__7247),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ));
    CascadeMux I__1404 (
            .O(N__7242),
            .I(\U712_BYTE_ENABLE.N_220_cascade_ ));
    IoInMux I__1403 (
            .O(N__7239),
            .I(N__7236));
    LocalMux I__1402 (
            .O(N__7236),
            .I(N__7233));
    IoSpan4Mux I__1401 (
            .O(N__7233),
            .I(N__7230));
    IoSpan4Mux I__1400 (
            .O(N__7230),
            .I(N__7227));
    Span4Mux_s3_h I__1399 (
            .O(N__7227),
            .I(N__7224));
    Sp12to4 I__1398 (
            .O(N__7224),
            .I(N__7221));
    Span12Mux_h I__1397 (
            .O(N__7221),
            .I(N__7218));
    Span12Mux_v I__1396 (
            .O(N__7218),
            .I(N__7215));
    Odrv12 I__1395 (
            .O(N__7215),
            .I(N_151_i));
    InMux I__1394 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1393 (
            .O(N__7209),
            .I(N__7205));
    InMux I__1392 (
            .O(N__7208),
            .I(N__7201));
    Span4Mux_h I__1391 (
            .O(N__7205),
            .I(N__7198));
    InMux I__1390 (
            .O(N__7204),
            .I(N__7195));
    LocalMux I__1389 (
            .O(N__7201),
            .I(N__7192));
    Odrv4 I__1388 (
            .O(N__7198),
            .I(\U712_CHIP_RAM.N_386 ));
    LocalMux I__1387 (
            .O(N__7195),
            .I(\U712_CHIP_RAM.N_386 ));
    Odrv4 I__1386 (
            .O(N__7192),
            .I(\U712_CHIP_RAM.N_386 ));
    CascadeMux I__1385 (
            .O(N__7185),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__1384 (
            .O(N__7182),
            .I(N__7176));
    InMux I__1383 (
            .O(N__7181),
            .I(N__7170));
    InMux I__1382 (
            .O(N__7180),
            .I(N__7167));
    InMux I__1381 (
            .O(N__7179),
            .I(N__7164));
    InMux I__1380 (
            .O(N__7176),
            .I(N__7159));
    InMux I__1379 (
            .O(N__7175),
            .I(N__7159));
    InMux I__1378 (
            .O(N__7174),
            .I(N__7149));
    CascadeMux I__1377 (
            .O(N__7173),
            .I(N__7146));
    LocalMux I__1376 (
            .O(N__7170),
            .I(N__7139));
    LocalMux I__1375 (
            .O(N__7167),
            .I(N__7139));
    LocalMux I__1374 (
            .O(N__7164),
            .I(N__7134));
    LocalMux I__1373 (
            .O(N__7159),
            .I(N__7134));
    InMux I__1372 (
            .O(N__7158),
            .I(N__7130));
    InMux I__1371 (
            .O(N__7157),
            .I(N__7125));
    InMux I__1370 (
            .O(N__7156),
            .I(N__7125));
    InMux I__1369 (
            .O(N__7155),
            .I(N__7122));
    InMux I__1368 (
            .O(N__7154),
            .I(N__7119));
    InMux I__1367 (
            .O(N__7153),
            .I(N__7114));
    InMux I__1366 (
            .O(N__7152),
            .I(N__7114));
    LocalMux I__1365 (
            .O(N__7149),
            .I(N__7111));
    InMux I__1364 (
            .O(N__7146),
            .I(N__7108));
    InMux I__1363 (
            .O(N__7145),
            .I(N__7105));
    InMux I__1362 (
            .O(N__7144),
            .I(N__7102));
    Span4Mux_v I__1361 (
            .O(N__7139),
            .I(N__7097));
    Span4Mux_v I__1360 (
            .O(N__7134),
            .I(N__7097));
    InMux I__1359 (
            .O(N__7133),
            .I(N__7094));
    LocalMux I__1358 (
            .O(N__7130),
            .I(N__7091));
    LocalMux I__1357 (
            .O(N__7125),
            .I(N__7088));
    LocalMux I__1356 (
            .O(N__7122),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1355 (
            .O(N__7119),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1354 (
            .O(N__7114),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1353 (
            .O(N__7111),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1352 (
            .O(N__7108),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1351 (
            .O(N__7105),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1350 (
            .O(N__7102),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1349 (
            .O(N__7097),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1348 (
            .O(N__7094),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1347 (
            .O(N__7091),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1346 (
            .O(N__7088),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1345 (
            .O(N__7065),
            .I(N__7061));
    CascadeMux I__1344 (
            .O(N__7064),
            .I(N__7055));
    InMux I__1343 (
            .O(N__7061),
            .I(N__7052));
    InMux I__1342 (
            .O(N__7060),
            .I(N__7046));
    InMux I__1341 (
            .O(N__7059),
            .I(N__7040));
    InMux I__1340 (
            .O(N__7058),
            .I(N__7034));
    InMux I__1339 (
            .O(N__7055),
            .I(N__7034));
    LocalMux I__1338 (
            .O(N__7052),
            .I(N__7031));
    InMux I__1337 (
            .O(N__7051),
            .I(N__7026));
    InMux I__1336 (
            .O(N__7050),
            .I(N__7026));
    InMux I__1335 (
            .O(N__7049),
            .I(N__7015));
    LocalMux I__1334 (
            .O(N__7046),
            .I(N__7012));
    InMux I__1333 (
            .O(N__7045),
            .I(N__7009));
    InMux I__1332 (
            .O(N__7044),
            .I(N__7004));
    InMux I__1331 (
            .O(N__7043),
            .I(N__7004));
    LocalMux I__1330 (
            .O(N__7040),
            .I(N__7001));
    InMux I__1329 (
            .O(N__7039),
            .I(N__6998));
    LocalMux I__1328 (
            .O(N__7034),
            .I(N__6995));
    Span4Mux_v I__1327 (
            .O(N__7031),
            .I(N__6990));
    LocalMux I__1326 (
            .O(N__7026),
            .I(N__6990));
    InMux I__1325 (
            .O(N__7025),
            .I(N__6985));
    InMux I__1324 (
            .O(N__7024),
            .I(N__6985));
    InMux I__1323 (
            .O(N__7023),
            .I(N__6976));
    InMux I__1322 (
            .O(N__7022),
            .I(N__6976));
    InMux I__1321 (
            .O(N__7021),
            .I(N__6976));
    InMux I__1320 (
            .O(N__7020),
            .I(N__6976));
    InMux I__1319 (
            .O(N__7019),
            .I(N__6971));
    InMux I__1318 (
            .O(N__7018),
            .I(N__6971));
    LocalMux I__1317 (
            .O(N__7015),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1316 (
            .O(N__7012),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1315 (
            .O(N__7009),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1314 (
            .O(N__7004),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1313 (
            .O(N__7001),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1312 (
            .O(N__6998),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1311 (
            .O(N__6995),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1310 (
            .O(N__6990),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1309 (
            .O(N__6985),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1308 (
            .O(N__6976),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1307 (
            .O(N__6971),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1306 (
            .O(N__6948),
            .I(N__6944));
    InMux I__1305 (
            .O(N__6947),
            .I(N__6938));
    InMux I__1304 (
            .O(N__6944),
            .I(N__6934));
    CascadeMux I__1303 (
            .O(N__6943),
            .I(N__6931));
    InMux I__1302 (
            .O(N__6942),
            .I(N__6926));
    InMux I__1301 (
            .O(N__6941),
            .I(N__6926));
    LocalMux I__1300 (
            .O(N__6938),
            .I(N__6923));
    InMux I__1299 (
            .O(N__6937),
            .I(N__6918));
    LocalMux I__1298 (
            .O(N__6934),
            .I(N__6915));
    InMux I__1297 (
            .O(N__6931),
            .I(N__6912));
    LocalMux I__1296 (
            .O(N__6926),
            .I(N__6909));
    Span4Mux_h I__1295 (
            .O(N__6923),
            .I(N__6906));
    InMux I__1294 (
            .O(N__6922),
            .I(N__6901));
    InMux I__1293 (
            .O(N__6921),
            .I(N__6901));
    LocalMux I__1292 (
            .O(N__6918),
            .I(\U712_CHIP_RAM.N_338 ));
    Odrv4 I__1291 (
            .O(N__6915),
            .I(\U712_CHIP_RAM.N_338 ));
    LocalMux I__1290 (
            .O(N__6912),
            .I(\U712_CHIP_RAM.N_338 ));
    Odrv4 I__1289 (
            .O(N__6909),
            .I(\U712_CHIP_RAM.N_338 ));
    Odrv4 I__1288 (
            .O(N__6906),
            .I(\U712_CHIP_RAM.N_338 ));
    LocalMux I__1287 (
            .O(N__6901),
            .I(\U712_CHIP_RAM.N_338 ));
    InMux I__1286 (
            .O(N__6888),
            .I(N__6884));
    InMux I__1285 (
            .O(N__6887),
            .I(N__6881));
    LocalMux I__1284 (
            .O(N__6884),
            .I(N__6876));
    LocalMux I__1283 (
            .O(N__6881),
            .I(N__6876));
    Span4Mux_h I__1282 (
            .O(N__6876),
            .I(N__6873));
    Odrv4 I__1281 (
            .O(N__6873),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2 ));
    InMux I__1280 (
            .O(N__6870),
            .I(N__6865));
    InMux I__1279 (
            .O(N__6869),
            .I(N__6862));
    InMux I__1278 (
            .O(N__6868),
            .I(N__6859));
    LocalMux I__1277 (
            .O(N__6865),
            .I(N__6856));
    LocalMux I__1276 (
            .O(N__6862),
            .I(N__6850));
    LocalMux I__1275 (
            .O(N__6859),
            .I(N__6850));
    Span4Mux_h I__1274 (
            .O(N__6856),
            .I(N__6847));
    InMux I__1273 (
            .O(N__6855),
            .I(N__6844));
    Span4Mux_h I__1272 (
            .O(N__6850),
            .I(N__6841));
    Odrv4 I__1271 (
            .O(N__6847),
            .I(\U712_CHIP_RAM.N_342 ));
    LocalMux I__1270 (
            .O(N__6844),
            .I(\U712_CHIP_RAM.N_342 ));
    Odrv4 I__1269 (
            .O(N__6841),
            .I(\U712_CHIP_RAM.N_342 ));
    CascadeMux I__1268 (
            .O(N__6834),
            .I(\U712_CHIP_RAM.N_293_cascade_ ));
    InMux I__1267 (
            .O(N__6831),
            .I(N__6828));
    LocalMux I__1266 (
            .O(N__6828),
            .I(\U712_CHIP_RAM.N_294 ));
    CascadeMux I__1265 (
            .O(N__6825),
            .I(N__6820));
    InMux I__1264 (
            .O(N__6824),
            .I(N__6817));
    InMux I__1263 (
            .O(N__6823),
            .I(N__6814));
    InMux I__1262 (
            .O(N__6820),
            .I(N__6811));
    LocalMux I__1261 (
            .O(N__6817),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1260 (
            .O(N__6814),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1259 (
            .O(N__6811),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    InMux I__1258 (
            .O(N__6804),
            .I(N__6801));
    LocalMux I__1257 (
            .O(N__6801),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3 ));
    InMux I__1256 (
            .O(N__6798),
            .I(N__6795));
    LocalMux I__1255 (
            .O(N__6795),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2 ));
    CascadeMux I__1254 (
            .O(N__6792),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    CascadeMux I__1253 (
            .O(N__6789),
            .I(N__6783));
    InMux I__1252 (
            .O(N__6788),
            .I(N__6779));
    InMux I__1251 (
            .O(N__6787),
            .I(N__6776));
    InMux I__1250 (
            .O(N__6786),
            .I(N__6773));
    InMux I__1249 (
            .O(N__6783),
            .I(N__6768));
    InMux I__1248 (
            .O(N__6782),
            .I(N__6768));
    LocalMux I__1247 (
            .O(N__6779),
            .I(N__6763));
    LocalMux I__1246 (
            .O(N__6776),
            .I(N__6763));
    LocalMux I__1245 (
            .O(N__6773),
            .I(N__6760));
    LocalMux I__1244 (
            .O(N__6768),
            .I(N__6757));
    Span4Mux_v I__1243 (
            .O(N__6763),
            .I(N__6752));
    Span4Mux_h I__1242 (
            .O(N__6760),
            .I(N__6752));
    Span4Mux_v I__1241 (
            .O(N__6757),
            .I(N__6749));
    Odrv4 I__1240 (
            .O(N__6752),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1239 (
            .O(N__6749),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1238 (
            .O(N__6744),
            .I(N__6741));
    LocalMux I__1237 (
            .O(N__6741),
            .I(N__6738));
    Odrv4 I__1236 (
            .O(N__6738),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0 ));
    InMux I__1235 (
            .O(N__6735),
            .I(N__6725));
    InMux I__1234 (
            .O(N__6734),
            .I(N__6725));
    InMux I__1233 (
            .O(N__6733),
            .I(N__6719));
    InMux I__1232 (
            .O(N__6732),
            .I(N__6719));
    InMux I__1231 (
            .O(N__6731),
            .I(N__6714));
    InMux I__1230 (
            .O(N__6730),
            .I(N__6714));
    LocalMux I__1229 (
            .O(N__6725),
            .I(N__6711));
    InMux I__1228 (
            .O(N__6724),
            .I(N__6708));
    LocalMux I__1227 (
            .O(N__6719),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1226 (
            .O(N__6714),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__1225 (
            .O(N__6711),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1224 (
            .O(N__6708),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__1223 (
            .O(N__6699),
            .I(N__6694));
    InMux I__1222 (
            .O(N__6698),
            .I(N__6691));
    InMux I__1221 (
            .O(N__6697),
            .I(N__6688));
    LocalMux I__1220 (
            .O(N__6694),
            .I(\U712_CHIP_RAM.N_207 ));
    LocalMux I__1219 (
            .O(N__6691),
            .I(\U712_CHIP_RAM.N_207 ));
    LocalMux I__1218 (
            .O(N__6688),
            .I(\U712_CHIP_RAM.N_207 ));
    InMux I__1217 (
            .O(N__6681),
            .I(N__6676));
    CascadeMux I__1216 (
            .O(N__6680),
            .I(N__6670));
    InMux I__1215 (
            .O(N__6679),
            .I(N__6667));
    LocalMux I__1214 (
            .O(N__6676),
            .I(N__6663));
    InMux I__1213 (
            .O(N__6675),
            .I(N__6655));
    InMux I__1212 (
            .O(N__6674),
            .I(N__6652));
    InMux I__1211 (
            .O(N__6673),
            .I(N__6649));
    InMux I__1210 (
            .O(N__6670),
            .I(N__6646));
    LocalMux I__1209 (
            .O(N__6667),
            .I(N__6643));
    InMux I__1208 (
            .O(N__6666),
            .I(N__6640));
    Span4Mux_h I__1207 (
            .O(N__6663),
            .I(N__6637));
    InMux I__1206 (
            .O(N__6662),
            .I(N__6634));
    InMux I__1205 (
            .O(N__6661),
            .I(N__6629));
    InMux I__1204 (
            .O(N__6660),
            .I(N__6629));
    InMux I__1203 (
            .O(N__6659),
            .I(N__6624));
    InMux I__1202 (
            .O(N__6658),
            .I(N__6624));
    LocalMux I__1201 (
            .O(N__6655),
            .I(N__6615));
    LocalMux I__1200 (
            .O(N__6652),
            .I(N__6615));
    LocalMux I__1199 (
            .O(N__6649),
            .I(N__6615));
    LocalMux I__1198 (
            .O(N__6646),
            .I(N__6615));
    Odrv4 I__1197 (
            .O(N__6643),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1196 (
            .O(N__6640),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1195 (
            .O(N__6637),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1194 (
            .O(N__6634),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1193 (
            .O(N__6629),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1192 (
            .O(N__6624),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1191 (
            .O(N__6615),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1190 (
            .O(N__6600),
            .I(N__6595));
    CascadeMux I__1189 (
            .O(N__6599),
            .I(N__6592));
    InMux I__1188 (
            .O(N__6598),
            .I(N__6587));
    InMux I__1187 (
            .O(N__6595),
            .I(N__6584));
    InMux I__1186 (
            .O(N__6592),
            .I(N__6576));
    InMux I__1185 (
            .O(N__6591),
            .I(N__6576));
    InMux I__1184 (
            .O(N__6590),
            .I(N__6576));
    LocalMux I__1183 (
            .O(N__6587),
            .I(N__6572));
    LocalMux I__1182 (
            .O(N__6584),
            .I(N__6569));
    CascadeMux I__1181 (
            .O(N__6583),
            .I(N__6566));
    LocalMux I__1180 (
            .O(N__6576),
            .I(N__6560));
    InMux I__1179 (
            .O(N__6575),
            .I(N__6557));
    Span4Mux_v I__1178 (
            .O(N__6572),
            .I(N__6552));
    Span4Mux_v I__1177 (
            .O(N__6569),
            .I(N__6552));
    InMux I__1176 (
            .O(N__6566),
            .I(N__6547));
    InMux I__1175 (
            .O(N__6565),
            .I(N__6547));
    InMux I__1174 (
            .O(N__6564),
            .I(N__6542));
    InMux I__1173 (
            .O(N__6563),
            .I(N__6542));
    Span4Mux_h I__1172 (
            .O(N__6560),
            .I(N__6539));
    LocalMux I__1171 (
            .O(N__6557),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1170 (
            .O(N__6552),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1169 (
            .O(N__6547),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1168 (
            .O(N__6542),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1167 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1166 (
            .O(N__6528),
            .I(N__6525));
    LocalMux I__1165 (
            .O(N__6525),
            .I(\U712_CHIP_RAM.N_262 ));
    CascadeMux I__1164 (
            .O(N__6522),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_ ));
    InMux I__1163 (
            .O(N__6519),
            .I(N__6516));
    LocalMux I__1162 (
            .O(N__6516),
            .I(N__6513));
    Odrv4 I__1161 (
            .O(N__6513),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0 ));
    CascadeMux I__1160 (
            .O(N__6510),
            .I(N__6507));
    InMux I__1159 (
            .O(N__6507),
            .I(N__6504));
    LocalMux I__1158 (
            .O(N__6504),
            .I(\U712_CHIP_RAM.N_237 ));
    CascadeMux I__1157 (
            .O(N__6501),
            .I(N__6497));
    CascadeMux I__1156 (
            .O(N__6500),
            .I(N__6493));
    InMux I__1155 (
            .O(N__6497),
            .I(N__6487));
    InMux I__1154 (
            .O(N__6496),
            .I(N__6482));
    InMux I__1153 (
            .O(N__6493),
            .I(N__6482));
    InMux I__1152 (
            .O(N__6492),
            .I(N__6476));
    InMux I__1151 (
            .O(N__6491),
            .I(N__6471));
    InMux I__1150 (
            .O(N__6490),
            .I(N__6471));
    LocalMux I__1149 (
            .O(N__6487),
            .I(N__6465));
    LocalMux I__1148 (
            .O(N__6482),
            .I(N__6465));
    InMux I__1147 (
            .O(N__6481),
            .I(N__6460));
    InMux I__1146 (
            .O(N__6480),
            .I(N__6457));
    InMux I__1145 (
            .O(N__6479),
            .I(N__6454));
    LocalMux I__1144 (
            .O(N__6476),
            .I(N__6451));
    LocalMux I__1143 (
            .O(N__6471),
            .I(N__6448));
    InMux I__1142 (
            .O(N__6470),
            .I(N__6445));
    Span4Mux_h I__1141 (
            .O(N__6465),
            .I(N__6442));
    InMux I__1140 (
            .O(N__6464),
            .I(N__6439));
    InMux I__1139 (
            .O(N__6463),
            .I(N__6436));
    LocalMux I__1138 (
            .O(N__6460),
            .I(N__6431));
    LocalMux I__1137 (
            .O(N__6457),
            .I(N__6431));
    LocalMux I__1136 (
            .O(N__6454),
            .I(N__6428));
    Span4Mux_h I__1135 (
            .O(N__6451),
            .I(N__6423));
    Span4Mux_v I__1134 (
            .O(N__6448),
            .I(N__6423));
    LocalMux I__1133 (
            .O(N__6445),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1132 (
            .O(N__6442),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1131 (
            .O(N__6439),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1130 (
            .O(N__6436),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1129 (
            .O(N__6431),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1128 (
            .O(N__6428),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1127 (
            .O(N__6423),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1126 (
            .O(N__6408),
            .I(N__6405));
    LocalMux I__1125 (
            .O(N__6405),
            .I(N__6402));
    Span4Mux_v I__1124 (
            .O(N__6402),
            .I(N__6399));
    Span4Mux_h I__1123 (
            .O(N__6399),
            .I(N__6396));
    Span4Mux_h I__1122 (
            .O(N__6396),
            .I(N__6393));
    Sp12to4 I__1121 (
            .O(N__6393),
            .I(N__6390));
    Odrv12 I__1120 (
            .O(N__6390),
            .I(A_c_4));
    InMux I__1119 (
            .O(N__6387),
            .I(N__6384));
    LocalMux I__1118 (
            .O(N__6384),
            .I(N__6381));
    Span12Mux_v I__1117 (
            .O(N__6381),
            .I(N__6378));
    Span12Mux_h I__1116 (
            .O(N__6378),
            .I(N__6375));
    Odrv12 I__1115 (
            .O(N__6375),
            .I(A_c_11));
    CascadeMux I__1114 (
            .O(N__6372),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    CascadeMux I__1113 (
            .O(N__6369),
            .I(N__6365));
    CascadeMux I__1112 (
            .O(N__6368),
            .I(N__6356));
    InMux I__1111 (
            .O(N__6365),
            .I(N__6352));
    InMux I__1110 (
            .O(N__6364),
            .I(N__6347));
    InMux I__1109 (
            .O(N__6363),
            .I(N__6347));
    InMux I__1108 (
            .O(N__6362),
            .I(N__6344));
    InMux I__1107 (
            .O(N__6361),
            .I(N__6339));
    CascadeMux I__1106 (
            .O(N__6360),
            .I(N__6336));
    InMux I__1105 (
            .O(N__6359),
            .I(N__6333));
    InMux I__1104 (
            .O(N__6356),
            .I(N__6328));
    InMux I__1103 (
            .O(N__6355),
            .I(N__6325));
    LocalMux I__1102 (
            .O(N__6352),
            .I(N__6318));
    LocalMux I__1101 (
            .O(N__6347),
            .I(N__6318));
    LocalMux I__1100 (
            .O(N__6344),
            .I(N__6318));
    InMux I__1099 (
            .O(N__6343),
            .I(N__6315));
    InMux I__1098 (
            .O(N__6342),
            .I(N__6312));
    LocalMux I__1097 (
            .O(N__6339),
            .I(N__6309));
    InMux I__1096 (
            .O(N__6336),
            .I(N__6306));
    LocalMux I__1095 (
            .O(N__6333),
            .I(N__6303));
    InMux I__1094 (
            .O(N__6332),
            .I(N__6298));
    InMux I__1093 (
            .O(N__6331),
            .I(N__6298));
    LocalMux I__1092 (
            .O(N__6328),
            .I(N__6295));
    LocalMux I__1091 (
            .O(N__6325),
            .I(N__6290));
    Span4Mux_v I__1090 (
            .O(N__6318),
            .I(N__6290));
    LocalMux I__1089 (
            .O(N__6315),
            .I(N__6287));
    LocalMux I__1088 (
            .O(N__6312),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1087 (
            .O(N__6309),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1086 (
            .O(N__6306),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1085 (
            .O(N__6303),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1084 (
            .O(N__6298),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1083 (
            .O(N__6295),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1082 (
            .O(N__6290),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1081 (
            .O(N__6287),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1080 (
            .O(N__6270),
            .I(N__6267));
    LocalMux I__1079 (
            .O(N__6267),
            .I(N__6264));
    Span4Mux_v I__1078 (
            .O(N__6264),
            .I(N__6260));
    InMux I__1077 (
            .O(N__6263),
            .I(N__6257));
    Odrv4 I__1076 (
            .O(N__6260),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0 ));
    LocalMux I__1075 (
            .O(N__6257),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0 ));
    CascadeMux I__1074 (
            .O(N__6252),
            .I(N__6249));
    InMux I__1073 (
            .O(N__6249),
            .I(N__6243));
    InMux I__1072 (
            .O(N__6248),
            .I(N__6240));
    InMux I__1071 (
            .O(N__6247),
            .I(N__6237));
    CascadeMux I__1070 (
            .O(N__6246),
            .I(N__6229));
    LocalMux I__1069 (
            .O(N__6243),
            .I(N__6226));
    LocalMux I__1068 (
            .O(N__6240),
            .I(N__6221));
    LocalMux I__1067 (
            .O(N__6237),
            .I(N__6221));
    InMux I__1066 (
            .O(N__6236),
            .I(N__6218));
    InMux I__1065 (
            .O(N__6235),
            .I(N__6215));
    InMux I__1064 (
            .O(N__6234),
            .I(N__6210));
    InMux I__1063 (
            .O(N__6233),
            .I(N__6210));
    InMux I__1062 (
            .O(N__6232),
            .I(N__6207));
    InMux I__1061 (
            .O(N__6229),
            .I(N__6204));
    Span4Mux_h I__1060 (
            .O(N__6226),
            .I(N__6199));
    Span4Mux_h I__1059 (
            .O(N__6221),
            .I(N__6199));
    LocalMux I__1058 (
            .O(N__6218),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__1057 (
            .O(N__6215),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__1056 (
            .O(N__6210),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__1055 (
            .O(N__6207),
            .I(\U712_CHIP_RAM.N_335 ));
    LocalMux I__1054 (
            .O(N__6204),
            .I(\U712_CHIP_RAM.N_335 ));
    Odrv4 I__1053 (
            .O(N__6199),
            .I(\U712_CHIP_RAM.N_335 ));
    CascadeMux I__1052 (
            .O(N__6186),
            .I(N__6182));
    InMux I__1051 (
            .O(N__6185),
            .I(N__6179));
    InMux I__1050 (
            .O(N__6182),
            .I(N__6176));
    LocalMux I__1049 (
            .O(N__6179),
            .I(\U712_CHIP_RAM.N_261 ));
    LocalMux I__1048 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.N_261 ));
    InMux I__1047 (
            .O(N__6171),
            .I(N__6167));
    InMux I__1046 (
            .O(N__6170),
            .I(N__6163));
    LocalMux I__1045 (
            .O(N__6167),
            .I(N__6156));
    InMux I__1044 (
            .O(N__6166),
            .I(N__6153));
    LocalMux I__1043 (
            .O(N__6163),
            .I(N__6149));
    InMux I__1042 (
            .O(N__6162),
            .I(N__6146));
    CascadeMux I__1041 (
            .O(N__6161),
            .I(N__6137));
    InMux I__1040 (
            .O(N__6160),
            .I(N__6131));
    InMux I__1039 (
            .O(N__6159),
            .I(N__6128));
    Span4Mux_v I__1038 (
            .O(N__6156),
            .I(N__6123));
    LocalMux I__1037 (
            .O(N__6153),
            .I(N__6123));
    InMux I__1036 (
            .O(N__6152),
            .I(N__6120));
    Span4Mux_h I__1035 (
            .O(N__6149),
            .I(N__6115));
    LocalMux I__1034 (
            .O(N__6146),
            .I(N__6115));
    InMux I__1033 (
            .O(N__6145),
            .I(N__6110));
    InMux I__1032 (
            .O(N__6144),
            .I(N__6110));
    InMux I__1031 (
            .O(N__6143),
            .I(N__6103));
    InMux I__1030 (
            .O(N__6142),
            .I(N__6103));
    InMux I__1029 (
            .O(N__6141),
            .I(N__6103));
    InMux I__1028 (
            .O(N__6140),
            .I(N__6098));
    InMux I__1027 (
            .O(N__6137),
            .I(N__6098));
    InMux I__1026 (
            .O(N__6136),
            .I(N__6095));
    InMux I__1025 (
            .O(N__6135),
            .I(N__6090));
    InMux I__1024 (
            .O(N__6134),
            .I(N__6090));
    LocalMux I__1023 (
            .O(N__6131),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1022 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.N_180 ));
    Odrv4 I__1021 (
            .O(N__6123),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1020 (
            .O(N__6120),
            .I(\U712_CHIP_RAM.N_180 ));
    Odrv4 I__1019 (
            .O(N__6115),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1018 (
            .O(N__6110),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1017 (
            .O(N__6103),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1016 (
            .O(N__6098),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1015 (
            .O(N__6095),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1014 (
            .O(N__6090),
            .I(\U712_CHIP_RAM.N_180 ));
    InMux I__1013 (
            .O(N__6069),
            .I(N__6066));
    LocalMux I__1012 (
            .O(N__6066),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0 ));
    CascadeMux I__1011 (
            .O(N__6063),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_ ));
    InMux I__1010 (
            .O(N__6060),
            .I(N__6057));
    LocalMux I__1009 (
            .O(N__6057),
            .I(\U712_BYTE_ENABLE.N_319 ));
    CascadeMux I__1008 (
            .O(N__6054),
            .I(N__6048));
    InMux I__1007 (
            .O(N__6053),
            .I(N__6042));
    InMux I__1006 (
            .O(N__6052),
            .I(N__6042));
    InMux I__1005 (
            .O(N__6051),
            .I(N__6038));
    InMux I__1004 (
            .O(N__6048),
            .I(N__6033));
    InMux I__1003 (
            .O(N__6047),
            .I(N__6033));
    LocalMux I__1002 (
            .O(N__6042),
            .I(N__6030));
    InMux I__1001 (
            .O(N__6041),
            .I(N__6027));
    LocalMux I__1000 (
            .O(N__6038),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__999 (
            .O(N__6033),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    Odrv4 I__998 (
            .O(N__6030),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__997 (
            .O(N__6027),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    InMux I__996 (
            .O(N__6018),
            .I(N__6015));
    LocalMux I__995 (
            .O(N__6015),
            .I(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0 ));
    InMux I__994 (
            .O(N__6012),
            .I(N__6009));
    LocalMux I__993 (
            .O(N__6009),
            .I(\U712_REG_SM.N_26 ));
    CascadeMux I__992 (
            .O(N__6006),
            .I(N__6003));
    InMux I__991 (
            .O(N__6003),
            .I(N__6000));
    LocalMux I__990 (
            .O(N__6000),
            .I(\U712_REG_SM.N_274 ));
    IoInMux I__989 (
            .O(N__5997),
            .I(N__5994));
    LocalMux I__988 (
            .O(N__5994),
            .I(N__5991));
    IoSpan4Mux I__987 (
            .O(N__5991),
            .I(N__5988));
    Span4Mux_s2_v I__986 (
            .O(N__5988),
            .I(N__5985));
    Span4Mux_v I__985 (
            .O(N__5985),
            .I(N__5982));
    Span4Mux_h I__984 (
            .O(N__5982),
            .I(N__5979));
    Odrv4 I__983 (
            .O(N__5979),
            .I(DMA_LATCH_EN_c));
    IoInMux I__982 (
            .O(N__5976),
            .I(N__5973));
    LocalMux I__981 (
            .O(N__5973),
            .I(N__5970));
    Span12Mux_s6_v I__980 (
            .O(N__5970),
            .I(N__5967));
    Odrv12 I__979 (
            .O(N__5967),
            .I(CONSTANT_ONE_NET));
    InMux I__978 (
            .O(N__5964),
            .I(N__5961));
    LocalMux I__977 (
            .O(N__5961),
            .I(N__5958));
    Span12Mux_v I__976 (
            .O(N__5958),
            .I(N__5955));
    Span12Mux_h I__975 (
            .O(N__5955),
            .I(N__5952));
    Odrv12 I__974 (
            .O(N__5952),
            .I(A_c_15));
    InMux I__973 (
            .O(N__5949),
            .I(N__5946));
    LocalMux I__972 (
            .O(N__5946),
            .I(N__5943));
    Span4Mux_v I__971 (
            .O(N__5943),
            .I(N__5940));
    Sp12to4 I__970 (
            .O(N__5940),
            .I(N__5937));
    Span12Mux_h I__969 (
            .O(N__5937),
            .I(N__5934));
    Odrv12 I__968 (
            .O(N__5934),
            .I(A_c_8));
    InMux I__967 (
            .O(N__5931),
            .I(N__5928));
    LocalMux I__966 (
            .O(N__5928),
            .I(N__5925));
    Span12Mux_v I__965 (
            .O(N__5925),
            .I(N__5922));
    Span12Mux_h I__964 (
            .O(N__5922),
            .I(N__5919));
    Odrv12 I__963 (
            .O(N__5919),
            .I(A_c_2));
    InMux I__962 (
            .O(N__5916),
            .I(N__5913));
    LocalMux I__961 (
            .O(N__5913),
            .I(N__5910));
    Span12Mux_h I__960 (
            .O(N__5910),
            .I(N__5907));
    Odrv12 I__959 (
            .O(N__5907),
            .I(A_c_9));
    InMux I__958 (
            .O(N__5904),
            .I(N__5901));
    LocalMux I__957 (
            .O(N__5901),
            .I(N__5898));
    Span4Mux_v I__956 (
            .O(N__5898),
            .I(N__5895));
    Odrv4 I__955 (
            .O(N__5895),
            .I(\U712_REG_SM.N_383 ));
    CascadeMux I__954 (
            .O(N__5892),
            .I(\U712_REG_SM.N_383_cascade_ ));
    InMux I__953 (
            .O(N__5889),
            .I(N__5885));
    InMux I__952 (
            .O(N__5888),
            .I(N__5873));
    LocalMux I__951 (
            .O(N__5885),
            .I(N__5870));
    InMux I__950 (
            .O(N__5884),
            .I(N__5867));
    InMux I__949 (
            .O(N__5883),
            .I(N__5864));
    InMux I__948 (
            .O(N__5882),
            .I(N__5861));
    InMux I__947 (
            .O(N__5881),
            .I(N__5858));
    InMux I__946 (
            .O(N__5880),
            .I(N__5853));
    InMux I__945 (
            .O(N__5879),
            .I(N__5853));
    InMux I__944 (
            .O(N__5878),
            .I(N__5846));
    InMux I__943 (
            .O(N__5877),
            .I(N__5846));
    InMux I__942 (
            .O(N__5876),
            .I(N__5846));
    LocalMux I__941 (
            .O(N__5873),
            .I(N__5843));
    Odrv4 I__940 (
            .O(N__5870),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__939 (
            .O(N__5867),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__938 (
            .O(N__5864),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__937 (
            .O(N__5861),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__936 (
            .O(N__5858),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__935 (
            .O(N__5853),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__934 (
            .O(N__5846),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__933 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__932 (
            .O(N__5826),
            .I(\U712_CYCLE_TERM.N_321_cascade_ ));
    CascadeMux I__931 (
            .O(N__5823),
            .I(N__5820));
    InMux I__930 (
            .O(N__5820),
            .I(N__5816));
    InMux I__929 (
            .O(N__5819),
            .I(N__5813));
    LocalMux I__928 (
            .O(N__5816),
            .I(N__5808));
    LocalMux I__927 (
            .O(N__5813),
            .I(N__5808));
    Odrv12 I__926 (
            .O(N__5808),
            .I(CPU_TACKm));
    IoInMux I__925 (
            .O(N__5805),
            .I(N__5802));
    LocalMux I__924 (
            .O(N__5802),
            .I(N__5799));
    IoSpan4Mux I__923 (
            .O(N__5799),
            .I(N__5796));
    Sp12to4 I__922 (
            .O(N__5796),
            .I(N__5793));
    Span12Mux_s7_v I__921 (
            .O(N__5793),
            .I(N__5790));
    Span12Mux_v I__920 (
            .O(N__5790),
            .I(N__5787));
    Odrv12 I__919 (
            .O(N__5787),
            .I(N_156_i));
    InMux I__918 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__917 (
            .O(N__5781),
            .I(N__5777));
    InMux I__916 (
            .O(N__5780),
            .I(N__5774));
    Odrv12 I__915 (
            .O(N__5777),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0 ));
    LocalMux I__914 (
            .O(N__5774),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0 ));
    IoInMux I__913 (
            .O(N__5769),
            .I(N__5766));
    LocalMux I__912 (
            .O(N__5766),
            .I(N__5763));
    Span12Mux_s5_h I__911 (
            .O(N__5763),
            .I(N__5760));
    Span12Mux_h I__910 (
            .O(N__5760),
            .I(N__5757));
    Span12Mux_v I__909 (
            .O(N__5757),
            .I(N__5754));
    Odrv12 I__908 (
            .O(N__5754),
            .I(N_126_i));
    CascadeMux I__907 (
            .O(N__5751),
            .I(N__5748));
    InMux I__906 (
            .O(N__5748),
            .I(N__5742));
    InMux I__905 (
            .O(N__5747),
            .I(N__5742));
    LocalMux I__904 (
            .O(N__5742),
            .I(\U712_BYTE_ENABLE.N_315 ));
    CascadeMux I__903 (
            .O(N__5739),
            .I(\U712_CHIP_RAM.N_184_cascade_ ));
    InMux I__902 (
            .O(N__5736),
            .I(N__5733));
    LocalMux I__901 (
            .O(N__5733),
            .I(N__5730));
    Odrv4 I__900 (
            .O(N__5730),
            .I(\U712_CHIP_RAM.N_304 ));
    InMux I__899 (
            .O(N__5727),
            .I(N__5724));
    LocalMux I__898 (
            .O(N__5724),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0 ));
    CascadeMux I__897 (
            .O(N__5721),
            .I(\U712_CHIP_RAM.N_392_cascade_ ));
    CEMux I__896 (
            .O(N__5718),
            .I(N__5714));
    CEMux I__895 (
            .O(N__5717),
            .I(N__5710));
    LocalMux I__894 (
            .O(N__5714),
            .I(N__5707));
    CEMux I__893 (
            .O(N__5713),
            .I(N__5704));
    LocalMux I__892 (
            .O(N__5710),
            .I(N__5701));
    Span4Mux_h I__891 (
            .O(N__5707),
            .I(N__5696));
    LocalMux I__890 (
            .O(N__5704),
            .I(N__5696));
    Sp12to4 I__889 (
            .O(N__5701),
            .I(N__5693));
    Sp12to4 I__888 (
            .O(N__5696),
            .I(N__5690));
    Odrv12 I__887 (
            .O(N__5693),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv12 I__886 (
            .O(N__5690),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__885 (
            .O(N__5685),
            .I(N__5682));
    LocalMux I__884 (
            .O(N__5682),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0 ));
    CascadeMux I__883 (
            .O(N__5679),
            .I(N__5676));
    InMux I__882 (
            .O(N__5676),
            .I(N__5672));
    InMux I__881 (
            .O(N__5675),
            .I(N__5669));
    LocalMux I__880 (
            .O(N__5672),
            .I(N__5664));
    LocalMux I__879 (
            .O(N__5669),
            .I(N__5664));
    Odrv4 I__878 (
            .O(N__5664),
            .I(\U712_REG_SM.N_196 ));
    CascadeMux I__877 (
            .O(N__5661),
            .I(N__5656));
    InMux I__876 (
            .O(N__5660),
            .I(N__5653));
    InMux I__875 (
            .O(N__5659),
            .I(N__5650));
    InMux I__874 (
            .O(N__5656),
            .I(N__5647));
    LocalMux I__873 (
            .O(N__5653),
            .I(\U712_CHIP_RAM.N_333 ));
    LocalMux I__872 (
            .O(N__5650),
            .I(\U712_CHIP_RAM.N_333 ));
    LocalMux I__871 (
            .O(N__5647),
            .I(\U712_CHIP_RAM.N_333 ));
    CascadeMux I__870 (
            .O(N__5640),
            .I(\U712_CHIP_RAM.N_310_cascade_ ));
    CascadeMux I__869 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ));
    CEMux I__868 (
            .O(N__5634),
            .I(N__5631));
    LocalMux I__867 (
            .O(N__5631),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ));
    InMux I__866 (
            .O(N__5628),
            .I(N__5624));
    InMux I__865 (
            .O(N__5627),
            .I(N__5620));
    LocalMux I__864 (
            .O(N__5624),
            .I(N__5617));
    InMux I__863 (
            .O(N__5623),
            .I(N__5614));
    LocalMux I__862 (
            .O(N__5620),
            .I(N__5606));
    Span4Mux_v I__861 (
            .O(N__5617),
            .I(N__5606));
    LocalMux I__860 (
            .O(N__5614),
            .I(N__5606));
    InMux I__859 (
            .O(N__5613),
            .I(N__5603));
    Span4Mux_h I__858 (
            .O(N__5606),
            .I(N__5599));
    LocalMux I__857 (
            .O(N__5603),
            .I(N__5596));
    InMux I__856 (
            .O(N__5602),
            .I(N__5593));
    Odrv4 I__855 (
            .O(N__5599),
            .I(DMA_CYCLEm));
    Odrv4 I__854 (
            .O(N__5596),
            .I(DMA_CYCLEm));
    LocalMux I__853 (
            .O(N__5593),
            .I(DMA_CYCLEm));
    IoInMux I__852 (
            .O(N__5586),
            .I(N__5583));
    LocalMux I__851 (
            .O(N__5583),
            .I(N__5580));
    Span4Mux_s3_v I__850 (
            .O(N__5580),
            .I(N__5575));
    InMux I__849 (
            .O(N__5579),
            .I(N__5572));
    InMux I__848 (
            .O(N__5578),
            .I(N__5569));
    Span4Mux_h I__847 (
            .O(N__5575),
            .I(N__5566));
    LocalMux I__846 (
            .O(N__5572),
            .I(N__5563));
    LocalMux I__845 (
            .O(N__5569),
            .I(N__5560));
    Sp12to4 I__844 (
            .O(N__5566),
            .I(N__5556));
    Span4Mux_v I__843 (
            .O(N__5563),
            .I(N__5553));
    Span4Mux_h I__842 (
            .O(N__5560),
            .I(N__5550));
    InMux I__841 (
            .O(N__5559),
            .I(N__5547));
    Odrv12 I__840 (
            .O(N__5556),
            .I(DBENn_c));
    Odrv4 I__839 (
            .O(N__5553),
            .I(DBENn_c));
    Odrv4 I__838 (
            .O(N__5550),
            .I(DBENn_c));
    LocalMux I__837 (
            .O(N__5547),
            .I(DBENn_c));
    InMux I__836 (
            .O(N__5538),
            .I(N__5535));
    LocalMux I__835 (
            .O(N__5535),
            .I(N__5531));
    InMux I__834 (
            .O(N__5534),
            .I(N__5528));
    Odrv4 I__833 (
            .O(N__5531),
            .I(\U712_CHIP_RAM.N_334 ));
    LocalMux I__832 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.N_334 ));
    InMux I__831 (
            .O(N__5523),
            .I(N__5520));
    LocalMux I__830 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.N_297 ));
    InMux I__829 (
            .O(N__5517),
            .I(N__5514));
    LocalMux I__828 (
            .O(N__5514),
            .I(N__5510));
    InMux I__827 (
            .O(N__5513),
            .I(N__5507));
    Span4Mux_v I__826 (
            .O(N__5510),
            .I(N__5502));
    LocalMux I__825 (
            .O(N__5507),
            .I(N__5502));
    Odrv4 I__824 (
            .O(N__5502),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0 ));
    InMux I__823 (
            .O(N__5499),
            .I(N__5495));
    InMux I__822 (
            .O(N__5498),
            .I(N__5492));
    LocalMux I__821 (
            .O(N__5495),
            .I(\U712_CHIP_RAM.N_202 ));
    LocalMux I__820 (
            .O(N__5492),
            .I(\U712_CHIP_RAM.N_202 ));
    InMux I__819 (
            .O(N__5487),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__818 (
            .O(N__5484),
            .I(N__5480));
    InMux I__817 (
            .O(N__5483),
            .I(N__5477));
    LocalMux I__816 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__815 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__814 (
            .O(N__5472),
            .I(N__5445));
    ClkMux I__813 (
            .O(N__5471),
            .I(N__5445));
    ClkMux I__812 (
            .O(N__5470),
            .I(N__5445));
    ClkMux I__811 (
            .O(N__5469),
            .I(N__5445));
    ClkMux I__810 (
            .O(N__5468),
            .I(N__5445));
    ClkMux I__809 (
            .O(N__5467),
            .I(N__5445));
    ClkMux I__808 (
            .O(N__5466),
            .I(N__5445));
    ClkMux I__807 (
            .O(N__5465),
            .I(N__5445));
    ClkMux I__806 (
            .O(N__5464),
            .I(N__5445));
    GlobalMux I__805 (
            .O(N__5445),
            .I(N__5442));
    gio2CtrlBuf I__804 (
            .O(N__5442),
            .I(C1_c_g));
    InMux I__803 (
            .O(N__5439),
            .I(N__5436));
    LocalMux I__802 (
            .O(N__5436),
            .I(\U712_CHIP_RAM.N_134 ));
    InMux I__801 (
            .O(N__5433),
            .I(N__5430));
    LocalMux I__800 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__799 (
            .O(N__5427),
            .I(N__5424));
    LocalMux I__798 (
            .O(N__5424),
            .I(N__5421));
    IoSpan4Mux I__797 (
            .O(N__5421),
            .I(N__5418));
    IoSpan4Mux I__796 (
            .O(N__5418),
            .I(N__5415));
    Span4Mux_s2_h I__795 (
            .O(N__5415),
            .I(N__5412));
    Sp12to4 I__794 (
            .O(N__5412),
            .I(N__5409));
    Span12Mux_s9_h I__793 (
            .O(N__5409),
            .I(N__5406));
    Odrv12 I__792 (
            .O(N__5406),
            .I(N_116_i));
    CascadeMux I__791 (
            .O(N__5403),
            .I(\U712_CHIP_RAM.N_207_cascade_ ));
    CascadeMux I__790 (
            .O(N__5400),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_ ));
    CascadeMux I__789 (
            .O(N__5397),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_ ));
    CascadeMux I__788 (
            .O(N__5394),
            .I(\U712_REG_SM.N_284_cascade_ ));
    InMux I__787 (
            .O(N__5391),
            .I(N__5387));
    InMux I__786 (
            .O(N__5390),
            .I(N__5384));
    LocalMux I__785 (
            .O(N__5387),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__784 (
            .O(N__5384),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__783 (
            .O(N__5379),
            .I(bfn_10_15_0_));
    InMux I__782 (
            .O(N__5376),
            .I(N__5372));
    InMux I__781 (
            .O(N__5375),
            .I(N__5369));
    LocalMux I__780 (
            .O(N__5372),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__779 (
            .O(N__5369),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__778 (
            .O(N__5364),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__777 (
            .O(N__5361),
            .I(N__5357));
    InMux I__776 (
            .O(N__5360),
            .I(N__5354));
    LocalMux I__775 (
            .O(N__5357),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__774 (
            .O(N__5354),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__773 (
            .O(N__5349),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__772 (
            .O(N__5346),
            .I(N__5342));
    InMux I__771 (
            .O(N__5345),
            .I(N__5339));
    LocalMux I__770 (
            .O(N__5342),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__769 (
            .O(N__5339),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__768 (
            .O(N__5334),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__767 (
            .O(N__5331),
            .I(N__5327));
    InMux I__766 (
            .O(N__5330),
            .I(N__5324));
    InMux I__765 (
            .O(N__5327),
            .I(N__5321));
    LocalMux I__764 (
            .O(N__5324),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__763 (
            .O(N__5321),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__762 (
            .O(N__5316),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__761 (
            .O(N__5313),
            .I(N__5309));
    InMux I__760 (
            .O(N__5312),
            .I(N__5306));
    LocalMux I__759 (
            .O(N__5309),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__758 (
            .O(N__5306),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__757 (
            .O(N__5301),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__756 (
            .O(N__5298),
            .I(N__5294));
    InMux I__755 (
            .O(N__5297),
            .I(N__5291));
    LocalMux I__754 (
            .O(N__5294),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__753 (
            .O(N__5291),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__752 (
            .O(N__5286),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__751 (
            .O(N__5283),
            .I(N__5280));
    LocalMux I__750 (
            .O(N__5280),
            .I(N__5277));
    Odrv4 I__749 (
            .O(N__5277),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18 ));
    InMux I__748 (
            .O(N__5274),
            .I(N__5264));
    InMux I__747 (
            .O(N__5273),
            .I(N__5264));
    InMux I__746 (
            .O(N__5272),
            .I(N__5264));
    InMux I__745 (
            .O(N__5271),
            .I(N__5261));
    LocalMux I__744 (
            .O(N__5264),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__743 (
            .O(N__5261),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__742 (
            .O(N__5256),
            .I(N__5253));
    LocalMux I__741 (
            .O(N__5253),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ));
    InMux I__740 (
            .O(N__5250),
            .I(N__5247));
    LocalMux I__739 (
            .O(N__5247),
            .I(\U712_REG_SM.N_222 ));
    CascadeMux I__738 (
            .O(N__5244),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ));
    CascadeMux I__737 (
            .O(N__5241),
            .I(N__5236));
    InMux I__736 (
            .O(N__5240),
            .I(N__5231));
    InMux I__735 (
            .O(N__5239),
            .I(N__5231));
    InMux I__734 (
            .O(N__5236),
            .I(N__5228));
    LocalMux I__733 (
            .O(N__5231),
            .I(N__5225));
    LocalMux I__732 (
            .O(N__5228),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__731 (
            .O(N__5225),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__730 (
            .O(N__5220),
            .I(N__5216));
    InMux I__729 (
            .O(N__5219),
            .I(N__5213));
    LocalMux I__728 (
            .O(N__5216),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    LocalMux I__727 (
            .O(N__5213),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__726 (
            .O(N__5208),
            .I(N__5205));
    LocalMux I__725 (
            .O(N__5205),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__724 (
            .O(N__5202),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__723 (
            .O(N__5199),
            .I(N__5195));
    InMux I__722 (
            .O(N__5198),
            .I(N__5192));
    LocalMux I__721 (
            .O(N__5195),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__720 (
            .O(N__5192),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__719 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__718 (
            .O(N__5184),
            .I(N__5180));
    InMux I__717 (
            .O(N__5183),
            .I(N__5177));
    LocalMux I__716 (
            .O(N__5180),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__715 (
            .O(N__5177),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__714 (
            .O(N__5172),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__713 (
            .O(N__5169),
            .I(N__5166));
    InMux I__712 (
            .O(N__5166),
            .I(N__5162));
    InMux I__711 (
            .O(N__5165),
            .I(N__5153));
    LocalMux I__710 (
            .O(N__5162),
            .I(N__5150));
    InMux I__709 (
            .O(N__5161),
            .I(N__5141));
    InMux I__708 (
            .O(N__5160),
            .I(N__5141));
    InMux I__707 (
            .O(N__5159),
            .I(N__5141));
    InMux I__706 (
            .O(N__5158),
            .I(N__5141));
    InMux I__705 (
            .O(N__5157),
            .I(N__5136));
    InMux I__704 (
            .O(N__5156),
            .I(N__5136));
    LocalMux I__703 (
            .O(N__5153),
            .I(N__5133));
    Odrv4 I__702 (
            .O(N__5150),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__701 (
            .O(N__5141),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__700 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.N_46 ));
    Odrv4 I__699 (
            .O(N__5133),
            .I(\U712_CHIP_RAM.N_46 ));
    InMux I__698 (
            .O(N__5124),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__697 (
            .O(N__5121),
            .I(N__5117));
    InMux I__696 (
            .O(N__5120),
            .I(N__5114));
    LocalMux I__695 (
            .O(N__5117),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__694 (
            .O(N__5114),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__693 (
            .O(N__5109),
            .I(N__5106));
    LocalMux I__692 (
            .O(N__5106),
            .I(\U712_CYCLE_TERM.N_217_i_0_en ));
    InMux I__691 (
            .O(N__5103),
            .I(N__5100));
    LocalMux I__690 (
            .O(N__5100),
            .I(\U712_REG_SM.START_RST_0_sqmuxa ));
    InMux I__689 (
            .O(N__5097),
            .I(N__5091));
    InMux I__688 (
            .O(N__5096),
            .I(N__5091));
    LocalMux I__687 (
            .O(N__5091),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    CascadeMux I__686 (
            .O(N__5088),
            .I(\U712_REG_SM.N_285_cascade_ ));
    CascadeMux I__685 (
            .O(N__5085),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ));
    InMux I__684 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__683 (
            .O(N__5079),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ));
    InMux I__682 (
            .O(N__5076),
            .I(N__5073));
    LocalMux I__681 (
            .O(N__5073),
            .I(\U712_CHIP_RAM.N_239 ));
    InMux I__680 (
            .O(N__5070),
            .I(N__5067));
    LocalMux I__679 (
            .O(N__5067),
            .I(\U712_CHIP_RAM.N_269 ));
    CascadeMux I__678 (
            .O(N__5064),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_ ));
    InMux I__677 (
            .O(N__5061),
            .I(N__5058));
    LocalMux I__676 (
            .O(N__5058),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__675 (
            .O(N__5055),
            .I(bfn_10_12_0_));
    InMux I__674 (
            .O(N__5052),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__673 (
            .O(N__5049),
            .I(N__5046));
    LocalMux I__672 (
            .O(N__5046),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__671 (
            .O(N__5043),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__670 (
            .O(N__5040),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__669 (
            .O(N__5037),
            .I(N__5034));
    LocalMux I__668 (
            .O(N__5034),
            .I(N__5031));
    Span4Mux_v I__667 (
            .O(N__5031),
            .I(N__5028));
    Odrv4 I__666 (
            .O(N__5028),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_3 ));
    CascadeMux I__665 (
            .O(N__5025),
            .I(N__5021));
    InMux I__664 (
            .O(N__5024),
            .I(N__5018));
    InMux I__663 (
            .O(N__5021),
            .I(N__5015));
    LocalMux I__662 (
            .O(N__5018),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    LocalMux I__661 (
            .O(N__5015),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    InMux I__660 (
            .O(N__5010),
            .I(N__5006));
    InMux I__659 (
            .O(N__5009),
            .I(N__5003));
    LocalMux I__658 (
            .O(N__5006),
            .I(N__5000));
    LocalMux I__657 (
            .O(N__5003),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__656 (
            .O(N__5000),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__655 (
            .O(N__4995),
            .I(N__4992));
    LocalMux I__654 (
            .O(N__4992),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__653 (
            .O(N__4989),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_ ));
    IoInMux I__652 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__651 (
            .O(N__4983),
            .I(N__4980));
    Span4Mux_s3_v I__650 (
            .O(N__4980),
            .I(N__4977));
    Span4Mux_v I__649 (
            .O(N__4977),
            .I(N__4974));
    Span4Mux_v I__648 (
            .O(N__4974),
            .I(N__4971));
    Span4Mux_v I__647 (
            .O(N__4971),
            .I(N__4967));
    InMux I__646 (
            .O(N__4970),
            .I(N__4964));
    Odrv4 I__645 (
            .O(N__4967),
            .I(BANK0_c));
    LocalMux I__644 (
            .O(N__4964),
            .I(BANK0_c));
    InMux I__643 (
            .O(N__4959),
            .I(N__4956));
    LocalMux I__642 (
            .O(N__4956),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_4 ));
    InMux I__641 (
            .O(N__4953),
            .I(N__4949));
    InMux I__640 (
            .O(N__4952),
            .I(N__4946));
    LocalMux I__639 (
            .O(N__4949),
            .I(\U712_CHIP_RAM.N_186 ));
    LocalMux I__638 (
            .O(N__4946),
            .I(\U712_CHIP_RAM.N_186 ));
    CascadeMux I__637 (
            .O(N__4941),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_ ));
    InMux I__636 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__635 (
            .O(N__4935),
            .I(\U712_CHIP_RAM.N_306 ));
    CascadeMux I__634 (
            .O(N__4932),
            .I(\U712_CHIP_RAM.N_333_cascade_ ));
    CascadeMux I__633 (
            .O(N__4929),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_ ));
    InMux I__632 (
            .O(N__4926),
            .I(N__4922));
    IoInMux I__631 (
            .O(N__4925),
            .I(N__4919));
    LocalMux I__630 (
            .O(N__4922),
            .I(N__4916));
    LocalMux I__629 (
            .O(N__4919),
            .I(N__4913));
    Span4Mux_v I__628 (
            .O(N__4916),
            .I(N__4910));
    IoSpan4Mux I__627 (
            .O(N__4913),
            .I(N__4907));
    Sp12to4 I__626 (
            .O(N__4910),
            .I(N__4904));
    IoSpan4Mux I__625 (
            .O(N__4907),
            .I(N__4901));
    Span12Mux_h I__624 (
            .O(N__4904),
            .I(N__4898));
    IoSpan4Mux I__623 (
            .O(N__4901),
            .I(N__4895));
    Odrv12 I__622 (
            .O(N__4898),
            .I(C1_c));
    Odrv4 I__621 (
            .O(N__4895),
            .I(C1_c));
    InMux I__620 (
            .O(N__4890),
            .I(N__4887));
    LocalMux I__619 (
            .O(N__4887),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__618 (
            .O(N__4884),
            .I(N__4880));
    InMux I__617 (
            .O(N__4883),
            .I(N__4877));
    LocalMux I__616 (
            .O(N__4880),
            .I(N__4874));
    LocalMux I__615 (
            .O(N__4877),
            .I(N__4871));
    Span4Mux_v I__614 (
            .O(N__4874),
            .I(N__4868));
    Span4Mux_h I__613 (
            .O(N__4871),
            .I(N__4865));
    Sp12to4 I__612 (
            .O(N__4868),
            .I(N__4862));
    Span4Mux_v I__611 (
            .O(N__4865),
            .I(N__4859));
    Span12Mux_h I__610 (
            .O(N__4862),
            .I(N__4856));
    IoSpan4Mux I__609 (
            .O(N__4859),
            .I(N__4853));
    Odrv12 I__608 (
            .O(N__4856),
            .I(TSn_c));
    Odrv4 I__607 (
            .O(N__4853),
            .I(TSn_c));
    InMux I__606 (
            .O(N__4848),
            .I(N__4845));
    LocalMux I__605 (
            .O(N__4845),
            .I(N__4842));
    Span4Mux_h I__604 (
            .O(N__4842),
            .I(N__4839));
    Span4Mux_v I__603 (
            .O(N__4839),
            .I(N__4836));
    Odrv4 I__602 (
            .O(N__4836),
            .I(RAMSPACEn_c));
    InMux I__601 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__600 (
            .O(N__4830),
            .I(N__4827));
    Span12Mux_v I__599 (
            .O(N__4827),
            .I(N__4824));
    Odrv12 I__598 (
            .O(N__4824),
            .I(\U712_CHIP_RAM.N_289 ));
    IoInMux I__597 (
            .O(N__4821),
            .I(N__4818));
    LocalMux I__596 (
            .O(N__4818),
            .I(N__4815));
    Span4Mux_s1_v I__595 (
            .O(N__4815),
            .I(N__4812));
    Span4Mux_v I__594 (
            .O(N__4812),
            .I(N__4809));
    Span4Mux_v I__593 (
            .O(N__4809),
            .I(N__4806));
    Span4Mux_v I__592 (
            .O(N__4806),
            .I(N__4803));
    Odrv4 I__591 (
            .O(N__4803),
            .I(CMA_c_1));
    InMux I__590 (
            .O(N__4800),
            .I(N__4797));
    LocalMux I__589 (
            .O(N__4797),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__588 (
            .O(N__4794),
            .I(N__4791));
    LocalMux I__587 (
            .O(N__4791),
            .I(N__4788));
    Span12Mux_v I__586 (
            .O(N__4788),
            .I(N__4785));
    Span12Mux_h I__585 (
            .O(N__4785),
            .I(N__4782));
    Odrv12 I__584 (
            .O(N__4782),
            .I(A_c_3));
    InMux I__583 (
            .O(N__4779),
            .I(N__4776));
    LocalMux I__582 (
            .O(N__4776),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    CascadeMux I__581 (
            .O(N__4773),
            .I(N__4770));
    InMux I__580 (
            .O(N__4770),
            .I(N__4764));
    InMux I__579 (
            .O(N__4769),
            .I(N__4764));
    LocalMux I__578 (
            .O(N__4764),
            .I(N__4761));
    Span12Mux_v I__577 (
            .O(N__4761),
            .I(N__4758));
    Span12Mux_h I__576 (
            .O(N__4758),
            .I(N__4755));
    Odrv12 I__575 (
            .O(N__4755),
            .I(A_c_10));
    InMux I__574 (
            .O(N__4752),
            .I(N__4749));
    LocalMux I__573 (
            .O(N__4749),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__572 (
            .O(N__4746),
            .I(N__4741));
    InMux I__571 (
            .O(N__4745),
            .I(N__4736));
    InMux I__570 (
            .O(N__4744),
            .I(N__4736));
    LocalMux I__569 (
            .O(N__4741),
            .I(\U712_CHIP_RAM.N_208 ));
    LocalMux I__568 (
            .O(N__4736),
            .I(\U712_CHIP_RAM.N_208 ));
    CEMux I__567 (
            .O(N__4731),
            .I(N__4728));
    LocalMux I__566 (
            .O(N__4728),
            .I(N__4725));
    Odrv4 I__565 (
            .O(N__4725),
            .I(\U712_CYCLE_TERM.N_217_i_0_en_0 ));
    IoInMux I__564 (
            .O(N__4722),
            .I(N__4719));
    LocalMux I__563 (
            .O(N__4719),
            .I(N__4715));
    IoInMux I__562 (
            .O(N__4718),
            .I(N__4712));
    Span12Mux_s1_v I__561 (
            .O(N__4715),
            .I(N__4709));
    LocalMux I__560 (
            .O(N__4712),
            .I(N__4706));
    Span12Mux_v I__559 (
            .O(N__4709),
            .I(N__4703));
    Span12Mux_s1_v I__558 (
            .O(N__4706),
            .I(N__4700));
    Span12Mux_h I__557 (
            .O(N__4703),
            .I(N__4694));
    Span12Mux_v I__556 (
            .O(N__4700),
            .I(N__4694));
    InMux I__555 (
            .O(N__4699),
            .I(N__4691));
    Odrv12 I__554 (
            .O(N__4694),
            .I(ASn_c));
    LocalMux I__553 (
            .O(N__4691),
            .I(ASn_c));
    InMux I__552 (
            .O(N__4686),
            .I(N__4682));
    InMux I__551 (
            .O(N__4685),
            .I(N__4679));
    LocalMux I__550 (
            .O(N__4682),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__549 (
            .O(N__4679),
            .I(\U712_REG_SM.START_RSTZ0 ));
    IoInMux I__548 (
            .O(N__4674),
            .I(N__4671));
    LocalMux I__547 (
            .O(N__4671),
            .I(N__4667));
    InMux I__546 (
            .O(N__4670),
            .I(N__4664));
    Span4Mux_s1_v I__545 (
            .O(N__4667),
            .I(N__4661));
    LocalMux I__544 (
            .O(N__4664),
            .I(N__4658));
    Sp12to4 I__543 (
            .O(N__4661),
            .I(N__4655));
    Span4Mux_v I__542 (
            .O(N__4658),
            .I(N__4652));
    Span12Mux_h I__541 (
            .O(N__4655),
            .I(N__4649));
    Sp12to4 I__540 (
            .O(N__4652),
            .I(N__4646));
    Span12Mux_v I__539 (
            .O(N__4649),
            .I(N__4641));
    Span12Mux_h I__538 (
            .O(N__4646),
            .I(N__4641));
    Span12Mux_v I__537 (
            .O(N__4641),
            .I(N__4638));
    Odrv12 I__536 (
            .O(N__4638),
            .I(RAMENn_c));
    CascadeMux I__535 (
            .O(N__4635),
            .I(\U712_REG_SM.N_270_cascade_ ));
    InMux I__534 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__533 (
            .O(N__4629),
            .I(N__4626));
    Odrv12 I__532 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_a2_2 ));
    CascadeMux I__531 (
            .O(N__4623),
            .I(N__4620));
    InMux I__530 (
            .O(N__4620),
            .I(N__4617));
    LocalMux I__529 (
            .O(N__4617),
            .I(N__4614));
    Odrv4 I__528 (
            .O(N__4614),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_a2_1 ));
    CascadeMux I__527 (
            .O(N__4611),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_cascade_ ));
    IoInMux I__526 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__525 (
            .O(N__4605),
            .I(N__4602));
    Span12Mux_s7_h I__524 (
            .O(N__4602),
            .I(N__4599));
    Span12Mux_h I__523 (
            .O(N__4599),
            .I(N__4595));
    InMux I__522 (
            .O(N__4598),
            .I(N__4592));
    Odrv12 I__521 (
            .O(N__4595),
            .I(CLK_EN_c));
    LocalMux I__520 (
            .O(N__4592),
            .I(CLK_EN_c));
    InMux I__519 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__518 (
            .O(N__4584),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ));
    InMux I__517 (
            .O(N__4581),
            .I(N__4578));
    LocalMux I__516 (
            .O(N__4578),
            .I(\U712_CHIP_RAM.N_385 ));
    CascadeMux I__515 (
            .O(N__4575),
            .I(\U712_CHIP_RAM.N_338_cascade_ ));
    CascadeMux I__514 (
            .O(N__4572),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    CascadeMux I__513 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.N_239_cascade_ ));
    CascadeMux I__512 (
            .O(N__4566),
            .I(N__4563));
    InMux I__511 (
            .O(N__4563),
            .I(N__4559));
    InMux I__510 (
            .O(N__4562),
            .I(N__4556));
    LocalMux I__509 (
            .O(N__4559),
            .I(N__4553));
    LocalMux I__508 (
            .O(N__4556),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    Odrv4 I__507 (
            .O(N__4553),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    InMux I__506 (
            .O(N__4548),
            .I(N__4543));
    InMux I__505 (
            .O(N__4547),
            .I(N__4540));
    InMux I__504 (
            .O(N__4546),
            .I(N__4537));
    LocalMux I__503 (
            .O(N__4543),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__502 (
            .O(N__4540),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    LocalMux I__501 (
            .O(N__4537),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    InMux I__500 (
            .O(N__4530),
            .I(N__4527));
    LocalMux I__499 (
            .O(N__4527),
            .I(\U712_CHIP_RAM.N_387 ));
    CascadeMux I__498 (
            .O(N__4524),
            .I(\U712_CHIP_RAM.N_385_cascade_ ));
    CascadeMux I__497 (
            .O(N__4521),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ));
    CascadeMux I__496 (
            .O(N__4518),
            .I(N__4515));
    InMux I__495 (
            .O(N__4515),
            .I(N__4512));
    LocalMux I__494 (
            .O(N__4512),
            .I(\U712_CHIP_RAM.N_223 ));
    CascadeMux I__493 (
            .O(N__4509),
            .I(\U712_CHIP_RAM.N_335_cascade_ ));
    CascadeMux I__492 (
            .O(N__4506),
            .I(\U712_CHIP_RAM.N_342_cascade_ ));
    InMux I__491 (
            .O(N__4503),
            .I(N__4500));
    LocalMux I__490 (
            .O(N__4500),
            .I(N__4497));
    Span4Mux_v I__489 (
            .O(N__4497),
            .I(N__4494));
    Span4Mux_h I__488 (
            .O(N__4494),
            .I(N__4491));
    Odrv4 I__487 (
            .O(N__4491),
            .I(TACK_EN_i_ess));
    IoInMux I__486 (
            .O(N__4488),
            .I(N__4485));
    LocalMux I__485 (
            .O(N__4485),
            .I(N__4482));
    IoSpan4Mux I__484 (
            .O(N__4482),
            .I(N__4479));
    Span4Mux_s0_h I__483 (
            .O(N__4479),
            .I(N__4476));
    Sp12to4 I__482 (
            .O(N__4476),
            .I(N__4473));
    Span12Mux_s11_h I__481 (
            .O(N__4473),
            .I(N__4469));
    InMux I__480 (
            .O(N__4472),
            .I(N__4466));
    Odrv12 I__479 (
            .O(N__4469),
            .I(TACK_OUTn));
    LocalMux I__478 (
            .O(N__4466),
            .I(TACK_OUTn));
    InMux I__477 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__476 (
            .O(N__4458),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__475 (
            .O(N__4455),
            .I(N__4452));
    LocalMux I__474 (
            .O(N__4452),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__473 (
            .O(N__4449),
            .I(N__4446));
    LocalMux I__472 (
            .O(N__4446),
            .I(N__4443));
    Span12Mux_s7_h I__471 (
            .O(N__4443),
            .I(N__4440));
    Span12Mux_h I__470 (
            .O(N__4440),
            .I(N__4437));
    Odrv12 I__469 (
            .O(N__4437),
            .I(CMA_c_5));
    CascadeMux I__468 (
            .O(N__4434),
            .I(\U712_CHIP_RAM.N_387_cascade_ ));
    InMux I__467 (
            .O(N__4431),
            .I(N__4428));
    LocalMux I__466 (
            .O(N__4428),
            .I(N__4424));
    InMux I__465 (
            .O(N__4427),
            .I(N__4421));
    Span4Mux_h I__464 (
            .O(N__4424),
            .I(N__4416));
    LocalMux I__463 (
            .O(N__4421),
            .I(N__4416));
    Span4Mux_v I__462 (
            .O(N__4416),
            .I(N__4413));
    Span4Mux_h I__461 (
            .O(N__4413),
            .I(N__4410));
    Sp12to4 I__460 (
            .O(N__4410),
            .I(N__4407));
    Odrv12 I__459 (
            .O(N__4407),
            .I(AWEn_c));
    InMux I__458 (
            .O(N__4404),
            .I(N__4395));
    InMux I__457 (
            .O(N__4403),
            .I(N__4395));
    InMux I__456 (
            .O(N__4402),
            .I(N__4395));
    LocalMux I__455 (
            .O(N__4395),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__454 (
            .O(N__4392),
            .I(\U712_CHIP_RAM.N_186_cascade_ ));
    InMux I__453 (
            .O(N__4389),
            .I(N__4386));
    LocalMux I__452 (
            .O(N__4386),
            .I(N__4383));
    Odrv4 I__451 (
            .O(N__4383),
            .I(DBR_SYNCZ0Z_0));
    InMux I__450 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__449 (
            .O(N__4377),
            .I(\U712_CHIP_RAM.DBENn_8_0 ));
    InMux I__448 (
            .O(N__4374),
            .I(N__4371));
    LocalMux I__447 (
            .O(N__4371),
            .I(N__4368));
    Odrv4 I__446 (
            .O(N__4368),
            .I(\U712_CHIP_RAM.N_341 ));
    CascadeMux I__445 (
            .O(N__4365),
            .I(\U712_CHIP_RAM.N_341_cascade_ ));
    InMux I__444 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__443 (
            .O(N__4359),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0 ));
    InMux I__442 (
            .O(N__4356),
            .I(N__4352));
    InMux I__441 (
            .O(N__4355),
            .I(N__4349));
    LocalMux I__440 (
            .O(N__4352),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ));
    LocalMux I__439 (
            .O(N__4349),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ));
    CEMux I__438 (
            .O(N__4344),
            .I(N__4341));
    LocalMux I__437 (
            .O(N__4341),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ));
    InMux I__436 (
            .O(N__4338),
            .I(N__4335));
    LocalMux I__435 (
            .O(N__4335),
            .I(N__4332));
    Span4Mux_h I__434 (
            .O(N__4332),
            .I(N__4329));
    Span4Mux_v I__433 (
            .O(N__4329),
            .I(N__4326));
    Sp12to4 I__432 (
            .O(N__4326),
            .I(N__4323));
    Odrv12 I__431 (
            .O(N__4323),
            .I(A_c_20));
    InMux I__430 (
            .O(N__4320),
            .I(N__4316));
    CascadeMux I__429 (
            .O(N__4319),
            .I(N__4313));
    LocalMux I__428 (
            .O(N__4316),
            .I(N__4310));
    InMux I__427 (
            .O(N__4313),
            .I(N__4307));
    Span4Mux_h I__426 (
            .O(N__4310),
            .I(N__4304));
    LocalMux I__425 (
            .O(N__4307),
            .I(N__4301));
    Odrv4 I__424 (
            .O(N__4304),
            .I(DBRn_c_i));
    Odrv4 I__423 (
            .O(N__4301),
            .I(DBRn_c_i));
    IoInMux I__422 (
            .O(N__4296),
            .I(N__4293));
    LocalMux I__421 (
            .O(N__4293),
            .I(N__4290));
    Span12Mux_s11_v I__420 (
            .O(N__4290),
            .I(N__4287));
    Odrv12 I__419 (
            .O(N__4287),
            .I(VBENn_c));
    InMux I__418 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__417 (
            .O(N__4281),
            .I(N__4278));
    Span4Mux_h I__416 (
            .O(N__4278),
            .I(N__4275));
    Sp12to4 I__415 (
            .O(N__4275),
            .I(N__4272));
    Span12Mux_v I__414 (
            .O(N__4272),
            .I(N__4269));
    Odrv12 I__413 (
            .O(N__4269),
            .I(A_c_14));
    InMux I__412 (
            .O(N__4266),
            .I(N__4263));
    LocalMux I__411 (
            .O(N__4263),
            .I(N__4260));
    Span4Mux_h I__410 (
            .O(N__4260),
            .I(N__4257));
    Span4Mux_v I__409 (
            .O(N__4257),
            .I(N__4254));
    Sp12to4 I__408 (
            .O(N__4254),
            .I(N__4251));
    Odrv12 I__407 (
            .O(N__4251),
            .I(A_c_7));
    CascadeMux I__406 (
            .O(N__4248),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ));
    CascadeMux I__405 (
            .O(N__4245),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ));
    IoInMux I__404 (
            .O(N__4242),
            .I(N__4239));
    LocalMux I__403 (
            .O(N__4239),
            .I(N__4236));
    Span4Mux_s3_v I__402 (
            .O(N__4236),
            .I(N__4233));
    Span4Mux_v I__401 (
            .O(N__4233),
            .I(N__4230));
    Sp12to4 I__400 (
            .O(N__4230),
            .I(N__4227));
    Span12Mux_s11_h I__399 (
            .O(N__4227),
            .I(N__4223));
    InMux I__398 (
            .O(N__4226),
            .I(N__4220));
    Odrv12 I__397 (
            .O(N__4223),
            .I(LATCH_CLK_c));
    LocalMux I__396 (
            .O(N__4220),
            .I(LATCH_CLK_c));
    InMux I__395 (
            .O(N__4215),
            .I(N__4212));
    LocalMux I__394 (
            .O(N__4212),
            .I(\U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0 ));
    IoInMux I__393 (
            .O(N__4209),
            .I(N__4206));
    LocalMux I__392 (
            .O(N__4206),
            .I(N__4203));
    Span4Mux_s3_v I__391 (
            .O(N__4203),
            .I(N__4200));
    Span4Mux_v I__390 (
            .O(N__4200),
            .I(N__4197));
    Span4Mux_v I__389 (
            .O(N__4197),
            .I(N__4194));
    Span4Mux_v I__388 (
            .O(N__4194),
            .I(N__4190));
    InMux I__387 (
            .O(N__4193),
            .I(N__4187));
    Odrv4 I__386 (
            .O(N__4190),
            .I(DBDIR_c));
    LocalMux I__385 (
            .O(N__4187),
            .I(DBDIR_c));
    IoInMux I__384 (
            .O(N__4182),
            .I(N__4179));
    LocalMux I__383 (
            .O(N__4179),
            .I(N__4176));
    Odrv12 I__382 (
            .O(N__4176),
            .I(DBRn_c_i_0));
    IoInMux I__381 (
            .O(N__4173),
            .I(N__4170));
    LocalMux I__380 (
            .O(N__4170),
            .I(N__4167));
    Span4Mux_s3_v I__379 (
            .O(N__4167),
            .I(N__4164));
    Span4Mux_h I__378 (
            .O(N__4164),
            .I(N__4161));
    Odrv4 I__377 (
            .O(N__4161),
            .I(CLK80_PLL_i_i));
    IoInMux I__376 (
            .O(N__4158),
            .I(N__4155));
    LocalMux I__375 (
            .O(N__4155),
            .I(N__4152));
    Span4Mux_s2_h I__374 (
            .O(N__4152),
            .I(N__4149));
    Span4Mux_h I__373 (
            .O(N__4149),
            .I(N__4146));
    Span4Mux_v I__372 (
            .O(N__4146),
            .I(N__4143));
    Odrv4 I__371 (
            .O(N__4143),
            .I(N_861_i));
    InMux I__370 (
            .O(N__4140),
            .I(N__4136));
    InMux I__369 (
            .O(N__4139),
            .I(N__4133));
    LocalMux I__368 (
            .O(N__4136),
            .I(N__4128));
    LocalMux I__367 (
            .O(N__4133),
            .I(N__4128));
    Span4Mux_v I__366 (
            .O(N__4128),
            .I(N__4125));
    Span4Mux_h I__365 (
            .O(N__4125),
            .I(N__4122));
    Sp12to4 I__364 (
            .O(N__4122),
            .I(N__4119));
    Span12Mux_v I__363 (
            .O(N__4119),
            .I(N__4116));
    Odrv12 I__362 (
            .O(N__4116),
            .I(DBRn_c));
    IoInMux I__361 (
            .O(N__4113),
            .I(N__4110));
    LocalMux I__360 (
            .O(N__4110),
            .I(N__4107));
    Span4Mux_s0_v I__359 (
            .O(N__4107),
            .I(N__4104));
    Span4Mux_v I__358 (
            .O(N__4104),
            .I(N__4101));
    Sp12to4 I__357 (
            .O(N__4101),
            .I(N__4098));
    Span12Mux_h I__356 (
            .O(N__4098),
            .I(N__4095));
    Span12Mux_v I__355 (
            .O(N__4095),
            .I(N__4092));
    Odrv12 I__354 (
            .O(N__4092),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__5467));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__5469));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__5470));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__5465));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__5466));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__5468));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__5471));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__5472));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4925),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7722),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4182),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__7308),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_2  (
            .in0(N__10017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4320),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10707),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_3_14_5.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_3_14_5.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_3_14_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_3_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4503),
            .lcout(N_861_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_10_1.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4139),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_6_10_5.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_6_10_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_6_10_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_6_10_5 (
            .in0(N__4140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10693),
            .ce(),
            .sr(N__9991));
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_7_10_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_7_10_0  (
            .in0(N__10325),
            .in1(N__9212),
            .in2(N__4319),
            .in3(N__5009),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__9984));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__8821),
            .in2(_gnd_net_),
            .in3(N__9842),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_8_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_8_8_1  (
            .in0(N__4284),
            .in1(N__4266),
            .in2(_gnd_net_),
            .in3(N__9396),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_8_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_8_2  (
            .in0(N__9397),
            .in1(N__8820),
            .in2(N__4248),
            .in3(N__8937),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_9_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_9_1  (
            .in0(N__4547),
            .in1(N__4374),
            .in2(N__6948),
            .in3(N__6270),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_9_2 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_8_9_2  (
            .in0(N__8194),
            .in1(N__4226),
            .in2(N__4245),
            .in3(N__4215),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10679),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_9_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__7179),
            .in2(_gnd_net_),
            .in3(N__5613),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_8_9_6 .LUT_INIT=16'b0000101001001010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_8_9_6  (
            .in0(N__10802),
            .in1(N__10952),
            .in2(N__9402),
            .in3(N__8787),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_10_1  (
            .in0(N__4427),
            .in1(N__4193),
            .in2(_gnd_net_),
            .in3(N__4548),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10684),
            .ce(),
            .sr(N__9978));
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_8_10_2  (
            .in0(N__5559),
            .in1(N__4356),
            .in2(_gnd_net_),
            .in3(N__4380),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10684),
            .ce(),
            .sr(N__9978));
    defparam DBR_SYNC_1_LC_8_10_4.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_8_10_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_8_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4389),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10684),
            .ce(),
            .sr(N__9978));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__10016),
            .in2(_gnd_net_),
            .in3(N__4355),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_8_11_3  (
            .in0(N__6236),
            .in1(N__6166),
            .in2(_gnd_net_),
            .in3(N__8922),
            .lcout(\U712_CHIP_RAM.DBENn_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_11_4  (
            .in0(N__7175),
            .in1(N__7050),
            .in2(N__6360),
            .in3(N__11096),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_8_11_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_8_11_6  (
            .in0(N__4746),
            .in1(N__7051),
            .in2(N__7182),
            .in3(N__6921),
            .lcout(\U712_CHIP_RAM.N_341 ),
            .ltout(\U712_CHIP_RAM.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIBTHEC_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIBTHEC_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIBTHEC_LC_8_11_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIBTHEC_LC_8_11_7  (
            .in0(N__6922),
            .in1(N__4546),
            .in2(N__4365),
            .in3(N__4362),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0  (
            .in0(N__6171),
            .in1(N__6492),
            .in2(N__6252),
            .in3(N__6598),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10694),
            .ce(N__4344),
            .sr(N__9965));
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_12_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_3_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__10326),
            .in2(_gnd_net_),
            .in3(N__4338),
            .lcout(\U712_CHIP_RAM.BANK0_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_0  (
            .in0(N__8195),
            .in1(N__7386),
            .in2(_gnd_net_),
            .in3(N__7416),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10698),
            .ce(N__4731),
            .sr(N__9958));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_14_0 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_14_0  (
            .in0(N__4472),
            .in1(N__8619),
            .in2(N__5241),
            .in3(N__7455),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10701),
            .ce(),
            .sr(N__9950));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_9_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_9_8_2  (
            .in0(N__4800),
            .in1(N__4461),
            .in2(_gnd_net_),
            .in3(N__4455),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10669),
            .ce(N__10565),
            .sr(N__9985));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_9_0  (
            .in0(N__6591),
            .in1(N__4403),
            .in2(N__6789),
            .in3(N__8435),
            .lcout(\U712_CHIP_RAM.N_387 ),
            .ltout(\U712_CHIP_RAM.N_387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_9_9_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__6235),
            .in2(N__4434),
            .in3(N__6162),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_2 .LUT_INIT=16'b0011010100110101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_2  (
            .in0(N__11341),
            .in1(N__4431),
            .in2(N__6599),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_3 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_3  (
            .in0(N__4404),
            .in1(N__4833),
            .in2(N__8213),
            .in3(N__8778),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10674),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_9_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__8434),
            .lcout(\U712_CHIP_RAM.N_186 ),
            .ltout(\U712_CHIP_RAM.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_9_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_9_5  (
            .in0(N__8202),
            .in1(N__6590),
            .in2(N__4392),
            .in3(N__6782),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_9_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_3_LC_9_9_6  (
            .in0(N__8777),
            .in1(N__7174),
            .in2(_gnd_net_),
            .in3(N__7059),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_9_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_9_9_7  (
            .in0(N__11100),
            .in1(N__6674),
            .in2(_gnd_net_),
            .in3(N__6361),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_9_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_9_10_0  (
            .in0(N__6563),
            .in1(N__6491),
            .in2(N__6246),
            .in3(N__6135),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_10_1 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_10_1  (
            .in0(N__7157),
            .in1(N__7019),
            .in2(N__6368),
            .in3(N__11094),
            .lcout(\U712_CHIP_RAM.N_385 ),
            .ltout(\U712_CHIP_RAM.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_10_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_10_2  (
            .in0(N__4530),
            .in1(N__6855),
            .in2(N__4524),
            .in3(N__6937),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_3  (
            .in0(N__8196),
            .in1(N__8788),
            .in2(N__4521),
            .in3(N__5024),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4  (
            .in0(N__11095),
            .in1(N__8197),
            .in2(N__4518),
            .in3(N__4562),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_3_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_3_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_3_LC_9_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_3_LC_9_10_5  (
            .in0(N__7156),
            .in1(N__6343),
            .in2(N__6680),
            .in3(N__7018),
            .lcout(\U712_CHIP_RAM.N_335 ),
            .ltout(\U712_CHIP_RAM.N_335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_10_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__6490),
            .in2(N__4509),
            .in3(N__6134),
            .lcout(\U712_CHIP_RAM.N_342 ),
            .ltout(\U712_CHIP_RAM.N_342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_9_10_7 .LUT_INIT=16'b1100000011010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_9_10_7  (
            .in0(N__4953),
            .in1(N__6564),
            .in2(N__4506),
            .in3(N__6787),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_11_0  (
            .in0(N__5880),
            .in1(N__4632),
            .in2(N__4623),
            .in3(N__6140),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CLK_EN_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_11_1 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_11_1  (
            .in0(N__4598),
            .in1(_gnd_net_),
            .in2(N__4611),
            .in3(N__4587),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10685),
            .ce(),
            .sr(N__9966));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_11_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_11_2  (
            .in0(N__7155),
            .in1(N__4745),
            .in2(N__6943),
            .in3(N__7044),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5O1M2_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5O1M2_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5O1M2_LC_9_11_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5O1M2_LC_9_11_3  (
            .in0(N__6662),
            .in1(N__5879),
            .in2(N__6161),
            .in3(N__6480),
            .lcout(\U712_CHIP_RAM.N_338 ),
            .ltout(\U712_CHIP_RAM.N_338_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_11_4 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_11_4  (
            .in0(N__4581),
            .in1(N__7043),
            .in2(N__4575),
            .in3(N__4744),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_11_5 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4572),
            .in3(N__8161),
            .lcout(\U712_CHIP_RAM.N_239 ),
            .ltout(\U712_CHIP_RAM.N_239_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_3_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_3_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_3_LC_9_11_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_3_LC_9_11_6  (
            .in0(N__5082),
            .in1(N__5659),
            .in2(N__4569),
            .in3(N__5538),
            .lcout(\U712_CHIP_RAM.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_9_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_9_12_1  (
            .in0(N__8188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6332),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_12_2  (
            .in0(N__5165),
            .in1(N__5049),
            .in2(N__4566),
            .in3(N__8187),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10690),
            .ce(N__5717),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_9_12_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__5602),
            .in2(_gnd_net_),
            .in3(N__6331),
            .lcout(\U712_CHIP_RAM.N_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_12_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_12_4  (
            .in0(N__7060),
            .in1(N__8186),
            .in2(_gnd_net_),
            .in3(N__7208),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_12_5  (
            .in0(N__6342),
            .in1(N__5883),
            .in2(_gnd_net_),
            .in3(N__5499),
            .lcout(\U712_CHIP_RAM.N_269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__10015),
            .in2(_gnd_net_),
            .in3(N__5109),
            .lcout(\U712_CYCLE_TERM.N_217_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_13_0 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_13_0  (
            .in0(N__5256),
            .in1(N__7353),
            .in2(N__8352),
            .in3(N__5675),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10695),
            .ce(),
            .sr(N__9951));
    defparam \U712_REG_SM.ASn_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_9_13_4 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \U712_REG_SM.ASn_LC_9_13_4  (
            .in0(N__8302),
            .in1(N__5250),
            .in2(N__8418),
            .in3(N__4699),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10695),
            .ce(),
            .sr(N__9951));
    defparam \U712_REG_SM.START_RST_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_9_13_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_9_13_6  (
            .in0(N__4686),
            .in1(N__5103),
            .in2(_gnd_net_),
            .in3(N__6051),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10695),
            .ce(),
            .sr(N__9951));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_14_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__4685),
            .in2(_gnd_net_),
            .in3(N__5271),
            .lcout(),
            .ltout(\U712_REG_SM.N_270_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_2 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_14_2  (
            .in0(N__8217),
            .in1(N__4670),
            .in2(N__4635),
            .in3(N__4884),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10699),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__8216),
            .in2(_gnd_net_),
            .in3(N__5220),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10699),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4890),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10702),
            .ce(),
            .sr(N__9945));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4926),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10703),
            .ce(),
            .sr(N__9944));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__4883),
            .in2(_gnd_net_),
            .in3(N__4848),
            .lcout(\U712_CHIP_RAM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7  (
            .in0(N__4752),
            .in1(N__4779),
            .in2(_gnd_net_),
            .in3(N__5433),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10666),
            .ce(N__10556),
            .sr(N__9979));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_9_0 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_9_0  (
            .in0(N__8774),
            .in1(N__10956),
            .in2(N__10819),
            .in3(N__9398),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_9_1  (
            .in0(N__4794),
            .in1(N__8773),
            .in2(_gnd_net_),
            .in3(N__8658),
            .lcout(\U712_CHIP_RAM.N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_9_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_9_2  (
            .in0(N__8775),
            .in1(N__4769),
            .in2(N__7957),
            .in3(N__8639),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_9_3 .LUT_INIT=16'b1110010011101100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_9_3  (
            .in0(N__8198),
            .in1(N__6575),
            .in2(N__7869),
            .in3(N__5623),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10670),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_9_5 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_9_5  (
            .in0(N__8640),
            .in1(N__7948),
            .in2(N__4773),
            .in3(N__8776),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_10_10_0 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_10_10_0  (
            .in0(N__5037),
            .in1(N__4959),
            .in2(N__5025),
            .in3(N__5010),
            .lcout(),
            .ltout(\U712_CHIP_RAM.BANK0_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_10_10_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_10_10_1  (
            .in0(N__4970),
            .in1(N__4995),
            .in2(N__4989),
            .in3(N__4938),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10675),
            .ce(),
            .sr(N__9967));
    defparam \U712_CHIP_RAM.BANK0_RNO_4_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_4_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_4_LC_10_10_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_4_LC_10_10_2  (
            .in0(N__6233),
            .in1(N__6152),
            .in2(_gnd_net_),
            .in3(N__6565),
            .lcout(\U712_CHIP_RAM.BANK0_RNOZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_10_10_3 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_10_10_3  (
            .in0(N__4952),
            .in1(N__6234),
            .in2(N__6583),
            .in3(N__6788),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_10_10_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4941),
            .in3(N__5660),
            .lcout(\U712_CHIP_RAM.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_10_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_10_5  (
            .in0(N__5888),
            .in1(N__6479),
            .in2(_gnd_net_),
            .in3(N__6136),
            .lcout(\U712_CHIP_RAM.N_333 ),
            .ltout(\U712_CHIP_RAM.N_333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI27TJ3_3_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI27TJ3_3_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI27TJ3_3_LC_10_10_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI27TJ3_3_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__6697),
            .in2(N__4932),
            .in3(N__6673),
            .lcout(\U712_CHIP_RAM.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_10_11_1  (
            .in0(N__6661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7025),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_10_11_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_10_11_2  (
            .in0(N__6698),
            .in1(N__5881),
            .in2(N__4929),
            .in3(N__6142),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER18 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7UUV6_4_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7UUV6_4_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7UUV6_4_LC_10_11_3 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7UUV6_4_LC_10_11_3  (
            .in0(N__6143),
            .in1(_gnd_net_),
            .in2(N__5085),
            .in3(N__6232),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_4 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_4  (
            .in0(N__5061),
            .in1(N__5076),
            .in2(N__5169),
            .in3(N__5070),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10681),
            .ce(N__5713),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_10_11_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_10_11_5  (
            .in0(N__6660),
            .in1(N__7144),
            .in2(_gnd_net_),
            .in3(N__7024),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_0_0_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_10_11_6 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_10_11_6  (
            .in0(N__6481),
            .in1(N__5534),
            .in2(N__5064),
            .in3(N__6141),
            .lcout(\U712_CHIP_RAM.N_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7  (
            .in0(N__5120),
            .in1(N__5183),
            .in2(_gnd_net_),
            .in3(N__5198),
            .lcout(\U712_CHIP_RAM.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__7045),
            .in2(_gnd_net_),
            .in3(N__5055),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_12_1  (
            .in0(N__5158),
            .in1(N__7154),
            .in2(_gnd_net_),
            .in3(N__5052),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__6355),
            .in2(_gnd_net_),
            .in3(N__5043),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_3  (
            .in0(N__5159),
            .in1(N__6675),
            .in2(_gnd_net_),
            .in3(N__5040),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_12_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_12_4  (
            .in0(N__5156),
            .in1(N__5884),
            .in2(_gnd_net_),
            .in3(N__5202),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_12_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_12_5  (
            .in0(N__5160),
            .in1(N__5199),
            .in2(_gnd_net_),
            .in3(N__5187),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_12_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_12_6  (
            .in0(N__5157),
            .in1(N__5184),
            .in2(_gnd_net_),
            .in3(N__5172),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_12_7  (
            .in0(N__5161),
            .in1(N__5121),
            .in2(_gnd_net_),
            .in3(N__5124),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10686),
            .ce(N__5718),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_10_13_0 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_10_13_0  (
            .in0(N__7466),
            .in1(N__8190),
            .in2(N__7415),
            .in3(N__7385),
            .lcout(\U712_CYCLE_TERM.N_217_i_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.START_RST_RNO_0_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_RNO_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.START_RST_RNO_0_LC_10_13_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.START_RST_RNO_0_LC_10_13_1  (
            .in0(N__5097),
            .in1(N__5273),
            .in2(N__8310),
            .in3(N__8413),
            .lcout(\U712_REG_SM.START_RST_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_13_2 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_13_2  (
            .in0(N__5272),
            .in1(N__5096),
            .in2(N__6054),
            .in3(N__8300),
            .lcout(),
            .ltout(\U712_REG_SM.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_13_3 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_10_13_3  (
            .in0(N__8301),
            .in1(N__8191),
            .in2(N__5088),
            .in3(N__8414),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10691),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_13_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_13_4  (
            .in0(N__5283),
            .in1(N__8189),
            .in2(_gnd_net_),
            .in3(N__6470),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10691),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_13_5  (
            .in0(N__6732),
            .in1(N__5274),
            .in2(_gnd_net_),
            .in3(N__8346),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_REG_SM.ASn_RNO_0_LC_10_13_6  (
            .in0(N__6047),
            .in1(N__6733),
            .in2(_gnd_net_),
            .in3(N__8296),
            .lcout(\U712_REG_SM.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_10_14_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_10_14_0  (
            .in0(N__8613),
            .in1(N__8193),
            .in2(_gnd_net_),
            .in3(N__7451),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_10_14_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_10_14_1  (
            .in0(N__5240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8214),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_14_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_14_2  (
            .in0(N__5484),
            .in1(N__5297),
            .in2(_gnd_net_),
            .in3(N__5312),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_14_3 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_14_3  (
            .in0(N__8192),
            .in1(N__5345),
            .in2(N__5244),
            .in3(N__5208),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__5239),
            .in2(_gnd_net_),
            .in3(N__5219),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_14_5 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_14_5  (
            .in0(N__5360),
            .in1(N__5390),
            .in2(N__5331),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_14_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_14_6  (
            .in0(N__8412),
            .in1(N__8486),
            .in2(_gnd_net_),
            .in3(N__8276),
            .lcout(),
            .ltout(\U712_REG_SM.N_284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_10_14_7  (
            .in0(N__7348),
            .in1(N__5904),
            .in2(N__5394),
            .in3(N__8215),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_15_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_15_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__5391),
            .in2(_gnd_net_),
            .in3(N__5379),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_15_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_15_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__5376),
            .in2(_gnd_net_),
            .in3(N__5364),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_15_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__5361),
            .in2(_gnd_net_),
            .in3(N__5349),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_15_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__5346),
            .in2(_gnd_net_),
            .in3(N__5334),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_15_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_15_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__5330),
            .in2(_gnd_net_),
            .in3(N__5316),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_15_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_15_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__5313),
            .in2(_gnd_net_),
            .in3(N__5301),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_15_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_15_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__5298),
            .in2(_gnd_net_),
            .in3(N__5286),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_15_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__5483),
            .in2(_gnd_net_),
            .in3(N__5487),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5464),
            .ce(),
            .sr(N__7494));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_9_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_9_1  (
            .in0(N__7663),
            .in1(N__9362),
            .in2(_gnd_net_),
            .in3(N__7612),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_0_LC_11_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_0_LC_11_9_3  (
            .in0(N__5579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5627),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_9_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_9_5  (
            .in0(N__9363),
            .in1(N__10803),
            .in2(_gnd_net_),
            .in3(N__5439),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_116_i_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_116_i_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_116_i_LC_11_10_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_116_i_LC_11_10_0  (
            .in0(N__11286),
            .in1(N__5780),
            .in2(N__7737),
            .in3(N__8810),
            .lcout(N_116_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_11_10_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__7158),
            .in2(_gnd_net_),
            .in3(N__6362),
            .lcout(\U712_CHIP_RAM.N_207 ),
            .ltout(\U712_CHIP_RAM.N_207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_10_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5403),
            .in3(N__8809),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_10_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_10_5  (
            .in0(N__11132),
            .in1(N__6679),
            .in2(N__5400),
            .in3(N__7049),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_6 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_6  (
            .in0(N__5523),
            .in1(N__5889),
            .in2(N__5397),
            .in3(N__6160),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10671),
            .ce(N__5634),
            .sr(N__9959));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_11_0  (
            .in0(N__6659),
            .in1(N__7022),
            .in2(N__5661),
            .in3(N__5517),
            .lcout(\U712_CHIP_RAM.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_1  (
            .in0(N__7021),
            .in1(N__7152),
            .in2(N__6369),
            .in3(N__6941),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_2  (
            .in0(N__6942),
            .in1(N__6263),
            .in2(N__5640),
            .in3(N__7204),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_3  (
            .in0(N__10014),
            .in1(_gnd_net_),
            .in2(N__5637),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_11_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_11_4  (
            .in0(N__5628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5578),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_11_5 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_11_5  (
            .in0(N__7023),
            .in1(N__11137),
            .in2(N__6501),
            .in3(N__6159),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_11_11_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_11_11_6  (
            .in0(N__6658),
            .in1(N__7133),
            .in2(_gnd_net_),
            .in3(N__7020),
            .lcout(\U712_CHIP_RAM.N_334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_11_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_11_7  (
            .in0(N__8830),
            .in1(N__11136),
            .in2(_gnd_net_),
            .in3(N__7153),
            .lcout(\U712_CHIP_RAM.N_297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_11_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_11_12_0  (
            .in0(N__5878),
            .in1(N__5513),
            .in2(_gnd_net_),
            .in3(N__5498),
            .lcout(\U712_CHIP_RAM.N_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISAAQ_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISAAQ_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISAAQ_LC_11_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISAAQ_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__5876),
            .in2(_gnd_net_),
            .in3(N__6463),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_12_2 .LUT_INIT=16'b0000001001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_12_2  (
            .in0(N__6359),
            .in1(N__6666),
            .in2(N__7173),
            .in3(N__7039),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_11_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_11_12_3  (
            .in0(N__6145),
            .in1(N__5685),
            .in2(N__5739),
            .in3(N__5877),
            .lcout(\U712_CHIP_RAM.N_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_12_4 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_12_4  (
            .in0(N__6069),
            .in1(N__5736),
            .in2(N__6825),
            .in3(N__7661),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_11_12_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_11_12_5  (
            .in0(N__6144),
            .in1(N__6247),
            .in2(_gnd_net_),
            .in3(N__8115),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_392_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4TF5A_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4TF5A_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4TF5A_LC_11_12_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4TF5A_LC_11_12_6  (
            .in0(N__5727),
            .in1(N__6888),
            .in2(N__5721),
            .in3(N__6869),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_13_0  (
            .in0(N__8347),
            .in1(N__6731),
            .in2(N__5679),
            .in3(N__8127),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10687),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__8478),
            .in2(_gnd_net_),
            .in3(N__6041),
            .lcout(\U712_REG_SM.N_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_11_13_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_11_13_3  (
            .in0(N__8126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6464),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_13_4 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_13_4  (
            .in0(N__8304),
            .in1(N__6730),
            .in2(_gnd_net_),
            .in3(N__8395),
            .lcout(\U712_REG_SM.N_196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_5  (
            .in0(N__8394),
            .in1(N__8303),
            .in2(_gnd_net_),
            .in3(N__8447),
            .lcout(\U712_REG_SM.N_383 ),
            .ltout(\U712_REG_SM.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_6  (
            .in0(N__8479),
            .in1(_gnd_net_),
            .in2(N__5892),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_281 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_13_7 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_13_7  (
            .in0(N__8125),
            .in1(N__5882),
            .in2(_gnd_net_),
            .in3(N__7145),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_14_0 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_14_0  (
            .in0(N__7377),
            .in1(N__7322),
            .in2(N__5823),
            .in3(N__7449),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_14_1 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_11_14_1  (
            .in0(N__8614),
            .in1(N__8128),
            .in2(N__5826),
            .in3(N__7378),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10692),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_11_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__7321),
            .in2(_gnd_net_),
            .in3(N__5819),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_156_i_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_156_i_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_156_i_LC_11_14_4 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_156_i_LC_11_14_4  (
            .in0(N__7259),
            .in1(N__6060),
            .in2(N__5751),
            .in3(N__11209),
            .lcout(N_156_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_126_i_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_126_i_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_126_i_LC_11_14_5 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \U712_BYTE_ENABLE.N_126_i_LC_11_14_5  (
            .in0(N__5784),
            .in1(N__5747),
            .in2(N__11211),
            .in3(N__7743),
            .lcout(N_126_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_11_15_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_11_15_1  (
            .in0(N__8848),
            .in1(N__9563),
            .in2(_gnd_net_),
            .in3(N__9482),
            .lcout(\U712_BYTE_ENABLE.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_11_15_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_11_15_2 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_11_15_2  (
            .in0(N__9712),
            .in1(N__9632),
            .in2(N__9564),
            .in3(N__8847),
            .lcout(\U712_BYTE_ENABLE.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_11_15_5 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_11_15_5  (
            .in0(N__11334),
            .in1(N__6734),
            .in2(_gnd_net_),
            .in3(N__8480),
            .lcout(\U712_REG_SM.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_11_15_6 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_11_15_6  (
            .in0(N__8482),
            .in1(N__6052),
            .in2(N__8306),
            .in3(N__8397),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_11_15_7 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_11_15_7  (
            .in0(N__6053),
            .in1(N__6735),
            .in2(N__8307),
            .in3(N__8481),
            .lcout(\U712_REG_SM.N_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_11_16_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_11_16_5 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \U712_REG_SM.DS_EN_LC_11_16_5  (
            .in0(N__6018),
            .in1(N__6012),
            .in2(N__6006),
            .in3(N__9743),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10700),
            .ce(),
            .sr(N__9942));
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_11_20_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_11_20_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_11_20_0  (
            .in0(N__11148),
            .in1(N__11266),
            .in2(_gnd_net_),
            .in3(N__11205),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_3  (
            .in0(N__9333),
            .in1(N__5964),
            .in2(_gnd_net_),
            .in3(N__5949),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4  (
            .in0(N__5931),
            .in1(N__5916),
            .in2(_gnd_net_),
            .in3(N__9332),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_11_1 .LUT_INIT=16'b1100111111001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_11_1  (
            .in0(N__7058),
            .in1(N__6699),
            .in2(N__6500),
            .in3(N__6681),
            .lcout(\U712_CHIP_RAM.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_11_2 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_11_2  (
            .in0(N__6744),
            .in1(N__6870),
            .in2(N__6600),
            .in3(N__6185),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_11_3 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_11_3  (
            .in0(N__6528),
            .in1(N__6824),
            .in2(N__6522),
            .in3(N__9360),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10668),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_11_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_11_4  (
            .in0(N__6364),
            .in1(N__6519),
            .in2(N__6510),
            .in3(N__6496),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_11_5  (
            .in0(N__6408),
            .in1(N__6387),
            .in2(_gnd_net_),
            .in3(N__9358),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_11_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_11_6  (
            .in0(N__9359),
            .in1(N__8826),
            .in2(N__6372),
            .in3(N__8913),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_1_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_1_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_1_LC_12_11_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_1_LC_12_11_7  (
            .in0(N__7180),
            .in1(N__6363),
            .in2(N__7064),
            .in3(N__11123),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_4_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_4_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_4_LC_12_12_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_4_LC_12_12_0  (
            .in0(N__8071),
            .in1(N__6248),
            .in2(N__6186),
            .in3(N__6170),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_12_12_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__8070),
            .in2(N__6063),
            .in3(N__7212),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_12_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__6823),
            .in2(N__7185),
            .in3(N__9030),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10673),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__7651),
            .in2(_gnd_net_),
            .in3(N__7593),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_12_4 .LUT_INIT=16'b0000001100110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_12_4  (
            .in0(N__7592),
            .in1(N__9029),
            .in2(N__7662),
            .in3(N__9320),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_12_12_5 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_12_12_5  (
            .in0(N__7181),
            .in1(N__8072),
            .in2(N__7065),
            .in3(N__6947),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_12_12_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_12_12_6  (
            .in0(N__6887),
            .in1(N__6868),
            .in2(N__6834),
            .in3(N__6831),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_12_7 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_12_7  (
            .in0(N__6804),
            .in1(N__6798),
            .in2(N__6792),
            .in3(N__7594),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10673),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__8073),
            .in2(_gnd_net_),
            .in3(N__6786),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_12_13_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_12_13_2  (
            .in0(N__6724),
            .in1(N__8396),
            .in2(_gnd_net_),
            .in3(N__8305),
            .lcout(\U712_REG_SM.N_235 ),
            .ltout(\U712_REG_SM.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_13_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__11345),
            .in2(N__7497),
            .in3(N__8341),
            .lcout(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_13_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_13_5  (
            .in0(N__7647),
            .in1(N__7591),
            .in2(N__9037),
            .in3(N__9361),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_12_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_12_13_7 .LUT_INIT=16'b1111100010111000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_12_13_7  (
            .in0(N__7482),
            .in1(N__8074),
            .in2(N__9829),
            .in3(N__7476),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_14_0 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_12_14_0  (
            .in0(N__7470),
            .in1(N__7450),
            .in2(N__7428),
            .in3(N__7408),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10683),
            .ce(),
            .sr(N__9943));
    defparam \U712_REG_SM.REG_TACK_LC_12_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_12_14_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_12_14_2  (
            .in0(N__7352),
            .in1(N__7332),
            .in2(N__7326),
            .in3(N__8223),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10683),
            .ce(),
            .sr(N__9943));
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7269),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10683),
            .ce(),
            .sr(N__9943));
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_12_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7292),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10683),
            .ce(),
            .sr(N__9943));
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_12_15_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_12_15_5 .LUT_INIT=16'b1100111000111011;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_i_o2_LC_12_15_5  (
            .in0(N__9713),
            .in1(N__9558),
            .in2(N__9650),
            .in3(N__9483),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_151_i_LC_12_15_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_151_i_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_151_i_LC_12_15_6 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_151_i_LC_12_15_6  (
            .in0(N__7263),
            .in1(N__11279),
            .in2(N__7242),
            .in3(N__8849),
            .lcout(N_151_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_15_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_12_15_7  (
            .in0(N__9641),
            .in1(N__9714),
            .in2(N__8853),
            .in3(N__9559),
            .lcout(\U712_BYTE_ENABLE.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_16_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_16_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_16_3  (
            .in0(N__9593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9702),
            .lcout(\U712_BYTE_ENABLE.UUBE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8095),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_13_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7613),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10658),
            .ce(),
            .sr(N__9986));
    defparam \U712_CHIP_RAM.RASn_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_6_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7677),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10658),
            .ce(),
            .sr(N__9986));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_7_5  (
            .in0(N__7676),
            .in1(N__9392),
            .in2(N__9051),
            .in3(N__7614),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10660),
            .ce(N__10560),
            .sr(N__9980));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_7_7 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_7_7  (
            .in0(N__7964),
            .in1(N__7503),
            .in2(N__8836),
            .in3(N__7545),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10660),
            .ce(N__10560),
            .sr(N__9980));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_0  (
            .in0(N__9213),
            .in1(N__10315),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10098),
            .ce(N__10059),
            .sr(N__9971));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_9_0  (
            .in0(N__7905),
            .in1(N__7887),
            .in2(_gnd_net_),
            .in3(N__9370),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__7857),
            .in2(_gnd_net_),
            .in3(N__8000),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_7  (
            .in0(N__8131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8001),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10667),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_10_0  (
            .in0(N__7851),
            .in1(N__7833),
            .in2(_gnd_net_),
            .in3(N__9342),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_10_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_10_5  (
            .in0(N__8794),
            .in1(N__7812),
            .in2(N__9380),
            .in3(N__8670),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__8792),
            .in2(_gnd_net_),
            .in3(N__9343),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_7  (
            .in0(N__8793),
            .in1(N__7806),
            .in2(N__9379),
            .in3(N__8646),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_11_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_13_11_6  (
            .in0(N__10850),
            .in1(N__8865),
            .in2(N__10798),
            .in3(N__7800),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10676),
            .ce(N__10543),
            .sr(N__9952));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_12_3  (
            .in0(N__7779),
            .in1(N__7761),
            .in2(_gnd_net_),
            .in3(N__9356),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_12_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_12_4  (
            .in0(N__9357),
            .in1(N__8825),
            .in2(N__8499),
            .in3(N__8625),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_12_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__10013),
            .in2(_gnd_net_),
            .in3(N__8496),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_13_0 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_13_0  (
            .in0(N__8490),
            .in1(N__8399),
            .in2(N__8351),
            .in3(N__8451),
            .lcout(),
            .ltout(\U712_REG_SM.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_13_1 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_13_13_1  (
            .in0(N__8400),
            .in1(N__8130),
            .in2(N__8421),
            .in3(N__8309),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10688),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_13_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_13_13_5 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_13_13_5  (
            .in0(N__8398),
            .in1(N__8342),
            .in2(_gnd_net_),
            .in3(N__8308),
            .lcout(\U712_REG_SM.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_7 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_13_13_7  (
            .in0(N__11210),
            .in1(N__8129),
            .in2(_gnd_net_),
            .in3(N__11272),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10688),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_7_7 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_7_7  (
            .in0(N__7989),
            .in1(N__8824),
            .in2(N__7968),
            .in3(N__9156),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10661),
            .ce(N__10555),
            .sr(N__9987));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_8_5  (
            .in0(N__10254),
            .in1(N__9208),
            .in2(_gnd_net_),
            .in3(N__9140),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10063),
            .sr(N__9981));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_4  (
            .in0(N__8822),
            .in1(N__8664),
            .in2(N__7914),
            .in3(N__9400),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_9_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_9_7  (
            .in0(N__9399),
            .in1(N__8823),
            .in2(N__8685),
            .in3(N__8676),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_10_0  (
            .in0(N__9139),
            .in1(N__10253),
            .in2(_gnd_net_),
            .in3(N__10418),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10056),
            .sr(N__9968));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_10_1  (
            .in0(N__10252),
            .in1(N__10464),
            .in2(_gnd_net_),
            .in3(N__10929),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10056),
            .sr(N__9968));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_11_2  (
            .in0(N__10372),
            .in1(N__10251),
            .in2(_gnd_net_),
            .in3(N__8901),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10054),
            .sr(N__9960));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_7  (
            .in0(N__8900),
            .in1(N__10250),
            .in2(_gnd_net_),
            .in3(N__11027),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10054),
            .sr(N__9960));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_6  (
            .in0(N__11028),
            .in1(N__10310),
            .in2(_gnd_net_),
            .in3(N__8899),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10096),
            .ce(N__10057),
            .sr(N__9953));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_13_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_13_3  (
            .in0(N__10149),
            .in1(N__10309),
            .in2(_gnd_net_),
            .in3(N__10923),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10060),
            .sr(N__9946));
    defparam pll_RNI8MQ3_LC_14_14_1.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_14_14_1.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_14_14_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8618),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_0 .LUT_INIT=16'b0000110111000000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_LC_14_20_0  (
            .in0(N__9648),
            .in1(N__9698),
            .in2(N__9528),
            .in3(N__9465),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_14_20_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_LC_14_20_4  (
            .in0(N__9649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9699),
            .lcout(U712_BYTE_ENABLE_UUBE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_15_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9050),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10659),
            .ce(),
            .sr(N__9993));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_8_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_15_8_6  (
            .in0(N__10877),
            .in1(N__9102),
            .in2(N__10827),
            .in3(N__8985),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10672),
            .ce(N__10566),
            .sr(N__9988));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_15_9_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_15_9_0  (
            .in0(N__10887),
            .in1(N__10876),
            .in2(N__10826),
            .in3(N__8958),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10677),
            .ce(N__10561),
            .sr(N__9982));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_7  (
            .in0(N__10311),
            .in1(N__10417),
            .in2(_gnd_net_),
            .in3(N__10463),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10061),
            .sr(N__9972));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_4  (
            .in0(N__10986),
            .in1(N__10300),
            .in2(_gnd_net_),
            .in3(N__11023),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10055),
            .sr(N__9969));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_12_5  (
            .in0(N__10148),
            .in1(N__10308),
            .in2(_gnd_net_),
            .in3(N__10374),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10062),
            .sr(N__9961));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_13_4  (
            .in0(N__10307),
            .in1(N__10373),
            .in2(_gnd_net_),
            .in3(N__8890),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10097),
            .ce(N__10064),
            .sr(N__9954));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_15_19_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_LC_15_19_3 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_LC_15_19_3  (
            .in0(N__9642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9755),
            .lcout(U712_BYTE_ENABLE_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_15_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_15_20_0 .LUT_INIT=16'b0001000100101010;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_LC_15_20_0  (
            .in0(N__9479),
            .in1(N__9700),
            .in2(N__9651),
            .in3(N__9542),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_15_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_15_20_2 .LUT_INIT=16'b0000111100101111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_15_20_2  (
            .in0(N__9481),
            .in1(N__9647),
            .in2(N__9759),
            .in3(N__9546),
            .lcout(N_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_220_i_LC_15_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_220_i_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_220_i_LC_15_20_3 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_220_i_LC_15_20_3  (
            .in0(N__9701),
            .in1(N__9646),
            .in2(N__9557),
            .in3(N__9480),
            .lcout(N_220_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_16_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9401),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10662),
            .ce(),
            .sr(N__9994));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_1  (
            .in0(N__9225),
            .in1(N__10299),
            .in2(_gnd_net_),
            .in3(N__9207),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10095),
            .ce(N__10068),
            .sr(N__9992));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_9_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_9_1  (
            .in0(N__9129),
            .in1(N__10298),
            .in2(_gnd_net_),
            .in3(N__10419),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10092),
            .ce(N__10065),
            .sr(N__9989));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_16_10_1  (
            .in0(N__10866),
            .in1(N__10380),
            .in2(N__10821),
            .in3(N__9096),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10689),
            .ce(N__10554),
            .sr(N__9983));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_16_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_16_10_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_16_10_3  (
            .in0(N__10865),
            .in1(N__10962),
            .in2(N__10820),
            .in3(N__9072),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10689),
            .ce(N__10554),
            .sr(N__9983));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_11_3  (
            .in0(N__10287),
            .in1(N__11022),
            .in2(_gnd_net_),
            .in3(N__10982),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10093),
            .ce(N__10058),
            .sr(N__9973));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_16_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_16_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_16_11_4  (
            .in0(N__10925),
            .in1(N__10455),
            .in2(_gnd_net_),
            .in3(N__10288),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10093),
            .ce(N__10058),
            .sr(N__9973));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7  (
            .in0(N__10146),
            .in1(N__10289),
            .in2(_gnd_net_),
            .in3(N__10924),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10093),
            .ce(N__10058),
            .sr(N__9973));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_16_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_16_12_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_16_12_1  (
            .in0(N__10878),
            .in1(N__10104),
            .in2(N__10825),
            .in3(N__10737),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10697),
            .ce(N__10547),
            .sr(N__9970));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_3  (
            .in0(N__10456),
            .in1(N__10297),
            .in2(_gnd_net_),
            .in3(N__10413),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10091),
            .ce(N__10066),
            .sr(N__9990));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_12_4  (
            .in0(N__10362),
            .in1(N__10296),
            .in2(_gnd_net_),
            .in3(N__10147),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10094),
            .ce(N__10067),
            .sr(N__9974));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_5  (
            .in0(N__11180),
            .in1(N__9843),
            .in2(_gnd_net_),
            .in3(N__11248),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_7 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_7  (
            .in0(N__11349),
            .in1(N__11247),
            .in2(N__11190),
            .in3(N__11147),
            .lcout(N_238),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

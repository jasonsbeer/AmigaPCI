// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 28 2025 22:04:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    SIZ,
    DRA,
    A,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [1:0] SIZ;
    input [9:0] DRA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11817;
    wire N__11816;
    wire N__11815;
    wire N__11808;
    wire N__11807;
    wire N__11806;
    wire N__11799;
    wire N__11798;
    wire N__11797;
    wire N__11790;
    wire N__11789;
    wire N__11788;
    wire N__11781;
    wire N__11780;
    wire N__11779;
    wire N__11772;
    wire N__11771;
    wire N__11770;
    wire N__11763;
    wire N__11762;
    wire N__11761;
    wire N__11754;
    wire N__11753;
    wire N__11752;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11691;
    wire N__11690;
    wire N__11689;
    wire N__11682;
    wire N__11681;
    wire N__11680;
    wire N__11673;
    wire N__11672;
    wire N__11671;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11637;
    wire N__11636;
    wire N__11635;
    wire N__11628;
    wire N__11627;
    wire N__11626;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11556;
    wire N__11555;
    wire N__11554;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11529;
    wire N__11528;
    wire N__11527;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11502;
    wire N__11501;
    wire N__11500;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11484;
    wire N__11483;
    wire N__11482;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11448;
    wire N__11447;
    wire N__11446;
    wire N__11439;
    wire N__11438;
    wire N__11437;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11421;
    wire N__11420;
    wire N__11419;
    wire N__11412;
    wire N__11411;
    wire N__11410;
    wire N__11403;
    wire N__11402;
    wire N__11401;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11385;
    wire N__11384;
    wire N__11383;
    wire N__11376;
    wire N__11375;
    wire N__11374;
    wire N__11367;
    wire N__11366;
    wire N__11365;
    wire N__11358;
    wire N__11357;
    wire N__11356;
    wire N__11349;
    wire N__11348;
    wire N__11347;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11331;
    wire N__11330;
    wire N__11329;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11313;
    wire N__11312;
    wire N__11311;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11295;
    wire N__11294;
    wire N__11293;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11241;
    wire N__11240;
    wire N__11239;
    wire N__11232;
    wire N__11231;
    wire N__11230;
    wire N__11223;
    wire N__11222;
    wire N__11221;
    wire N__11214;
    wire N__11213;
    wire N__11212;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11196;
    wire N__11195;
    wire N__11194;
    wire N__11187;
    wire N__11186;
    wire N__11185;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11169;
    wire N__11168;
    wire N__11167;
    wire N__11160;
    wire N__11159;
    wire N__11158;
    wire N__11151;
    wire N__11150;
    wire N__11149;
    wire N__11142;
    wire N__11141;
    wire N__11140;
    wire N__11133;
    wire N__11132;
    wire N__11131;
    wire N__11124;
    wire N__11123;
    wire N__11122;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11106;
    wire N__11105;
    wire N__11104;
    wire N__11097;
    wire N__11096;
    wire N__11095;
    wire N__11088;
    wire N__11087;
    wire N__11086;
    wire N__11079;
    wire N__11078;
    wire N__11077;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11061;
    wire N__11060;
    wire N__11059;
    wire N__11052;
    wire N__11051;
    wire N__11050;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10972;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10962;
    wire N__10959;
    wire N__10958;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10954;
    wire N__10953;
    wire N__10952;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10946;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10936;
    wire N__10935;
    wire N__10934;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10843;
    wire N__10840;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10780;
    wire N__10777;
    wire N__10776;
    wire N__10773;
    wire N__10772;
    wire N__10769;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10745;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10715;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10659;
    wire N__10654;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10633;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10583;
    wire N__10580;
    wire N__10575;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10544;
    wire N__10541;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10510;
    wire N__10507;
    wire N__10502;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10461;
    wire N__10460;
    wire N__10459;
    wire N__10454;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10448;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10363;
    wire N__10362;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10300;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10285;
    wire N__10282;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10193;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10178;
    wire N__10177;
    wire N__10176;
    wire N__10175;
    wire N__10174;
    wire N__10171;
    wire N__10170;
    wire N__10165;
    wire N__10162;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10125;
    wire N__10122;
    wire N__10117;
    wire N__10114;
    wire N__10109;
    wire N__10106;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10087;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10057;
    wire N__10056;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10036;
    wire N__10033;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10015;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10004;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9941;
    wire N__9936;
    wire N__9933;
    wire N__9926;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9911;
    wire N__9908;
    wire N__9907;
    wire N__9906;
    wire N__9905;
    wire N__9904;
    wire N__9903;
    wire N__9900;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9863;
    wire N__9862;
    wire N__9857;
    wire N__9852;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9830;
    wire N__9827;
    wire N__9822;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9784;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9769;
    wire N__9766;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9747;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9712;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9707;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9679;
    wire N__9678;
    wire N__9677;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9616;
    wire N__9615;
    wire N__9614;
    wire N__9611;
    wire N__9606;
    wire N__9603;
    wire N__9598;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9461;
    wire N__9460;
    wire N__9457;
    wire N__9456;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9449;
    wire N__9448;
    wire N__9447;
    wire N__9444;
    wire N__9443;
    wire N__9442;
    wire N__9441;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9413;
    wire N__9410;
    wire N__9405;
    wire N__9400;
    wire N__9397;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9385;
    wire N__9380;
    wire N__9375;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9355;
    wire N__9350;
    wire N__9345;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9334;
    wire N__9325;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9115;
    wire N__9114;
    wire N__9113;
    wire N__9112;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9104;
    wire N__9103;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9084;
    wire N__9079;
    wire N__9078;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9070;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9062;
    wire N__9061;
    wire N__9060;
    wire N__9059;
    wire N__9058;
    wire N__9055;
    wire N__9054;
    wire N__9053;
    wire N__9050;
    wire N__9045;
    wire N__9038;
    wire N__9035;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9020;
    wire N__9015;
    wire N__9010;
    wire N__9009;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8972;
    wire N__8967;
    wire N__8960;
    wire N__8957;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8897;
    wire N__8896;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8884;
    wire N__8879;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8864;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8688;
    wire N__8687;
    wire N__8686;
    wire N__8685;
    wire N__8684;
    wire N__8683;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8670;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8662;
    wire N__8661;
    wire N__8660;
    wire N__8659;
    wire N__8658;
    wire N__8657;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8522;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8501;
    wire N__8498;
    wire N__8497;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8482;
    wire N__8481;
    wire N__8480;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8247;
    wire N__8244;
    wire N__8235;
    wire N__8232;
    wire N__8225;
    wire N__8224;
    wire N__8223;
    wire N__8220;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8205;
    wire N__8204;
    wire N__8201;
    wire N__8200;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8181;
    wire N__8174;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8166;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8146;
    wire N__8143;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8032;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7810;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7693;
    wire N__7692;
    wire N__7691;
    wire N__7690;
    wire N__7689;
    wire N__7688;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7628;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7616;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7583;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7571;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7556;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7534;
    wire N__7533;
    wire N__7532;
    wire N__7531;
    wire N__7530;
    wire N__7529;
    wire N__7528;
    wire N__7527;
    wire N__7526;
    wire N__7523;
    wire N__7522;
    wire N__7521;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7517;
    wire N__7516;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7499;
    wire N__7496;
    wire N__7495;
    wire N__7492;
    wire N__7485;
    wire N__7482;
    wire N__7481;
    wire N__7478;
    wire N__7477;
    wire N__7476;
    wire N__7471;
    wire N__7468;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7450;
    wire N__7447;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7437;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7421;
    wire N__7416;
    wire N__7409;
    wire N__7404;
    wire N__7393;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7165;
    wire N__7164;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7156;
    wire N__7155;
    wire N__7148;
    wire N__7141;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7074;
    wire N__7069;
    wire N__7066;
    wire N__7061;
    wire N__7060;
    wire N__7055;
    wire N__7052;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7041;
    wire N__7040;
    wire N__7039;
    wire N__7038;
    wire N__7037;
    wire N__7036;
    wire N__7031;
    wire N__7022;
    wire N__7013;
    wire N__7010;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6998;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6980;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6973;
    wire N__6968;
    wire N__6963;
    wire N__6956;
    wire N__6953;
    wire N__6952;
    wire N__6951;
    wire N__6950;
    wire N__6945;
    wire N__6940;
    wire N__6935;
    wire N__6934;
    wire N__6931;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6896;
    wire N__6893;
    wire N__6892;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6884;
    wire N__6883;
    wire N__6882;
    wire N__6879;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6857;
    wire N__6852;
    wire N__6849;
    wire N__6848;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6829;
    wire N__6826;
    wire N__6821;
    wire N__6816;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6762;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6724;
    wire N__6723;
    wire N__6722;
    wire N__6721;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6699;
    wire N__6696;
    wire N__6691;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6673;
    wire N__6666;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6618;
    wire N__6615;
    wire N__6610;
    wire N__6609;
    wire N__6608;
    wire N__6605;
    wire N__6604;
    wire N__6603;
    wire N__6602;
    wire N__6601;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6585;
    wire N__6584;
    wire N__6581;
    wire N__6576;
    wire N__6571;
    wire N__6568;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6548;
    wire N__6545;
    wire N__6544;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6517;
    wire N__6508;
    wire N__6505;
    wire N__6500;
    wire N__6493;
    wire N__6470;
    wire N__6469;
    wire N__6468;
    wire N__6467;
    wire N__6466;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6443;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6403;
    wire N__6400;
    wire N__6393;
    wire N__6390;
    wire N__6371;
    wire N__6368;
    wire N__6367;
    wire N__6366;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6349;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6323;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6311;
    wire N__6310;
    wire N__6305;
    wire N__6300;
    wire N__6295;
    wire N__6294;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6276;
    wire N__6271;
    wire N__6264;
    wire N__6259;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6182;
    wire N__6179;
    wire N__6178;
    wire N__6175;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6129;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6115;
    wire N__6112;
    wire N__6107;
    wire N__6102;
    wire N__6095;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6079;
    wire N__6078;
    wire N__6073;
    wire N__6070;
    wire N__6069;
    wire N__6068;
    wire N__6063;
    wire N__6060;
    wire N__6055;
    wire N__6050;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5939;
    wire N__5938;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5930;
    wire N__5927;
    wire N__5922;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5904;
    wire N__5903;
    wire N__5902;
    wire N__5897;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5860;
    wire N__5843;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5835;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5818;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5796;
    wire N__5793;
    wire N__5788;
    wire N__5777;
    wire N__5774;
    wire N__5767;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5564;
    wire N__5561;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5497;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5456;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5448;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5435;
    wire N__5432;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5402;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5333;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5284;
    wire N__5283;
    wire N__5282;
    wire N__5279;
    wire N__5274;
    wire N__5271;
    wire N__5264;
    wire N__5263;
    wire N__5262;
    wire N__5261;
    wire N__5260;
    wire N__5257;
    wire N__5252;
    wire N__5247;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5212;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5149;
    wire N__5146;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5108;
    wire N__5107;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5081;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5073;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5016;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__4994;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4949;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4937;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4922;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4892;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4884;
    wire N__4883;
    wire N__4882;
    wire N__4879;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4850;
    wire N__4849;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4688;
    wire N__4685;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4616;
    wire N__4613;
    wire N__4612;
    wire N__4607;
    wire N__4604;
    wire N__4603;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4577;
    wire N__4574;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4485;
    wire N__4484;
    wire N__4483;
    wire N__4482;
    wire N__4481;
    wire N__4474;
    wire N__4471;
    wire N__4464;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4397;
    wire N__4396;
    wire N__4393;
    wire N__4392;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4333;
    wire N__4332;
    wire N__4329;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4315;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4097;
    wire N__4094;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4082;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire N_996_i;
    wire CLK80_PLL_i_i;
    wire \U712_CHIP_RAM.N_186_cascade_ ;
    wire DBDIR_c;
    wire TACK_OUTn;
    wire CLK40_PLL_i_i;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_265_cascade_ ;
    wire \U712_CHIP_RAM.N_265 ;
    wire \U712_CHIP_RAM.N_236_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire \U712_CHIP_RAM.N_426_cascade_ ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0 ;
    wire \U712_CHIP_RAM.N_350_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ;
    wire \U712_CHIP_RAM.N_350 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_287 ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire TACK_EN_i_ess;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_300_cascade_ ;
    wire \U712_CHIP_RAM.N_301 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1 ;
    wire bfn_8_6_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_236 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1 ;
    wire \U712_CHIP_RAM.N_348 ;
    wire \U712_CHIP_RAM.N_437 ;
    wire \U712_CHIP_RAM.N_426 ;
    wire \U712_CHIP_RAM.N_76_cascade_ ;
    wire \U712_CHIP_RAM.N_328 ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.N_438_cascade_ ;
    wire \U712_CHIP_RAM.N_336 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_438 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_247 ;
    wire \U712_CHIP_RAM.N_247_cascade_ ;
    wire \U712_CHIP_RAM.N_244 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0 ;
    wire C3_c;
    wire DBRn_c;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_269_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_269_i_0_en_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire N_249_i;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_ ;
    wire \U712_CHIP_RAM.N_325_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ;
    wire \U712_CHIP_RAM.N_325 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.N_241_cascade_ ;
    wire \U712_CHIP_RAM.N_388_cascade_ ;
    wire \U712_CHIP_RAM.N_325_1 ;
    wire \U712_CHIP_RAM.N_381 ;
    wire \U712_CHIP_RAM.N_386 ;
    wire \U712_CHIP_RAM.N_434_cascade_ ;
    wire \U712_CHIP_RAM.N_439 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_335 ;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_351_cascade_ ;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire DBR_SYNCZ0Z_0;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.m17_i_0_o2_1_cascade_ ;
    wire A_c_7;
    wire \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.m15_i_0_a2_0_0_cascade_ ;
    wire \U712_REG_SM.N_289 ;
    wire \U712_REG_SM.N_358_cascade_ ;
    wire \U712_REG_SM.N_360 ;
    wire \U712_REG_SM.N_359 ;
    wire \U712_REG_SM.N_270_i ;
    wire \U712_REG_SM.REG_TACK_7 ;
    wire REG_TACK;
    wire C1_c;
    wire \U712_REG_SM.N_340_cascade_ ;
    wire REGSPACEn_c;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.N_345 ;
    wire \U712_BYTE_ENABLE.N_374_cascade_ ;
    wire N_51_i;
    wire CONSTANT_ONE_NET;
    wire A_c_10;
    wire A_c_3;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_322_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_CHIP_RAM.N_388 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_271_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1 ;
    wire \U712_CHIP_RAM.N_317 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_434 ;
    wire \U712_CHIP_RAM.N_13 ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_300 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_241 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_360_1_cascade_ ;
    wire \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1 ;
    wire \U712_REG_SM.m17_i_0_o2_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.m17_i_0_o2_1 ;
    wire \U712_REG_SM.N_435 ;
    wire \U712_REG_SM.N_435_cascade_ ;
    wire \U712_REG_SM.N_363 ;
    wire ASn_c;
    wire \U712_REG_SM.ASn_0_sqmuxa ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.m17_i_0_o2 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire RnW_c;
    wire WRITE_CYCLEm;
    wire N_276;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire A_c_16;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_5_0_a2_0 ;
    wire \U712_CHIP_RAM.N_112 ;
    wire CLK_EN_c;
    wire bfn_11_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.N_392 ;
    wire A_c_13;
    wire A_c_6;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_BYTE_ENABLE.N_370 ;
    wire \U712_BYTE_ENABLE.N_369_cascade_ ;
    wire N_55_i;
    wire WEn_c;
    wire CRCSn_c;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0 ;
    wire N_53_i;
    wire \U712_BYTE_ENABLE.N_303 ;
    wire UMBE_0_o2_i;
    wire U712_BYTE_ENABLE_UUBE_i;
    wire CASn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_5;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0 ;
    wire CPU_CYCLEm;
    wire N_57_i;
    wire \U712_BYTE_ENABLE.UUBE ;
    wire N_185;
    wire N_44;
    wire A_c_1;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire N_303_i;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DS_ENm;
    wire A_c_0;
    wire N_337_i;
    wire DRA_c_6;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire AGNUS_REV_c;
    wire RAS0n_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire CASUn_c;
    wire CASLn_c;
    wire DRDENn_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3986),
            .RESETB(N__5729),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11817),
            .DIN(N__11816),
            .DOUT(N__11815),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11817),
            .PADOUT(N__11816),
            .PADIN(N__11815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5501),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11808),
            .DIN(N__11807),
            .DOUT(N__11806),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11808),
            .PADOUT(N__11807),
            .PADIN(N__11806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11799),
            .DIN(N__11798),
            .DOUT(N__11797),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11799),
            .PADOUT(N__11798),
            .PADIN(N__11797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9209),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11790),
            .DIN(N__11789),
            .DOUT(N__11788),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11790),
            .PADOUT(N__11789),
            .PADIN(N__11788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11781),
            .DIN(N__11780),
            .DOUT(N__11779),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11781),
            .PADOUT(N__11780),
            .PADIN(N__11779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11772),
            .DIN(N__11771),
            .DOUT(N__11770),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11772),
            .PADOUT(N__11771),
            .PADIN(N__11770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11763),
            .DIN(N__11762),
            .DOUT(N__11761),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11763),
            .PADOUT(N__11762),
            .PADIN(N__11761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11754),
            .DIN(N__11753),
            .DOUT(N__11752),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11754),
            .PADOUT(N__11753),
            .PADIN(N__11752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11745),
            .DIN(N__11744),
            .DOUT(N__11743),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11745),
            .PADOUT(N__11744),
            .PADIN(N__11743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11736),
            .DIN(N__11735),
            .DOUT(N__11734),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11736),
            .PADOUT(N__11735),
            .PADIN(N__11734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11727),
            .DIN(N__11726),
            .DOUT(N__11725),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11727),
            .PADOUT(N__11726),
            .PADIN(N__11725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8915),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11718),
            .DIN(N__11717),
            .DOUT(N__11716),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11718),
            .PADOUT(N__11717),
            .PADIN(N__11716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8285),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11709),
            .DIN(N__11708),
            .DOUT(N__11707),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11709),
            .PADOUT(N__11708),
            .PADIN(N__11707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11700),
            .DIN(N__11699),
            .DOUT(N__11698),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11700),
            .PADOUT(N__11699),
            .PADIN(N__11698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11691),
            .DIN(N__11690),
            .DOUT(N__11689),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11691),
            .PADOUT(N__11690),
            .PADIN(N__11689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11682),
            .DIN(N__11681),
            .DOUT(N__11680),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11682),
            .PADOUT(N__11681),
            .PADIN(N__11680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4295),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11673),
            .DIN(N__11672),
            .DOUT(N__11671),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11673),
            .PADOUT(N__11672),
            .PADIN(N__11671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11664),
            .DIN(N__11663),
            .DOUT(N__11662),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11664),
            .PADOUT(N__11663),
            .PADIN(N__11662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11655),
            .DIN(N__11654),
            .DOUT(N__11653),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11655),
            .PADOUT(N__11654),
            .PADIN(N__11653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11646),
            .DIN(N__11645),
            .DOUT(N__11644),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11646),
            .PADOUT(N__11645),
            .PADIN(N__11644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11637),
            .DIN(N__11636),
            .DOUT(N__11635),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11637),
            .PADOUT(N__11636),
            .PADIN(N__11635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7901),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11628),
            .DIN(N__11627),
            .DOUT(N__11626),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11628),
            .PADOUT(N__11627),
            .PADIN(N__11626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11619),
            .DIN(N__11618),
            .DOUT(N__11617),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11619),
            .PADOUT(N__11618),
            .PADIN(N__11617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9242),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11610),
            .DIN(N__11609),
            .DOUT(N__11608),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11610),
            .PADOUT(N__11609),
            .PADIN(N__11608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11601),
            .DIN(N__11600),
            .DOUT(N__11599),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11601),
            .PADOUT(N__11600),
            .PADIN(N__11599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11592),
            .DIN(N__11591),
            .DOUT(N__11590),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11592),
            .PADOUT(N__11591),
            .PADIN(N__11590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11583),
            .DIN(N__11582),
            .DOUT(N__11581),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11583),
            .PADOUT(N__11582),
            .PADIN(N__11581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11574),
            .DIN(N__11573),
            .DOUT(N__11572),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11574),
            .PADOUT(N__11573),
            .PADIN(N__11572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11565),
            .DIN(N__11564),
            .DOUT(N__11563),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11565),
            .PADOUT(N__11564),
            .PADIN(N__11563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11556),
            .DIN(N__11555),
            .DOUT(N__11554),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11556),
            .PADOUT(N__11555),
            .PADIN(N__11554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11547),
            .DIN(N__11546),
            .DOUT(N__11545),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11547),
            .PADOUT(N__11546),
            .PADIN(N__11545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11538),
            .DIN(N__11537),
            .DOUT(N__11536),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11538),
            .PADOUT(N__11537),
            .PADIN(N__11536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11529),
            .DIN(N__11528),
            .DOUT(N__11527),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11529),
            .PADOUT(N__11528),
            .PADIN(N__11527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11520),
            .DIN(N__11519),
            .DOUT(N__11518),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11520),
            .PADOUT(N__11519),
            .PADIN(N__11518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11511),
            .DIN(N__11510),
            .DOUT(N__11509),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11511),
            .PADOUT(N__11510),
            .PADIN(N__11509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7883),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11502),
            .DIN(N__11501),
            .DOUT(N__11500),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11502),
            .PADOUT(N__11501),
            .PADIN(N__11500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11493),
            .DIN(N__11492),
            .DOUT(N__11491),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11493),
            .PADOUT(N__11492),
            .PADIN(N__11491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4172),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11484),
            .DIN(N__11483),
            .DOUT(N__11482),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11484),
            .PADOUT(N__11483),
            .PADIN(N__11482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11475),
            .DIN(N__11474),
            .DOUT(N__11473),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11475),
            .PADOUT(N__11474),
            .PADIN(N__11473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4004),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11466),
            .DIN(N__11465),
            .DOUT(N__11464),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11466),
            .PADOUT(N__11465),
            .PADIN(N__11464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11457),
            .DIN(N__11456),
            .DOUT(N__11455),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11457),
            .PADOUT(N__11456),
            .PADIN(N__11455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7112),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11448),
            .DIN(N__11447),
            .DOUT(N__11446),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11448),
            .PADOUT(N__11447),
            .PADIN(N__11446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8081),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuft_iopad (
            .OE(N__11439),
            .DIN(N__11438),
            .DOUT(N__11437),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO RAMENn_obuft_preio (
            .PADOEN(N__11439),
            .PADOUT(N__11438),
            .PADIN(N__11437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11430),
            .DIN(N__11429),
            .DOUT(N__11428),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11430),
            .PADOUT(N__11429),
            .PADIN(N__11428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11421),
            .DIN(N__11420),
            .DOUT(N__11419),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11421),
            .PADOUT(N__11420),
            .PADIN(N__11419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11412),
            .DIN(N__11411),
            .DOUT(N__11410),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11412),
            .PADOUT(N__11411),
            .PADIN(N__11410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11403),
            .DIN(N__11402),
            .DOUT(N__11401),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11403),
            .PADOUT(N__11402),
            .PADIN(N__11401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11394),
            .DIN(N__11393),
            .DOUT(N__11392),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11394),
            .PADOUT(N__11393),
            .PADIN(N__11392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8138),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11385),
            .DIN(N__11384),
            .DOUT(N__11383),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11385),
            .PADOUT(N__11384),
            .PADIN(N__11383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11376),
            .DIN(N__11375),
            .DOUT(N__11374),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11376),
            .PADOUT(N__11375),
            .PADIN(N__11374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4081),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11367),
            .DIN(N__11366),
            .DOUT(N__11365),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11367),
            .PADOUT(N__11366),
            .PADIN(N__11365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9182),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11358),
            .DIN(N__11357),
            .DOUT(N__11356),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11358),
            .PADOUT(N__11357),
            .PADIN(N__11356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11349),
            .DIN(N__11348),
            .DOUT(N__11347),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11349),
            .PADOUT(N__11348),
            .PADIN(N__11347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5750),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11340),
            .DIN(N__11339),
            .DOUT(N__11338),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11340),
            .PADOUT(N__11339),
            .PADIN(N__11338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11331),
            .DIN(N__11330),
            .DOUT(N__11329),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11331),
            .PADOUT(N__11330),
            .PADIN(N__11329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11322),
            .DIN(N__11321),
            .DOUT(N__11320),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11322),
            .PADOUT(N__11321),
            .PADIN(N__11320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11313),
            .DIN(N__11312),
            .DOUT(N__11311),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11313),
            .PADOUT(N__11312),
            .PADIN(N__11311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11304),
            .DIN(N__11303),
            .DOUT(N__11302),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11304),
            .PADOUT(N__11303),
            .PADIN(N__11302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8330),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11295),
            .DIN(N__11294),
            .DOUT(N__11293),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11295),
            .PADOUT(N__11294),
            .PADIN(N__11293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7919),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11286),
            .DIN(N__11285),
            .DOUT(N__11284),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11286),
            .PADOUT(N__11285),
            .PADIN(N__11284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4142),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11277),
            .DIN(N__11276),
            .DOUT(N__11275),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11277),
            .PADOUT(N__11276),
            .PADIN(N__11275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7943),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11268),
            .DIN(N__11267),
            .DOUT(N__11266),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11268),
            .PADOUT(N__11267),
            .PADIN(N__11266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11259),
            .DIN(N__11258),
            .DOUT(N__11257),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11259),
            .PADOUT(N__11258),
            .PADIN(N__11257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11250),
            .DIN(N__11249),
            .DOUT(N__11248),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11250),
            .PADOUT(N__11249),
            .PADIN(N__11248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11241),
            .DIN(N__11240),
            .DOUT(N__11239),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11241),
            .PADOUT(N__11240),
            .PADIN(N__11239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11232),
            .DIN(N__11231),
            .DOUT(N__11230),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11232),
            .PADOUT(N__11231),
            .PADIN(N__11230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7307),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11223),
            .DIN(N__11222),
            .DOUT(N__11221),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11223),
            .PADOUT(N__11222),
            .PADIN(N__11221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11214),
            .DIN(N__11213),
            .DOUT(N__11212),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11214),
            .PADOUT(N__11213),
            .PADIN(N__11212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11205),
            .DIN(N__11204),
            .DOUT(N__11203),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11205),
            .PADOUT(N__11204),
            .PADIN(N__11203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11196),
            .DIN(N__11195),
            .DOUT(N__11194),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11196),
            .PADOUT(N__11195),
            .PADIN(N__11194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4022),
            .DIN0(),
            .DOUT0(N__4121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11187),
            .DIN(N__11186),
            .DOUT(N__11185),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11187),
            .PADOUT(N__11186),
            .PADIN(N__11185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11178),
            .DIN(N__11177),
            .DOUT(N__11176),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11178),
            .PADOUT(N__11177),
            .PADIN(N__11176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11169),
            .DIN(N__11168),
            .DOUT(N__11167),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11169),
            .PADOUT(N__11168),
            .PADIN(N__11167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11160),
            .DIN(N__11159),
            .DOUT(N__11158),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11160),
            .PADOUT(N__11159),
            .PADIN(N__11158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9140),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11151),
            .DIN(N__11150),
            .DOUT(N__11149),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11151),
            .PADOUT(N__11150),
            .PADIN(N__11149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11142),
            .DIN(N__11141),
            .DOUT(N__11140),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11142),
            .PADOUT(N__11141),
            .PADIN(N__11140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11133),
            .DIN(N__11132),
            .DOUT(N__11131),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11133),
            .PADOUT(N__11132),
            .PADIN(N__11131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11124),
            .DIN(N__11123),
            .DOUT(N__11122),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11124),
            .PADOUT(N__11123),
            .PADIN(N__11122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11115),
            .DIN(N__11114),
            .DOUT(N__11113),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11115),
            .PADOUT(N__11114),
            .PADIN(N__11113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11106),
            .DIN(N__11105),
            .DOUT(N__11104),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11106),
            .PADOUT(N__11105),
            .PADIN(N__11104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10082),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11097),
            .DIN(N__11096),
            .DOUT(N__11095),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11097),
            .PADOUT(N__11096),
            .PADIN(N__11095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11088),
            .DIN(N__11087),
            .DOUT(N__11086),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11088),
            .PADOUT(N__11087),
            .PADIN(N__11086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7232),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11079),
            .DIN(N__11078),
            .DOUT(N__11077),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11079),
            .PADOUT(N__11078),
            .PADIN(N__11077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11070),
            .DIN(N__11069),
            .DOUT(N__11068),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11070),
            .PADOUT(N__11069),
            .PADIN(N__11068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11061),
            .DIN(N__11060),
            .DOUT(N__11059),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11061),
            .PADOUT(N__11060),
            .PADIN(N__11059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8939),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11052),
            .DIN(N__11051),
            .DOUT(N__11050),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11052),
            .PADOUT(N__11051),
            .PADIN(N__11050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11043),
            .DIN(N__11042),
            .DOUT(N__11041),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11043),
            .PADOUT(N__11042),
            .PADIN(N__11041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11034),
            .DIN(N__11033),
            .DOUT(N__11032),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11034),
            .PADOUT(N__11033),
            .PADIN(N__11032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4643),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11025),
            .DIN(N__11024),
            .DOUT(N__11023),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11025),
            .PADOUT(N__11024),
            .PADIN(N__11023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9227),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11016),
            .DIN(N__11015),
            .DOUT(N__11014),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11016),
            .PADOUT(N__11015),
            .PADIN(N__11014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4097),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2687 (
            .O(N__10997),
            .I(N__10991));
    InMux I__2686 (
            .O(N__10996),
            .I(N__10988));
    InMux I__2685 (
            .O(N__10995),
            .I(N__10985));
    InMux I__2684 (
            .O(N__10994),
            .I(N__10982));
    LocalMux I__2683 (
            .O(N__10991),
            .I(N__10979));
    LocalMux I__2682 (
            .O(N__10988),
            .I(N__10969));
    LocalMux I__2681 (
            .O(N__10985),
            .I(N__10959));
    LocalMux I__2680 (
            .O(N__10982),
            .I(N__10946));
    Glb2LocalMux I__2679 (
            .O(N__10979),
            .I(N__10853));
    SRMux I__2678 (
            .O(N__10978),
            .I(N__10853));
    SRMux I__2677 (
            .O(N__10977),
            .I(N__10853));
    SRMux I__2676 (
            .O(N__10976),
            .I(N__10853));
    SRMux I__2675 (
            .O(N__10975),
            .I(N__10853));
    SRMux I__2674 (
            .O(N__10974),
            .I(N__10853));
    SRMux I__2673 (
            .O(N__10973),
            .I(N__10853));
    SRMux I__2672 (
            .O(N__10972),
            .I(N__10853));
    Glb2LocalMux I__2671 (
            .O(N__10969),
            .I(N__10853));
    SRMux I__2670 (
            .O(N__10968),
            .I(N__10853));
    SRMux I__2669 (
            .O(N__10967),
            .I(N__10853));
    SRMux I__2668 (
            .O(N__10966),
            .I(N__10853));
    SRMux I__2667 (
            .O(N__10965),
            .I(N__10853));
    SRMux I__2666 (
            .O(N__10964),
            .I(N__10853));
    SRMux I__2665 (
            .O(N__10963),
            .I(N__10853));
    SRMux I__2664 (
            .O(N__10962),
            .I(N__10853));
    Glb2LocalMux I__2663 (
            .O(N__10959),
            .I(N__10853));
    SRMux I__2662 (
            .O(N__10958),
            .I(N__10853));
    SRMux I__2661 (
            .O(N__10957),
            .I(N__10853));
    SRMux I__2660 (
            .O(N__10956),
            .I(N__10853));
    SRMux I__2659 (
            .O(N__10955),
            .I(N__10853));
    SRMux I__2658 (
            .O(N__10954),
            .I(N__10853));
    SRMux I__2657 (
            .O(N__10953),
            .I(N__10853));
    SRMux I__2656 (
            .O(N__10952),
            .I(N__10853));
    SRMux I__2655 (
            .O(N__10951),
            .I(N__10853));
    SRMux I__2654 (
            .O(N__10950),
            .I(N__10853));
    SRMux I__2653 (
            .O(N__10949),
            .I(N__10853));
    Glb2LocalMux I__2652 (
            .O(N__10946),
            .I(N__10853));
    SRMux I__2651 (
            .O(N__10945),
            .I(N__10853));
    SRMux I__2650 (
            .O(N__10944),
            .I(N__10853));
    SRMux I__2649 (
            .O(N__10943),
            .I(N__10853));
    SRMux I__2648 (
            .O(N__10942),
            .I(N__10853));
    SRMux I__2647 (
            .O(N__10941),
            .I(N__10853));
    SRMux I__2646 (
            .O(N__10940),
            .I(N__10853));
    SRMux I__2645 (
            .O(N__10939),
            .I(N__10853));
    SRMux I__2644 (
            .O(N__10938),
            .I(N__10853));
    SRMux I__2643 (
            .O(N__10937),
            .I(N__10853));
    SRMux I__2642 (
            .O(N__10936),
            .I(N__10853));
    SRMux I__2641 (
            .O(N__10935),
            .I(N__10853));
    SRMux I__2640 (
            .O(N__10934),
            .I(N__10853));
    GlobalMux I__2639 (
            .O(N__10853),
            .I(N__10850));
    gio2CtrlBuf I__2638 (
            .O(N__10850),
            .I(RESETn_c_i_g));
    InMux I__2637 (
            .O(N__10847),
            .I(N__10844));
    LocalMux I__2636 (
            .O(N__10844),
            .I(N__10840));
    InMux I__2635 (
            .O(N__10843),
            .I(N__10836));
    Sp12to4 I__2634 (
            .O(N__10840),
            .I(N__10833));
    InMux I__2633 (
            .O(N__10839),
            .I(N__10830));
    LocalMux I__2632 (
            .O(N__10836),
            .I(N__10827));
    Span12Mux_v I__2631 (
            .O(N__10833),
            .I(N__10823));
    LocalMux I__2630 (
            .O(N__10830),
            .I(N__10820));
    Span4Mux_v I__2629 (
            .O(N__10827),
            .I(N__10817));
    InMux I__2628 (
            .O(N__10826),
            .I(N__10813));
    Span12Mux_h I__2627 (
            .O(N__10823),
            .I(N__10810));
    Span12Mux_v I__2626 (
            .O(N__10820),
            .I(N__10807));
    Span4Mux_v I__2625 (
            .O(N__10817),
            .I(N__10804));
    InMux I__2624 (
            .O(N__10816),
            .I(N__10801));
    LocalMux I__2623 (
            .O(N__10813),
            .I(N__10798));
    Odrv12 I__2622 (
            .O(N__10810),
            .I(REG_CYCLEm));
    Odrv12 I__2621 (
            .O(N__10807),
            .I(REG_CYCLEm));
    Odrv4 I__2620 (
            .O(N__10804),
            .I(REG_CYCLEm));
    LocalMux I__2619 (
            .O(N__10801),
            .I(REG_CYCLEm));
    Odrv4 I__2618 (
            .O(N__10798),
            .I(REG_CYCLEm));
    InMux I__2617 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__2616 (
            .O(N__10784),
            .I(N__10781));
    Span4Mux_h I__2615 (
            .O(N__10781),
            .I(N__10777));
    InMux I__2614 (
            .O(N__10780),
            .I(N__10773));
    Span4Mux_h I__2613 (
            .O(N__10777),
            .I(N__10769));
    InMux I__2612 (
            .O(N__10776),
            .I(N__10765));
    LocalMux I__2611 (
            .O(N__10773),
            .I(N__10762));
    InMux I__2610 (
            .O(N__10772),
            .I(N__10759));
    Span4Mux_h I__2609 (
            .O(N__10769),
            .I(N__10756));
    InMux I__2608 (
            .O(N__10768),
            .I(N__10753));
    LocalMux I__2607 (
            .O(N__10765),
            .I(N__10750));
    Sp12to4 I__2606 (
            .O(N__10762),
            .I(N__10745));
    LocalMux I__2605 (
            .O(N__10759),
            .I(N__10745));
    Span4Mux_h I__2604 (
            .O(N__10756),
            .I(N__10740));
    LocalMux I__2603 (
            .O(N__10753),
            .I(N__10740));
    Span12Mux_h I__2602 (
            .O(N__10750),
            .I(N__10737));
    Span12Mux_v I__2601 (
            .O(N__10745),
            .I(N__10734));
    Span4Mux_h I__2600 (
            .O(N__10740),
            .I(N__10731));
    Span12Mux_v I__2599 (
            .O(N__10737),
            .I(N__10728));
    Span12Mux_h I__2598 (
            .O(N__10734),
            .I(N__10725));
    Span4Mux_v I__2597 (
            .O(N__10731),
            .I(N__10722));
    Odrv12 I__2596 (
            .O(N__10728),
            .I(CASUn_c));
    Odrv12 I__2595 (
            .O(N__10725),
            .I(CASUn_c));
    Odrv4 I__2594 (
            .O(N__10722),
            .I(CASUn_c));
    InMux I__2593 (
            .O(N__10715),
            .I(N__10711));
    InMux I__2592 (
            .O(N__10714),
            .I(N__10708));
    LocalMux I__2591 (
            .O(N__10711),
            .I(N__10705));
    LocalMux I__2590 (
            .O(N__10708),
            .I(N__10702));
    Span4Mux_v I__2589 (
            .O(N__10705),
            .I(N__10695));
    Span4Mux_v I__2588 (
            .O(N__10702),
            .I(N__10695));
    InMux I__2587 (
            .O(N__10701),
            .I(N__10692));
    InMux I__2586 (
            .O(N__10700),
            .I(N__10689));
    Sp12to4 I__2585 (
            .O(N__10695),
            .I(N__10685));
    LocalMux I__2584 (
            .O(N__10692),
            .I(N__10682));
    LocalMux I__2583 (
            .O(N__10689),
            .I(N__10679));
    InMux I__2582 (
            .O(N__10688),
            .I(N__10676));
    Span12Mux_h I__2581 (
            .O(N__10685),
            .I(N__10673));
    Span12Mux_v I__2580 (
            .O(N__10682),
            .I(N__10670));
    Span12Mux_v I__2579 (
            .O(N__10679),
            .I(N__10667));
    LocalMux I__2578 (
            .O(N__10676),
            .I(N__10664));
    Span12Mux_v I__2577 (
            .O(N__10673),
            .I(N__10659));
    Span12Mux_h I__2576 (
            .O(N__10670),
            .I(N__10659));
    Span12Mux_h I__2575 (
            .O(N__10667),
            .I(N__10654));
    Span12Mux_v I__2574 (
            .O(N__10664),
            .I(N__10654));
    Odrv12 I__2573 (
            .O(N__10659),
            .I(CASLn_c));
    Odrv12 I__2572 (
            .O(N__10654),
            .I(CASLn_c));
    IoInMux I__2571 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__2570 (
            .O(N__10646),
            .I(N__10643));
    Span4Mux_s3_v I__2569 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_v I__2568 (
            .O(N__10640),
            .I(N__10637));
    Odrv4 I__2567 (
            .O(N__10637),
            .I(DRDENn_c));
    InMux I__2566 (
            .O(N__10634),
            .I(N__10629));
    InMux I__2565 (
            .O(N__10633),
            .I(N__10625));
    InMux I__2564 (
            .O(N__10632),
            .I(N__10622));
    LocalMux I__2563 (
            .O(N__10629),
            .I(N__10616));
    InMux I__2562 (
            .O(N__10628),
            .I(N__10613));
    LocalMux I__2561 (
            .O(N__10625),
            .I(N__10610));
    LocalMux I__2560 (
            .O(N__10622),
            .I(N__10607));
    InMux I__2559 (
            .O(N__10621),
            .I(N__10602));
    InMux I__2558 (
            .O(N__10620),
            .I(N__10602));
    InMux I__2557 (
            .O(N__10619),
            .I(N__10599));
    Span4Mux_v I__2556 (
            .O(N__10616),
            .I(N__10596));
    LocalMux I__2555 (
            .O(N__10613),
            .I(N__10593));
    Span4Mux_v I__2554 (
            .O(N__10610),
            .I(N__10590));
    Span4Mux_v I__2553 (
            .O(N__10607),
            .I(N__10587));
    LocalMux I__2552 (
            .O(N__10602),
            .I(N__10584));
    LocalMux I__2551 (
            .O(N__10599),
            .I(N__10580));
    Span4Mux_v I__2550 (
            .O(N__10596),
            .I(N__10575));
    Span4Mux_v I__2549 (
            .O(N__10593),
            .I(N__10575));
    Span4Mux_v I__2548 (
            .O(N__10590),
            .I(N__10568));
    Span4Mux_v I__2547 (
            .O(N__10587),
            .I(N__10568));
    Span4Mux_v I__2546 (
            .O(N__10584),
            .I(N__10568));
    InMux I__2545 (
            .O(N__10583),
            .I(N__10565));
    Span12Mux_v I__2544 (
            .O(N__10580),
            .I(N__10562));
    Sp12to4 I__2543 (
            .O(N__10575),
            .I(N__10555));
    Sp12to4 I__2542 (
            .O(N__10568),
            .I(N__10555));
    LocalMux I__2541 (
            .O(N__10565),
            .I(N__10555));
    Span12Mux_h I__2540 (
            .O(N__10562),
            .I(N__10552));
    Span12Mux_h I__2539 (
            .O(N__10555),
            .I(N__10549));
    Odrv12 I__2538 (
            .O(N__10552),
            .I(A_c_1));
    Odrv12 I__2537 (
            .O(N__10549),
            .I(A_c_1));
    InMux I__2536 (
            .O(N__10544),
            .I(N__10541));
    LocalMux I__2535 (
            .O(N__10541),
            .I(N__10535));
    InMux I__2534 (
            .O(N__10540),
            .I(N__10532));
    InMux I__2533 (
            .O(N__10539),
            .I(N__10529));
    CascadeMux I__2532 (
            .O(N__10538),
            .I(N__10525));
    Span4Mux_v I__2531 (
            .O(N__10535),
            .I(N__10521));
    LocalMux I__2530 (
            .O(N__10532),
            .I(N__10518));
    LocalMux I__2529 (
            .O(N__10529),
            .I(N__10515));
    InMux I__2528 (
            .O(N__10528),
            .I(N__10510));
    InMux I__2527 (
            .O(N__10525),
            .I(N__10510));
    InMux I__2526 (
            .O(N__10524),
            .I(N__10507));
    Span4Mux_h I__2525 (
            .O(N__10521),
            .I(N__10502));
    Span4Mux_v I__2524 (
            .O(N__10518),
            .I(N__10502));
    Span4Mux_v I__2523 (
            .O(N__10515),
            .I(N__10495));
    LocalMux I__2522 (
            .O(N__10510),
            .I(N__10495));
    LocalMux I__2521 (
            .O(N__10507),
            .I(N__10495));
    Span4Mux_v I__2520 (
            .O(N__10502),
            .I(N__10492));
    Span4Mux_h I__2519 (
            .O(N__10495),
            .I(N__10489));
    Span4Mux_v I__2518 (
            .O(N__10492),
            .I(N__10486));
    Span4Mux_v I__2517 (
            .O(N__10489),
            .I(N__10483));
    Sp12to4 I__2516 (
            .O(N__10486),
            .I(N__10478));
    Sp12to4 I__2515 (
            .O(N__10483),
            .I(N__10478));
    Span12Mux_h I__2514 (
            .O(N__10478),
            .I(N__10475));
    Odrv12 I__2513 (
            .O(N__10475),
            .I(SIZ_c_0));
    CascadeMux I__2512 (
            .O(N__10472),
            .I(N__10469));
    InMux I__2511 (
            .O(N__10469),
            .I(N__10465));
    InMux I__2510 (
            .O(N__10468),
            .I(N__10462));
    LocalMux I__2509 (
            .O(N__10465),
            .I(N__10454));
    LocalMux I__2508 (
            .O(N__10462),
            .I(N__10454));
    CascadeMux I__2507 (
            .O(N__10461),
            .I(N__10448));
    InMux I__2506 (
            .O(N__10460),
            .I(N__10443));
    InMux I__2505 (
            .O(N__10459),
            .I(N__10443));
    Span4Mux_v I__2504 (
            .O(N__10454),
            .I(N__10440));
    InMux I__2503 (
            .O(N__10453),
            .I(N__10437));
    InMux I__2502 (
            .O(N__10452),
            .I(N__10432));
    InMux I__2501 (
            .O(N__10451),
            .I(N__10432));
    InMux I__2500 (
            .O(N__10448),
            .I(N__10429));
    LocalMux I__2499 (
            .O(N__10443),
            .I(N__10426));
    Span4Mux_v I__2498 (
            .O(N__10440),
            .I(N__10423));
    LocalMux I__2497 (
            .O(N__10437),
            .I(N__10416));
    LocalMux I__2496 (
            .O(N__10432),
            .I(N__10416));
    LocalMux I__2495 (
            .O(N__10429),
            .I(N__10416));
    Sp12to4 I__2494 (
            .O(N__10426),
            .I(N__10413));
    Span4Mux_v I__2493 (
            .O(N__10423),
            .I(N__10410));
    Sp12to4 I__2492 (
            .O(N__10416),
            .I(N__10407));
    Span12Mux_v I__2491 (
            .O(N__10413),
            .I(N__10404));
    Sp12to4 I__2490 (
            .O(N__10410),
            .I(N__10399));
    Span12Mux_v I__2489 (
            .O(N__10407),
            .I(N__10399));
    Span12Mux_h I__2488 (
            .O(N__10404),
            .I(N__10396));
    Span12Mux_h I__2487 (
            .O(N__10399),
            .I(N__10393));
    Odrv12 I__2486 (
            .O(N__10396),
            .I(SIZ_c_1));
    Odrv12 I__2485 (
            .O(N__10393),
            .I(SIZ_c_1));
    IoInMux I__2484 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__2483 (
            .O(N__10385),
            .I(N__10382));
    Span4Mux_s2_v I__2482 (
            .O(N__10382),
            .I(N__10379));
    Span4Mux_v I__2481 (
            .O(N__10379),
            .I(N__10376));
    Odrv4 I__2480 (
            .O(N__10376),
            .I(N_303_i));
    InMux I__2479 (
            .O(N__10373),
            .I(N__10370));
    LocalMux I__2478 (
            .O(N__10370),
            .I(N__10367));
    Odrv4 I__2477 (
            .O(N__10367),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2476 (
            .O(N__10364),
            .I(N__10358));
    InMux I__2475 (
            .O(N__10363),
            .I(N__10355));
    InMux I__2474 (
            .O(N__10362),
            .I(N__10352));
    InMux I__2473 (
            .O(N__10361),
            .I(N__10349));
    LocalMux I__2472 (
            .O(N__10358),
            .I(N__10340));
    LocalMux I__2471 (
            .O(N__10355),
            .I(N__10340));
    LocalMux I__2470 (
            .O(N__10352),
            .I(N__10340));
    LocalMux I__2469 (
            .O(N__10349),
            .I(N__10340));
    Span4Mux_v I__2468 (
            .O(N__10340),
            .I(N__10337));
    Sp12to4 I__2467 (
            .O(N__10337),
            .I(N__10334));
    Span12Mux_h I__2466 (
            .O(N__10334),
            .I(N__10331));
    Odrv12 I__2465 (
            .O(N__10331),
            .I(DRA_c_8));
    InMux I__2464 (
            .O(N__10328),
            .I(N__10325));
    LocalMux I__2463 (
            .O(N__10325),
            .I(N__10322));
    Span4Mux_h I__2462 (
            .O(N__10322),
            .I(N__10319));
    Odrv4 I__2461 (
            .O(N__10319),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2460 (
            .O(N__10316),
            .I(N__10313));
    LocalMux I__2459 (
            .O(N__10313),
            .I(N__10310));
    Span12Mux_v I__2458 (
            .O(N__10310),
            .I(N__10307));
    Odrv12 I__2457 (
            .O(N__10307),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2456 (
            .O(N__10304),
            .I(N__10301));
    LocalMux I__2455 (
            .O(N__10301),
            .I(N__10296));
    InMux I__2454 (
            .O(N__10300),
            .I(N__10293));
    InMux I__2453 (
            .O(N__10299),
            .I(N__10290));
    Span4Mux_v I__2452 (
            .O(N__10296),
            .I(N__10285));
    LocalMux I__2451 (
            .O(N__10293),
            .I(N__10285));
    LocalMux I__2450 (
            .O(N__10290),
            .I(N__10282));
    Span4Mux_v I__2449 (
            .O(N__10285),
            .I(N__10278));
    Span4Mux_v I__2448 (
            .O(N__10282),
            .I(N__10275));
    InMux I__2447 (
            .O(N__10281),
            .I(N__10272));
    Sp12to4 I__2446 (
            .O(N__10278),
            .I(N__10269));
    Sp12to4 I__2445 (
            .O(N__10275),
            .I(N__10264));
    LocalMux I__2444 (
            .O(N__10272),
            .I(N__10264));
    Span12Mux_v I__2443 (
            .O(N__10269),
            .I(N__10261));
    Span12Mux_h I__2442 (
            .O(N__10264),
            .I(N__10258));
    Span12Mux_h I__2441 (
            .O(N__10261),
            .I(N__10253));
    Span12Mux_v I__2440 (
            .O(N__10258),
            .I(N__10253));
    Odrv12 I__2439 (
            .O(N__10253),
            .I(DRA_c_1));
    InMux I__2438 (
            .O(N__10250),
            .I(N__10247));
    LocalMux I__2437 (
            .O(N__10247),
            .I(N__10243));
    InMux I__2436 (
            .O(N__10246),
            .I(N__10240));
    Span4Mux_h I__2435 (
            .O(N__10243),
            .I(N__10235));
    LocalMux I__2434 (
            .O(N__10240),
            .I(N__10235));
    Sp12to4 I__2433 (
            .O(N__10235),
            .I(N__10232));
    Span12Mux_v I__2432 (
            .O(N__10232),
            .I(N__10229));
    Span12Mux_h I__2431 (
            .O(N__10229),
            .I(N__10226));
    Odrv12 I__2430 (
            .O(N__10226),
            .I(DRA_c_0));
    InMux I__2429 (
            .O(N__10223),
            .I(N__10220));
    LocalMux I__2428 (
            .O(N__10220),
            .I(N__10217));
    Odrv4 I__2427 (
            .O(N__10217),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2426 (
            .O(N__10214),
            .I(N__10211));
    LocalMux I__2425 (
            .O(N__10211),
            .I(N__10207));
    CascadeMux I__2424 (
            .O(N__10210),
            .I(N__10204));
    Span4Mux_h I__2423 (
            .O(N__10207),
            .I(N__10201));
    InMux I__2422 (
            .O(N__10204),
            .I(N__10198));
    Sp12to4 I__2421 (
            .O(N__10201),
            .I(N__10193));
    LocalMux I__2420 (
            .O(N__10198),
            .I(N__10193));
    Span12Mux_v I__2419 (
            .O(N__10193),
            .I(N__10189));
    InMux I__2418 (
            .O(N__10192),
            .I(N__10186));
    Odrv12 I__2417 (
            .O(N__10189),
            .I(DS_ENm));
    LocalMux I__2416 (
            .O(N__10186),
            .I(DS_ENm));
    CascadeMux I__2415 (
            .O(N__10181),
            .I(N__10171));
    InMux I__2414 (
            .O(N__10180),
            .I(N__10165));
    InMux I__2413 (
            .O(N__10179),
            .I(N__10165));
    InMux I__2412 (
            .O(N__10178),
            .I(N__10162));
    InMux I__2411 (
            .O(N__10177),
            .I(N__10158));
    InMux I__2410 (
            .O(N__10176),
            .I(N__10155));
    InMux I__2409 (
            .O(N__10175),
            .I(N__10150));
    InMux I__2408 (
            .O(N__10174),
            .I(N__10150));
    InMux I__2407 (
            .O(N__10171),
            .I(N__10147));
    CascadeMux I__2406 (
            .O(N__10170),
            .I(N__10144));
    LocalMux I__2405 (
            .O(N__10165),
            .I(N__10141));
    LocalMux I__2404 (
            .O(N__10162),
            .I(N__10138));
    InMux I__2403 (
            .O(N__10161),
            .I(N__10135));
    LocalMux I__2402 (
            .O(N__10158),
            .I(N__10132));
    LocalMux I__2401 (
            .O(N__10155),
            .I(N__10125));
    LocalMux I__2400 (
            .O(N__10150),
            .I(N__10125));
    LocalMux I__2399 (
            .O(N__10147),
            .I(N__10125));
    InMux I__2398 (
            .O(N__10144),
            .I(N__10122));
    Span4Mux_v I__2397 (
            .O(N__10141),
            .I(N__10117));
    Span4Mux_v I__2396 (
            .O(N__10138),
            .I(N__10117));
    LocalMux I__2395 (
            .O(N__10135),
            .I(N__10114));
    Span4Mux_v I__2394 (
            .O(N__10132),
            .I(N__10109));
    Span4Mux_v I__2393 (
            .O(N__10125),
            .I(N__10109));
    LocalMux I__2392 (
            .O(N__10122),
            .I(N__10106));
    Sp12to4 I__2391 (
            .O(N__10117),
            .I(N__10101));
    Span12Mux_v I__2390 (
            .O(N__10114),
            .I(N__10101));
    Sp12to4 I__2389 (
            .O(N__10109),
            .I(N__10098));
    Span4Mux_v I__2388 (
            .O(N__10106),
            .I(N__10095));
    Span12Mux_h I__2387 (
            .O(N__10101),
            .I(N__10092));
    Span12Mux_h I__2386 (
            .O(N__10098),
            .I(N__10087));
    Sp12to4 I__2385 (
            .O(N__10095),
            .I(N__10087));
    Odrv12 I__2384 (
            .O(N__10092),
            .I(A_c_0));
    Odrv12 I__2383 (
            .O(N__10087),
            .I(A_c_0));
    IoInMux I__2382 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__2381 (
            .O(N__10079),
            .I(N__10076));
    Span4Mux_s3_v I__2380 (
            .O(N__10076),
            .I(N__10073));
    Span4Mux_h I__2379 (
            .O(N__10073),
            .I(N__10070));
    Span4Mux_h I__2378 (
            .O(N__10070),
            .I(N__10067));
    Odrv4 I__2377 (
            .O(N__10067),
            .I(N_337_i));
    InMux I__2376 (
            .O(N__10064),
            .I(N__10061));
    LocalMux I__2375 (
            .O(N__10061),
            .I(N__10058));
    Span4Mux_v I__2374 (
            .O(N__10058),
            .I(N__10052));
    InMux I__2373 (
            .O(N__10057),
            .I(N__10049));
    InMux I__2372 (
            .O(N__10056),
            .I(N__10046));
    InMux I__2371 (
            .O(N__10055),
            .I(N__10043));
    Span4Mux_v I__2370 (
            .O(N__10052),
            .I(N__10036));
    LocalMux I__2369 (
            .O(N__10049),
            .I(N__10036));
    LocalMux I__2368 (
            .O(N__10046),
            .I(N__10036));
    LocalMux I__2367 (
            .O(N__10043),
            .I(N__10033));
    Span4Mux_h I__2366 (
            .O(N__10036),
            .I(N__10028));
    Span4Mux_v I__2365 (
            .O(N__10033),
            .I(N__10028));
    Span4Mux_v I__2364 (
            .O(N__10028),
            .I(N__10025));
    Sp12to4 I__2363 (
            .O(N__10025),
            .I(N__10022));
    Odrv12 I__2362 (
            .O(N__10022),
            .I(DRA_c_6));
    CascadeMux I__2361 (
            .O(N__10019),
            .I(N__10016));
    InMux I__2360 (
            .O(N__10016),
            .I(N__10011));
    InMux I__2359 (
            .O(N__10015),
            .I(N__10008));
    InMux I__2358 (
            .O(N__10014),
            .I(N__10005));
    LocalMux I__2357 (
            .O(N__10011),
            .I(N__9997));
    LocalMux I__2356 (
            .O(N__10008),
            .I(N__9997));
    LocalMux I__2355 (
            .O(N__10005),
            .I(N__9997));
    InMux I__2354 (
            .O(N__10004),
            .I(N__9994));
    Span4Mux_v I__2353 (
            .O(N__9997),
            .I(N__9991));
    LocalMux I__2352 (
            .O(N__9994),
            .I(N__9988));
    Sp12to4 I__2351 (
            .O(N__9991),
            .I(N__9983));
    Span12Mux_v I__2350 (
            .O(N__9988),
            .I(N__9983));
    Span12Mux_h I__2349 (
            .O(N__9983),
            .I(N__9980));
    Odrv12 I__2348 (
            .O(N__9980),
            .I(DRA_c_7));
    InMux I__2347 (
            .O(N__9977),
            .I(N__9974));
    LocalMux I__2346 (
            .O(N__9974),
            .I(N__9971));
    Span4Mux_h I__2345 (
            .O(N__9971),
            .I(N__9968));
    Odrv4 I__2344 (
            .O(N__9968),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2343 (
            .O(N__9965),
            .I(N__9960));
    CascadeMux I__2342 (
            .O(N__9964),
            .I(N__9954));
    CascadeMux I__2341 (
            .O(N__9963),
            .I(N__9951));
    LocalMux I__2340 (
            .O(N__9960),
            .I(N__9941));
    InMux I__2339 (
            .O(N__9959),
            .I(N__9936));
    InMux I__2338 (
            .O(N__9958),
            .I(N__9936));
    InMux I__2337 (
            .O(N__9957),
            .I(N__9933));
    InMux I__2336 (
            .O(N__9954),
            .I(N__9926));
    InMux I__2335 (
            .O(N__9951),
            .I(N__9926));
    InMux I__2334 (
            .O(N__9950),
            .I(N__9926));
    InMux I__2333 (
            .O(N__9949),
            .I(N__9921));
    InMux I__2332 (
            .O(N__9948),
            .I(N__9921));
    InMux I__2331 (
            .O(N__9947),
            .I(N__9918));
    InMux I__2330 (
            .O(N__9946),
            .I(N__9915));
    InMux I__2329 (
            .O(N__9945),
            .I(N__9912));
    InMux I__2328 (
            .O(N__9944),
            .I(N__9908));
    Span4Mux_v I__2327 (
            .O(N__9941),
            .I(N__9900));
    LocalMux I__2326 (
            .O(N__9936),
            .I(N__9887));
    LocalMux I__2325 (
            .O(N__9933),
            .I(N__9887));
    LocalMux I__2324 (
            .O(N__9926),
            .I(N__9887));
    LocalMux I__2323 (
            .O(N__9921),
            .I(N__9887));
    LocalMux I__2322 (
            .O(N__9918),
            .I(N__9887));
    LocalMux I__2321 (
            .O(N__9915),
            .I(N__9887));
    LocalMux I__2320 (
            .O(N__9912),
            .I(N__9884));
    InMux I__2319 (
            .O(N__9911),
            .I(N__9881));
    LocalMux I__2318 (
            .O(N__9908),
            .I(N__9878));
    InMux I__2317 (
            .O(N__9907),
            .I(N__9873));
    InMux I__2316 (
            .O(N__9906),
            .I(N__9873));
    InMux I__2315 (
            .O(N__9905),
            .I(N__9870));
    InMux I__2314 (
            .O(N__9904),
            .I(N__9867));
    InMux I__2313 (
            .O(N__9903),
            .I(N__9864));
    Span4Mux_h I__2312 (
            .O(N__9900),
            .I(N__9857));
    Span4Mux_v I__2311 (
            .O(N__9887),
            .I(N__9857));
    Span4Mux_v I__2310 (
            .O(N__9884),
            .I(N__9852));
    LocalMux I__2309 (
            .O(N__9881),
            .I(N__9852));
    Span4Mux_v I__2308 (
            .O(N__9878),
            .I(N__9841));
    LocalMux I__2307 (
            .O(N__9873),
            .I(N__9841));
    LocalMux I__2306 (
            .O(N__9870),
            .I(N__9841));
    LocalMux I__2305 (
            .O(N__9867),
            .I(N__9841));
    LocalMux I__2304 (
            .O(N__9864),
            .I(N__9841));
    InMux I__2303 (
            .O(N__9863),
            .I(N__9838));
    InMux I__2302 (
            .O(N__9862),
            .I(N__9835));
    Span4Mux_h I__2301 (
            .O(N__9857),
            .I(N__9830));
    Span4Mux_v I__2300 (
            .O(N__9852),
            .I(N__9830));
    Span4Mux_v I__2299 (
            .O(N__9841),
            .I(N__9827));
    LocalMux I__2298 (
            .O(N__9838),
            .I(N__9822));
    LocalMux I__2297 (
            .O(N__9835),
            .I(N__9822));
    Sp12to4 I__2296 (
            .O(N__9830),
            .I(N__9817));
    Sp12to4 I__2295 (
            .O(N__9827),
            .I(N__9817));
    Span12Mux_h I__2294 (
            .O(N__9822),
            .I(N__9814));
    Span12Mux_h I__2293 (
            .O(N__9817),
            .I(N__9811));
    Span12Mux_v I__2292 (
            .O(N__9814),
            .I(N__9808));
    Span12Mux_v I__2291 (
            .O(N__9811),
            .I(N__9805));
    Odrv12 I__2290 (
            .O(N__9808),
            .I(AGNUS_REV_c));
    Odrv12 I__2289 (
            .O(N__9805),
            .I(AGNUS_REV_c));
    InMux I__2288 (
            .O(N__9800),
            .I(N__9797));
    LocalMux I__2287 (
            .O(N__9797),
            .I(N__9794));
    Span4Mux_v I__2286 (
            .O(N__9794),
            .I(N__9791));
    Sp12to4 I__2285 (
            .O(N__9791),
            .I(N__9788));
    Odrv12 I__2284 (
            .O(N__9788),
            .I(RAS0n_c));
    InMux I__2283 (
            .O(N__9785),
            .I(N__9780));
    InMux I__2282 (
            .O(N__9784),
            .I(N__9777));
    CascadeMux I__2281 (
            .O(N__9783),
            .I(N__9774));
    LocalMux I__2280 (
            .O(N__9780),
            .I(N__9769));
    LocalMux I__2279 (
            .O(N__9777),
            .I(N__9769));
    InMux I__2278 (
            .O(N__9774),
            .I(N__9766));
    Span4Mux_v I__2277 (
            .O(N__9769),
            .I(N__9762));
    LocalMux I__2276 (
            .O(N__9766),
            .I(N__9759));
    InMux I__2275 (
            .O(N__9765),
            .I(N__9756));
    Span4Mux_v I__2274 (
            .O(N__9762),
            .I(N__9753));
    Span4Mux_v I__2273 (
            .O(N__9759),
            .I(N__9750));
    LocalMux I__2272 (
            .O(N__9756),
            .I(N__9747));
    Sp12to4 I__2271 (
            .O(N__9753),
            .I(N__9742));
    Sp12to4 I__2270 (
            .O(N__9750),
            .I(N__9742));
    Sp12to4 I__2269 (
            .O(N__9747),
            .I(N__9739));
    Span12Mux_h I__2268 (
            .O(N__9742),
            .I(N__9736));
    Span12Mux_v I__2267 (
            .O(N__9739),
            .I(N__9733));
    Span12Mux_v I__2266 (
            .O(N__9736),
            .I(N__9730));
    Span12Mux_v I__2265 (
            .O(N__9733),
            .I(N__9727));
    Odrv12 I__2264 (
            .O(N__9730),
            .I(DRA_c_9));
    Odrv12 I__2263 (
            .O(N__9727),
            .I(DRA_c_9));
    InMux I__2262 (
            .O(N__9722),
            .I(N__9719));
    LocalMux I__2261 (
            .O(N__9719),
            .I(N__9716));
    Odrv4 I__2260 (
            .O(N__9716),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2259 (
            .O(N__9713),
            .I(N__9692));
    ClkMux I__2258 (
            .O(N__9712),
            .I(N__9692));
    ClkMux I__2257 (
            .O(N__9711),
            .I(N__9692));
    ClkMux I__2256 (
            .O(N__9710),
            .I(N__9692));
    ClkMux I__2255 (
            .O(N__9709),
            .I(N__9692));
    ClkMux I__2254 (
            .O(N__9708),
            .I(N__9692));
    ClkMux I__2253 (
            .O(N__9707),
            .I(N__9692));
    GlobalMux I__2252 (
            .O(N__9692),
            .I(N__9689));
    gio2CtrlBuf I__2251 (
            .O(N__9689),
            .I(C3_c_g));
    CEMux I__2250 (
            .O(N__9686),
            .I(N__9644));
    CEMux I__2249 (
            .O(N__9685),
            .I(N__9644));
    CEMux I__2248 (
            .O(N__9684),
            .I(N__9644));
    CEMux I__2247 (
            .O(N__9683),
            .I(N__9644));
    CEMux I__2246 (
            .O(N__9682),
            .I(N__9644));
    CEMux I__2245 (
            .O(N__9681),
            .I(N__9644));
    CEMux I__2244 (
            .O(N__9680),
            .I(N__9644));
    CEMux I__2243 (
            .O(N__9679),
            .I(N__9644));
    CEMux I__2242 (
            .O(N__9678),
            .I(N__9644));
    CEMux I__2241 (
            .O(N__9677),
            .I(N__9644));
    CEMux I__2240 (
            .O(N__9676),
            .I(N__9644));
    CEMux I__2239 (
            .O(N__9675),
            .I(N__9644));
    CEMux I__2238 (
            .O(N__9674),
            .I(N__9644));
    CEMux I__2237 (
            .O(N__9673),
            .I(N__9644));
    GlobalMux I__2236 (
            .O(N__9644),
            .I(N__9641));
    gio2CtrlBuf I__2235 (
            .O(N__9641),
            .I(DBRn_c_i_0_g));
    InMux I__2234 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__2233 (
            .O(N__9635),
            .I(N__9632));
    Odrv4 I__2232 (
            .O(N__9632),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2231 (
            .O(N__9629),
            .I(N__9626));
    LocalMux I__2230 (
            .O(N__9626),
            .I(N__9623));
    Odrv4 I__2229 (
            .O(N__9623),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2228 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__2227 (
            .O(N__9617),
            .I(N__9611));
    InMux I__2226 (
            .O(N__9616),
            .I(N__9606));
    InMux I__2225 (
            .O(N__9615),
            .I(N__9606));
    InMux I__2224 (
            .O(N__9614),
            .I(N__9603));
    Span4Mux_h I__2223 (
            .O(N__9611),
            .I(N__9598));
    LocalMux I__2222 (
            .O(N__9606),
            .I(N__9598));
    LocalMux I__2221 (
            .O(N__9603),
            .I(N__9593));
    Sp12to4 I__2220 (
            .O(N__9598),
            .I(N__9593));
    Span12Mux_v I__2219 (
            .O(N__9593),
            .I(N__9590));
    Span12Mux_h I__2218 (
            .O(N__9590),
            .I(N__9587));
    Odrv12 I__2217 (
            .O(N__9587),
            .I(DRA_c_5));
    InMux I__2216 (
            .O(N__9584),
            .I(N__9578));
    InMux I__2215 (
            .O(N__9583),
            .I(N__9575));
    InMux I__2214 (
            .O(N__9582),
            .I(N__9572));
    InMux I__2213 (
            .O(N__9581),
            .I(N__9569));
    LocalMux I__2212 (
            .O(N__9578),
            .I(N__9564));
    LocalMux I__2211 (
            .O(N__9575),
            .I(N__9564));
    LocalMux I__2210 (
            .O(N__9572),
            .I(N__9561));
    LocalMux I__2209 (
            .O(N__9569),
            .I(N__9558));
    Span4Mux_v I__2208 (
            .O(N__9564),
            .I(N__9555));
    Span4Mux_v I__2207 (
            .O(N__9561),
            .I(N__9552));
    Span4Mux_h I__2206 (
            .O(N__9558),
            .I(N__9549));
    Span4Mux_v I__2205 (
            .O(N__9555),
            .I(N__9546));
    Span4Mux_v I__2204 (
            .O(N__9552),
            .I(N__9543));
    Sp12to4 I__2203 (
            .O(N__9549),
            .I(N__9540));
    Sp12to4 I__2202 (
            .O(N__9546),
            .I(N__9537));
    Sp12to4 I__2201 (
            .O(N__9543),
            .I(N__9532));
    Span12Mux_v I__2200 (
            .O(N__9540),
            .I(N__9532));
    Span12Mux_h I__2199 (
            .O(N__9537),
            .I(N__9529));
    Span12Mux_h I__2198 (
            .O(N__9532),
            .I(N__9526));
    Odrv12 I__2197 (
            .O(N__9529),
            .I(DRA_c_4));
    Odrv12 I__2196 (
            .O(N__9526),
            .I(DRA_c_4));
    InMux I__2195 (
            .O(N__9521),
            .I(N__9518));
    LocalMux I__2194 (
            .O(N__9518),
            .I(N__9515));
    Odrv12 I__2193 (
            .O(N__9515),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2192 (
            .O(N__9512),
            .I(N__9509));
    LocalMux I__2191 (
            .O(N__9509),
            .I(N__9506));
    Span4Mux_h I__2190 (
            .O(N__9506),
            .I(N__9503));
    Span4Mux_h I__2189 (
            .O(N__9503),
            .I(N__9500));
    Odrv4 I__2188 (
            .O(N__9500),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2187 (
            .O(N__9497),
            .I(N__9493));
    InMux I__2186 (
            .O(N__9496),
            .I(N__9490));
    LocalMux I__2185 (
            .O(N__9493),
            .I(N__9487));
    LocalMux I__2184 (
            .O(N__9490),
            .I(N__9484));
    Span4Mux_h I__2183 (
            .O(N__9487),
            .I(N__9479));
    Span4Mux_v I__2182 (
            .O(N__9484),
            .I(N__9479));
    Odrv4 I__2181 (
            .O(N__9479),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0 ));
    CascadeMux I__2180 (
            .O(N__9476),
            .I(N__9471));
    CascadeMux I__2179 (
            .O(N__9475),
            .I(N__9465));
    CascadeMux I__2178 (
            .O(N__9474),
            .I(N__9462));
    InMux I__2177 (
            .O(N__9471),
            .I(N__9457));
    CascadeMux I__2176 (
            .O(N__9470),
            .I(N__9449));
    CascadeMux I__2175 (
            .O(N__9469),
            .I(N__9444));
    InMux I__2174 (
            .O(N__9468),
            .I(N__9437));
    InMux I__2173 (
            .O(N__9465),
            .I(N__9434));
    InMux I__2172 (
            .O(N__9462),
            .I(N__9431));
    InMux I__2171 (
            .O(N__9461),
            .I(N__9426));
    InMux I__2170 (
            .O(N__9460),
            .I(N__9426));
    LocalMux I__2169 (
            .O(N__9457),
            .I(N__9423));
    InMux I__2168 (
            .O(N__9456),
            .I(N__9420));
    InMux I__2167 (
            .O(N__9455),
            .I(N__9417));
    InMux I__2166 (
            .O(N__9454),
            .I(N__9414));
    InMux I__2165 (
            .O(N__9453),
            .I(N__9410));
    InMux I__2164 (
            .O(N__9452),
            .I(N__9405));
    InMux I__2163 (
            .O(N__9449),
            .I(N__9405));
    InMux I__2162 (
            .O(N__9448),
            .I(N__9400));
    InMux I__2161 (
            .O(N__9447),
            .I(N__9400));
    InMux I__2160 (
            .O(N__9444),
            .I(N__9397));
    InMux I__2159 (
            .O(N__9443),
            .I(N__9392));
    InMux I__2158 (
            .O(N__9442),
            .I(N__9392));
    InMux I__2157 (
            .O(N__9441),
            .I(N__9389));
    InMux I__2156 (
            .O(N__9440),
            .I(N__9386));
    LocalMux I__2155 (
            .O(N__9437),
            .I(N__9380));
    LocalMux I__2154 (
            .O(N__9434),
            .I(N__9380));
    LocalMux I__2153 (
            .O(N__9431),
            .I(N__9375));
    LocalMux I__2152 (
            .O(N__9426),
            .I(N__9375));
    Span4Mux_v I__2151 (
            .O(N__9423),
            .I(N__9368));
    LocalMux I__2150 (
            .O(N__9420),
            .I(N__9368));
    LocalMux I__2149 (
            .O(N__9417),
            .I(N__9368));
    LocalMux I__2148 (
            .O(N__9414),
            .I(N__9365));
    InMux I__2147 (
            .O(N__9413),
            .I(N__9362));
    LocalMux I__2146 (
            .O(N__9410),
            .I(N__9355));
    LocalMux I__2145 (
            .O(N__9405),
            .I(N__9355));
    LocalMux I__2144 (
            .O(N__9400),
            .I(N__9355));
    LocalMux I__2143 (
            .O(N__9397),
            .I(N__9350));
    LocalMux I__2142 (
            .O(N__9392),
            .I(N__9350));
    LocalMux I__2141 (
            .O(N__9389),
            .I(N__9345));
    LocalMux I__2140 (
            .O(N__9386),
            .I(N__9345));
    InMux I__2139 (
            .O(N__9385),
            .I(N__9342));
    Span4Mux_v I__2138 (
            .O(N__9380),
            .I(N__9334));
    Span4Mux_v I__2137 (
            .O(N__9375),
            .I(N__9334));
    Span4Mux_v I__2136 (
            .O(N__9368),
            .I(N__9325));
    Span4Mux_v I__2135 (
            .O(N__9365),
            .I(N__9325));
    LocalMux I__2134 (
            .O(N__9362),
            .I(N__9325));
    Span4Mux_h I__2133 (
            .O(N__9355),
            .I(N__9325));
    Span4Mux_h I__2132 (
            .O(N__9350),
            .I(N__9322));
    Span4Mux_v I__2131 (
            .O(N__9345),
            .I(N__9317));
    LocalMux I__2130 (
            .O(N__9342),
            .I(N__9314));
    InMux I__2129 (
            .O(N__9341),
            .I(N__9311));
    InMux I__2128 (
            .O(N__9340),
            .I(N__9306));
    InMux I__2127 (
            .O(N__9339),
            .I(N__9306));
    Span4Mux_h I__2126 (
            .O(N__9334),
            .I(N__9303));
    Span4Mux_h I__2125 (
            .O(N__9325),
            .I(N__9300));
    Span4Mux_h I__2124 (
            .O(N__9322),
            .I(N__9297));
    InMux I__2123 (
            .O(N__9321),
            .I(N__9294));
    InMux I__2122 (
            .O(N__9320),
            .I(N__9291));
    Odrv4 I__2121 (
            .O(N__9317),
            .I(CPU_CYCLEm));
    Odrv12 I__2120 (
            .O(N__9314),
            .I(CPU_CYCLEm));
    LocalMux I__2119 (
            .O(N__9311),
            .I(CPU_CYCLEm));
    LocalMux I__2118 (
            .O(N__9306),
            .I(CPU_CYCLEm));
    Odrv4 I__2117 (
            .O(N__9303),
            .I(CPU_CYCLEm));
    Odrv4 I__2116 (
            .O(N__9300),
            .I(CPU_CYCLEm));
    Odrv4 I__2115 (
            .O(N__9297),
            .I(CPU_CYCLEm));
    LocalMux I__2114 (
            .O(N__9294),
            .I(CPU_CYCLEm));
    LocalMux I__2113 (
            .O(N__9291),
            .I(CPU_CYCLEm));
    IoInMux I__2112 (
            .O(N__9272),
            .I(N__9269));
    LocalMux I__2111 (
            .O(N__9269),
            .I(N__9266));
    Span4Mux_s3_h I__2110 (
            .O(N__9266),
            .I(N__9263));
    Span4Mux_v I__2109 (
            .O(N__9263),
            .I(N__9260));
    Span4Mux_v I__2108 (
            .O(N__9260),
            .I(N__9257));
    Sp12to4 I__2107 (
            .O(N__9257),
            .I(N__9254));
    Odrv12 I__2106 (
            .O(N__9254),
            .I(N_57_i));
    CascadeMux I__2105 (
            .O(N__9251),
            .I(N__9248));
    InMux I__2104 (
            .O(N__9248),
            .I(N__9245));
    LocalMux I__2103 (
            .O(N__9245),
            .I(\U712_BYTE_ENABLE.UUBE ));
    IoInMux I__2102 (
            .O(N__9242),
            .I(N__9239));
    LocalMux I__2101 (
            .O(N__9239),
            .I(N__9236));
    Span4Mux_s3_v I__2100 (
            .O(N__9236),
            .I(N__9233));
    Span4Mux_v I__2099 (
            .O(N__9233),
            .I(N__9230));
    Odrv4 I__2098 (
            .O(N__9230),
            .I(N_185));
    IoInMux I__2097 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__2096 (
            .O(N__9224),
            .I(N__9221));
    Span4Mux_s3_v I__2095 (
            .O(N__9221),
            .I(N__9218));
    Sp12to4 I__2094 (
            .O(N__9218),
            .I(N__9215));
    Span12Mux_h I__2093 (
            .O(N__9215),
            .I(N__9212));
    Odrv12 I__2092 (
            .O(N__9212),
            .I(N_44));
    IoInMux I__2091 (
            .O(N__9209),
            .I(N__9206));
    LocalMux I__2090 (
            .O(N__9206),
            .I(N__9203));
    IoSpan4Mux I__2089 (
            .O(N__9203),
            .I(N__9200));
    Span4Mux_s2_v I__2088 (
            .O(N__9200),
            .I(N__9197));
    Span4Mux_v I__2087 (
            .O(N__9197),
            .I(N__9194));
    Span4Mux_h I__2086 (
            .O(N__9194),
            .I(N__9191));
    Odrv4 I__2085 (
            .O(N__9191),
            .I(CASn_c));
    InMux I__2084 (
            .O(N__9188),
            .I(N__9185));
    LocalMux I__2083 (
            .O(N__9185),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__2082 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__2081 (
            .O(N__9179),
            .I(N__9176));
    IoSpan4Mux I__2080 (
            .O(N__9176),
            .I(N__9173));
    Span4Mux_s3_h I__2079 (
            .O(N__9173),
            .I(N__9170));
    Sp12to4 I__2078 (
            .O(N__9170),
            .I(N__9167));
    Span12Mux_h I__2077 (
            .O(N__9167),
            .I(N__9164));
    Odrv12 I__2076 (
            .O(N__9164),
            .I(CMA_c_4));
    InMux I__2075 (
            .O(N__9161),
            .I(N__9158));
    LocalMux I__2074 (
            .O(N__9158),
            .I(N__9155));
    Span4Mux_v I__2073 (
            .O(N__9155),
            .I(N__9152));
    Span4Mux_v I__2072 (
            .O(N__9152),
            .I(N__9149));
    Sp12to4 I__2071 (
            .O(N__9149),
            .I(N__9146));
    Span12Mux_h I__2070 (
            .O(N__9146),
            .I(N__9143));
    Odrv12 I__2069 (
            .O(N__9143),
            .I(A_c_17));
    IoInMux I__2068 (
            .O(N__9140),
            .I(N__9137));
    LocalMux I__2067 (
            .O(N__9137),
            .I(N__9134));
    Span12Mux_s2_h I__2066 (
            .O(N__9134),
            .I(N__9131));
    Span12Mux_h I__2065 (
            .O(N__9131),
            .I(N__9128));
    Odrv12 I__2064 (
            .O(N__9128),
            .I(CMA_c_8));
    InMux I__2063 (
            .O(N__9125),
            .I(N__9122));
    LocalMux I__2062 (
            .O(N__9122),
            .I(N__9119));
    Odrv12 I__2061 (
            .O(N__9119),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    CascadeMux I__2060 (
            .O(N__9116),
            .I(N__9108));
    CascadeMux I__2059 (
            .O(N__9115),
            .I(N__9105));
    CascadeMux I__2058 (
            .O(N__9114),
            .I(N__9099));
    CascadeMux I__2057 (
            .O(N__9113),
            .I(N__9096));
    InMux I__2056 (
            .O(N__9112),
            .I(N__9092));
    InMux I__2055 (
            .O(N__9111),
            .I(N__9089));
    InMux I__2054 (
            .O(N__9108),
            .I(N__9084));
    InMux I__2053 (
            .O(N__9105),
            .I(N__9084));
    InMux I__2052 (
            .O(N__9104),
            .I(N__9079));
    InMux I__2051 (
            .O(N__9103),
            .I(N__9079));
    CascadeMux I__2050 (
            .O(N__9102),
            .I(N__9075));
    InMux I__2049 (
            .O(N__9099),
            .I(N__9070));
    InMux I__2048 (
            .O(N__9096),
            .I(N__9066));
    CascadeMux I__2047 (
            .O(N__9095),
            .I(N__9063));
    LocalMux I__2046 (
            .O(N__9092),
            .I(N__9055));
    LocalMux I__2045 (
            .O(N__9089),
            .I(N__9050));
    LocalMux I__2044 (
            .O(N__9084),
            .I(N__9045));
    LocalMux I__2043 (
            .O(N__9079),
            .I(N__9045));
    InMux I__2042 (
            .O(N__9078),
            .I(N__9038));
    InMux I__2041 (
            .O(N__9075),
            .I(N__9038));
    InMux I__2040 (
            .O(N__9074),
            .I(N__9038));
    InMux I__2039 (
            .O(N__9073),
            .I(N__9035));
    LocalMux I__2038 (
            .O(N__9070),
            .I(N__9031));
    InMux I__2037 (
            .O(N__9069),
            .I(N__9028));
    LocalMux I__2036 (
            .O(N__9066),
            .I(N__9025));
    InMux I__2035 (
            .O(N__9063),
            .I(N__9020));
    InMux I__2034 (
            .O(N__9062),
            .I(N__9020));
    InMux I__2033 (
            .O(N__9061),
            .I(N__9015));
    InMux I__2032 (
            .O(N__9060),
            .I(N__9015));
    InMux I__2031 (
            .O(N__9059),
            .I(N__9010));
    InMux I__2030 (
            .O(N__9058),
            .I(N__9010));
    Span4Mux_v I__2029 (
            .O(N__9055),
            .I(N__9005));
    InMux I__2028 (
            .O(N__9054),
            .I(N__9002));
    InMux I__2027 (
            .O(N__9053),
            .I(N__8999));
    Span4Mux_h I__2026 (
            .O(N__9050),
            .I(N__8990));
    Span4Mux_v I__2025 (
            .O(N__9045),
            .I(N__8990));
    LocalMux I__2024 (
            .O(N__9038),
            .I(N__8990));
    LocalMux I__2023 (
            .O(N__9035),
            .I(N__8990));
    InMux I__2022 (
            .O(N__9034),
            .I(N__8987));
    Span4Mux_h I__2021 (
            .O(N__9031),
            .I(N__8984));
    LocalMux I__2020 (
            .O(N__9028),
            .I(N__8981));
    Sp12to4 I__2019 (
            .O(N__9025),
            .I(N__8972));
    LocalMux I__2018 (
            .O(N__9020),
            .I(N__8972));
    LocalMux I__2017 (
            .O(N__9015),
            .I(N__8972));
    LocalMux I__2016 (
            .O(N__9010),
            .I(N__8972));
    InMux I__2015 (
            .O(N__9009),
            .I(N__8967));
    InMux I__2014 (
            .O(N__9008),
            .I(N__8967));
    Span4Mux_h I__2013 (
            .O(N__9005),
            .I(N__8960));
    LocalMux I__2012 (
            .O(N__9002),
            .I(N__8960));
    LocalMux I__2011 (
            .O(N__8999),
            .I(N__8960));
    Span4Mux_h I__2010 (
            .O(N__8990),
            .I(N__8957));
    LocalMux I__2009 (
            .O(N__8987),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2008 (
            .O(N__8984),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2007 (
            .O(N__8981),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2006 (
            .O(N__8972),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2005 (
            .O(N__8967),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2004 (
            .O(N__8960),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2003 (
            .O(N__8957),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__2002 (
            .O(N__8942),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ));
    IoInMux I__2001 (
            .O(N__8939),
            .I(N__8936));
    LocalMux I__2000 (
            .O(N__8936),
            .I(N__8933));
    Span12Mux_s2_h I__1999 (
            .O(N__8933),
            .I(N__8930));
    Span12Mux_h I__1998 (
            .O(N__8930),
            .I(N__8927));
    Odrv12 I__1997 (
            .O(N__8927),
            .I(CMA_c_6));
    InMux I__1996 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1995 (
            .O(N__8921),
            .I(N__8918));
    Odrv12 I__1994 (
            .O(N__8918),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1993 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__1992 (
            .O(N__8912),
            .I(N__8909));
    Span12Mux_s2_h I__1991 (
            .O(N__8909),
            .I(N__8906));
    Span12Mux_h I__1990 (
            .O(N__8906),
            .I(N__8903));
    Odrv12 I__1989 (
            .O(N__8903),
            .I(CMA_c_7));
    InMux I__1988 (
            .O(N__8900),
            .I(N__8892));
    InMux I__1987 (
            .O(N__8899),
            .I(N__8889));
    InMux I__1986 (
            .O(N__8898),
            .I(N__8884));
    InMux I__1985 (
            .O(N__8897),
            .I(N__8884));
    InMux I__1984 (
            .O(N__8896),
            .I(N__8879));
    InMux I__1983 (
            .O(N__8895),
            .I(N__8879));
    LocalMux I__1982 (
            .O(N__8892),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__1981 (
            .O(N__8889),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__1980 (
            .O(N__8884),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__1979 (
            .O(N__8879),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    CascadeMux I__1978 (
            .O(N__8870),
            .I(N__8864));
    CascadeMux I__1977 (
            .O(N__8869),
            .I(N__8860));
    CascadeMux I__1976 (
            .O(N__8868),
            .I(N__8857));
    CascadeMux I__1975 (
            .O(N__8867),
            .I(N__8853));
    InMux I__1974 (
            .O(N__8864),
            .I(N__8850));
    InMux I__1973 (
            .O(N__8863),
            .I(N__8847));
    InMux I__1972 (
            .O(N__8860),
            .I(N__8844));
    InMux I__1971 (
            .O(N__8857),
            .I(N__8841));
    InMux I__1970 (
            .O(N__8856),
            .I(N__8838));
    InMux I__1969 (
            .O(N__8853),
            .I(N__8835));
    LocalMux I__1968 (
            .O(N__8850),
            .I(N__8832));
    LocalMux I__1967 (
            .O(N__8847),
            .I(N__8827));
    LocalMux I__1966 (
            .O(N__8844),
            .I(N__8827));
    LocalMux I__1965 (
            .O(N__8841),
            .I(N__8822));
    LocalMux I__1964 (
            .O(N__8838),
            .I(N__8815));
    LocalMux I__1963 (
            .O(N__8835),
            .I(N__8815));
    Span4Mux_h I__1962 (
            .O(N__8832),
            .I(N__8815));
    Span4Mux_h I__1961 (
            .O(N__8827),
            .I(N__8812));
    InMux I__1960 (
            .O(N__8826),
            .I(N__8809));
    InMux I__1959 (
            .O(N__8825),
            .I(N__8806));
    Odrv4 I__1958 (
            .O(N__8822),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1957 (
            .O(N__8815),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1956 (
            .O(N__8812),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1955 (
            .O(N__8809),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1954 (
            .O(N__8806),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__1953 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__1952 (
            .O(N__8792),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1951 (
            .O(N__8789),
            .I(N__8786));
    LocalMux I__1950 (
            .O(N__8786),
            .I(N__8783));
    Span4Mux_s3_v I__1949 (
            .O(N__8783),
            .I(N__8780));
    Span4Mux_v I__1948 (
            .O(N__8780),
            .I(N__8777));
    Span4Mux_v I__1947 (
            .O(N__8777),
            .I(N__8774));
    Odrv4 I__1946 (
            .O(N__8774),
            .I(CMA_c_0));
    InMux I__1945 (
            .O(N__8771),
            .I(N__8767));
    InMux I__1944 (
            .O(N__8770),
            .I(N__8764));
    LocalMux I__1943 (
            .O(N__8767),
            .I(N__8759));
    LocalMux I__1942 (
            .O(N__8764),
            .I(N__8756));
    InMux I__1941 (
            .O(N__8763),
            .I(N__8751));
    InMux I__1940 (
            .O(N__8762),
            .I(N__8751));
    Span4Mux_v I__1939 (
            .O(N__8759),
            .I(N__8746));
    Span4Mux_v I__1938 (
            .O(N__8756),
            .I(N__8746));
    LocalMux I__1937 (
            .O(N__8751),
            .I(N__8743));
    Odrv4 I__1936 (
            .O(N__8746),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv4 I__1935 (
            .O(N__8743),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1934 (
            .O(N__8738),
            .I(N__8735));
    LocalMux I__1933 (
            .O(N__8735),
            .I(N__8732));
    Span4Mux_h I__1932 (
            .O(N__8732),
            .I(N__8729));
    Sp12to4 I__1931 (
            .O(N__8729),
            .I(N__8726));
    Span12Mux_v I__1930 (
            .O(N__8726),
            .I(N__8723));
    Span12Mux_h I__1929 (
            .O(N__8723),
            .I(N__8720));
    Odrv12 I__1928 (
            .O(N__8720),
            .I(A_c_19));
    IoInMux I__1927 (
            .O(N__8717),
            .I(N__8714));
    LocalMux I__1926 (
            .O(N__8714),
            .I(N__8711));
    IoSpan4Mux I__1925 (
            .O(N__8711),
            .I(N__8708));
    IoSpan4Mux I__1924 (
            .O(N__8708),
            .I(N__8705));
    Sp12to4 I__1923 (
            .O(N__8705),
            .I(N__8702));
    Span12Mux_s7_h I__1922 (
            .O(N__8702),
            .I(N__8699));
    Odrv12 I__1921 (
            .O(N__8699),
            .I(CMA_c_9));
    InMux I__1920 (
            .O(N__8696),
            .I(N__8693));
    LocalMux I__1919 (
            .O(N__8693),
            .I(N__8662));
    ClkMux I__1918 (
            .O(N__8692),
            .I(N__8579));
    ClkMux I__1917 (
            .O(N__8691),
            .I(N__8579));
    ClkMux I__1916 (
            .O(N__8690),
            .I(N__8579));
    ClkMux I__1915 (
            .O(N__8689),
            .I(N__8579));
    ClkMux I__1914 (
            .O(N__8688),
            .I(N__8579));
    ClkMux I__1913 (
            .O(N__8687),
            .I(N__8579));
    ClkMux I__1912 (
            .O(N__8686),
            .I(N__8579));
    ClkMux I__1911 (
            .O(N__8685),
            .I(N__8579));
    ClkMux I__1910 (
            .O(N__8684),
            .I(N__8579));
    ClkMux I__1909 (
            .O(N__8683),
            .I(N__8579));
    ClkMux I__1908 (
            .O(N__8682),
            .I(N__8579));
    ClkMux I__1907 (
            .O(N__8681),
            .I(N__8579));
    ClkMux I__1906 (
            .O(N__8680),
            .I(N__8579));
    ClkMux I__1905 (
            .O(N__8679),
            .I(N__8579));
    ClkMux I__1904 (
            .O(N__8678),
            .I(N__8579));
    ClkMux I__1903 (
            .O(N__8677),
            .I(N__8579));
    ClkMux I__1902 (
            .O(N__8676),
            .I(N__8579));
    ClkMux I__1901 (
            .O(N__8675),
            .I(N__8579));
    ClkMux I__1900 (
            .O(N__8674),
            .I(N__8579));
    ClkMux I__1899 (
            .O(N__8673),
            .I(N__8579));
    ClkMux I__1898 (
            .O(N__8672),
            .I(N__8579));
    ClkMux I__1897 (
            .O(N__8671),
            .I(N__8579));
    ClkMux I__1896 (
            .O(N__8670),
            .I(N__8579));
    ClkMux I__1895 (
            .O(N__8669),
            .I(N__8579));
    ClkMux I__1894 (
            .O(N__8668),
            .I(N__8579));
    ClkMux I__1893 (
            .O(N__8667),
            .I(N__8579));
    ClkMux I__1892 (
            .O(N__8666),
            .I(N__8579));
    ClkMux I__1891 (
            .O(N__8665),
            .I(N__8579));
    Glb2LocalMux I__1890 (
            .O(N__8662),
            .I(N__8579));
    ClkMux I__1889 (
            .O(N__8661),
            .I(N__8579));
    ClkMux I__1888 (
            .O(N__8660),
            .I(N__8579));
    ClkMux I__1887 (
            .O(N__8659),
            .I(N__8579));
    ClkMux I__1886 (
            .O(N__8658),
            .I(N__8579));
    ClkMux I__1885 (
            .O(N__8657),
            .I(N__8579));
    ClkMux I__1884 (
            .O(N__8656),
            .I(N__8579));
    ClkMux I__1883 (
            .O(N__8655),
            .I(N__8579));
    ClkMux I__1882 (
            .O(N__8654),
            .I(N__8579));
    GlobalMux I__1881 (
            .O(N__8579),
            .I(CLK80_PLL));
    CEMux I__1880 (
            .O(N__8576),
            .I(N__8573));
    LocalMux I__1879 (
            .O(N__8573),
            .I(N__8567));
    CEMux I__1878 (
            .O(N__8572),
            .I(N__8564));
    CEMux I__1877 (
            .O(N__8571),
            .I(N__8560));
    CEMux I__1876 (
            .O(N__8570),
            .I(N__8557));
    Span4Mux_v I__1875 (
            .O(N__8567),
            .I(N__8554));
    LocalMux I__1874 (
            .O(N__8564),
            .I(N__8551));
    CEMux I__1873 (
            .O(N__8563),
            .I(N__8548));
    LocalMux I__1872 (
            .O(N__8560),
            .I(N__8543));
    LocalMux I__1871 (
            .O(N__8557),
            .I(N__8540));
    Span4Mux_h I__1870 (
            .O(N__8554),
            .I(N__8533));
    Span4Mux_h I__1869 (
            .O(N__8551),
            .I(N__8533));
    LocalMux I__1868 (
            .O(N__8548),
            .I(N__8533));
    CEMux I__1867 (
            .O(N__8547),
            .I(N__8530));
    CEMux I__1866 (
            .O(N__8546),
            .I(N__8527));
    Span4Mux_v I__1865 (
            .O(N__8543),
            .I(N__8522));
    Span4Mux_v I__1864 (
            .O(N__8540),
            .I(N__8522));
    Span4Mux_v I__1863 (
            .O(N__8533),
            .I(N__8517));
    LocalMux I__1862 (
            .O(N__8530),
            .I(N__8517));
    LocalMux I__1861 (
            .O(N__8527),
            .I(N__8514));
    Span4Mux_h I__1860 (
            .O(N__8522),
            .I(N__8511));
    Span4Mux_v I__1859 (
            .O(N__8517),
            .I(N__8508));
    Odrv4 I__1858 (
            .O(N__8514),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1857 (
            .O(N__8511),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1856 (
            .O(N__8508),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    CascadeMux I__1855 (
            .O(N__8501),
            .I(N__8498));
    InMux I__1854 (
            .O(N__8498),
            .I(N__8492));
    InMux I__1853 (
            .O(N__8497),
            .I(N__8492));
    LocalMux I__1852 (
            .O(N__8492),
            .I(N__8489));
    Span4Mux_v I__1851 (
            .O(N__8489),
            .I(N__8486));
    Odrv4 I__1850 (
            .O(N__8486),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1849 (
            .O(N__8483),
            .I(N__8475));
    InMux I__1848 (
            .O(N__8482),
            .I(N__8475));
    InMux I__1847 (
            .O(N__8481),
            .I(N__8472));
    InMux I__1846 (
            .O(N__8480),
            .I(N__8469));
    LocalMux I__1845 (
            .O(N__8475),
            .I(N__8462));
    LocalMux I__1844 (
            .O(N__8472),
            .I(N__8462));
    LocalMux I__1843 (
            .O(N__8469),
            .I(N__8462));
    Span4Mux_v I__1842 (
            .O(N__8462),
            .I(N__8459));
    Span4Mux_v I__1841 (
            .O(N__8459),
            .I(N__8456));
    Sp12to4 I__1840 (
            .O(N__8456),
            .I(N__8453));
    Span12Mux_h I__1839 (
            .O(N__8453),
            .I(N__8450));
    Odrv12 I__1838 (
            .O(N__8450),
            .I(DRA_c_3));
    CascadeMux I__1837 (
            .O(N__8447),
            .I(N__8444));
    InMux I__1836 (
            .O(N__8444),
            .I(N__8441));
    LocalMux I__1835 (
            .O(N__8441),
            .I(N__8438));
    Odrv4 I__1834 (
            .O(N__8438),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1833 (
            .O(N__8435),
            .I(N__8432));
    LocalMux I__1832 (
            .O(N__8432),
            .I(N__8429));
    Span4Mux_h I__1831 (
            .O(N__8429),
            .I(N__8426));
    Odrv4 I__1830 (
            .O(N__8426),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1829 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__1828 (
            .O(N__8420),
            .I(N__8417));
    Odrv4 I__1827 (
            .O(N__8417),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1826 (
            .O(N__8414),
            .I(N__8409));
    InMux I__1825 (
            .O(N__8413),
            .I(N__8406));
    InMux I__1824 (
            .O(N__8412),
            .I(N__8403));
    LocalMux I__1823 (
            .O(N__8409),
            .I(N__8399));
    LocalMux I__1822 (
            .O(N__8406),
            .I(N__8396));
    LocalMux I__1821 (
            .O(N__8403),
            .I(N__8393));
    InMux I__1820 (
            .O(N__8402),
            .I(N__8390));
    Span4Mux_v I__1819 (
            .O(N__8399),
            .I(N__8387));
    Span4Mux_h I__1818 (
            .O(N__8396),
            .I(N__8380));
    Span4Mux_v I__1817 (
            .O(N__8393),
            .I(N__8380));
    LocalMux I__1816 (
            .O(N__8390),
            .I(N__8380));
    Sp12to4 I__1815 (
            .O(N__8387),
            .I(N__8377));
    Sp12to4 I__1814 (
            .O(N__8380),
            .I(N__8374));
    Span12Mux_h I__1813 (
            .O(N__8377),
            .I(N__8371));
    Span12Mux_v I__1812 (
            .O(N__8374),
            .I(N__8368));
    Span12Mux_v I__1811 (
            .O(N__8371),
            .I(N__8365));
    Span12Mux_h I__1810 (
            .O(N__8368),
            .I(N__8362));
    Odrv12 I__1809 (
            .O(N__8365),
            .I(DRA_c_2));
    Odrv12 I__1808 (
            .O(N__8362),
            .I(DRA_c_2));
    InMux I__1807 (
            .O(N__8357),
            .I(N__8354));
    LocalMux I__1806 (
            .O(N__8354),
            .I(N__8351));
    Odrv4 I__1805 (
            .O(N__8351),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1804 (
            .O(N__8348),
            .I(N__8345));
    LocalMux I__1803 (
            .O(N__8345),
            .I(N__8342));
    Span4Mux_h I__1802 (
            .O(N__8342),
            .I(N__8338));
    InMux I__1801 (
            .O(N__8341),
            .I(N__8335));
    Odrv4 I__1800 (
            .O(N__8338),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0 ));
    LocalMux I__1799 (
            .O(N__8335),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0 ));
    IoInMux I__1798 (
            .O(N__8330),
            .I(N__8327));
    LocalMux I__1797 (
            .O(N__8327),
            .I(N__8324));
    Span4Mux_s3_h I__1796 (
            .O(N__8324),
            .I(N__8321));
    Sp12to4 I__1795 (
            .O(N__8321),
            .I(N__8318));
    Span12Mux_v I__1794 (
            .O(N__8318),
            .I(N__8315));
    Span12Mux_h I__1793 (
            .O(N__8315),
            .I(N__8312));
    Odrv12 I__1792 (
            .O(N__8312),
            .I(N_53_i));
    InMux I__1791 (
            .O(N__8309),
            .I(N__8306));
    LocalMux I__1790 (
            .O(N__8306),
            .I(\U712_BYTE_ENABLE.N_303 ));
    IoInMux I__1789 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__1788 (
            .O(N__8300),
            .I(N__8297));
    Span4Mux_s3_v I__1787 (
            .O(N__8297),
            .I(N__8294));
    Span4Mux_h I__1786 (
            .O(N__8294),
            .I(N__8291));
    Span4Mux_h I__1785 (
            .O(N__8291),
            .I(N__8288));
    Odrv4 I__1784 (
            .O(N__8288),
            .I(UMBE_0_o2_i));
    IoInMux I__1783 (
            .O(N__8285),
            .I(N__8282));
    LocalMux I__1782 (
            .O(N__8282),
            .I(N__8279));
    Span4Mux_s2_v I__1781 (
            .O(N__8279),
            .I(N__8276));
    Span4Mux_v I__1780 (
            .O(N__8276),
            .I(N__8273));
    Odrv4 I__1779 (
            .O(N__8273),
            .I(U712_BYTE_ENABLE_UUBE_i));
    InMux I__1778 (
            .O(N__8270),
            .I(N__8266));
    InMux I__1777 (
            .O(N__8269),
            .I(N__8263));
    LocalMux I__1776 (
            .O(N__8266),
            .I(N__8257));
    LocalMux I__1775 (
            .O(N__8263),
            .I(N__8254));
    InMux I__1774 (
            .O(N__8262),
            .I(N__8251));
    InMux I__1773 (
            .O(N__8261),
            .I(N__8248));
    InMux I__1772 (
            .O(N__8260),
            .I(N__8244));
    Span4Mux_v I__1771 (
            .O(N__8257),
            .I(N__8235));
    Span4Mux_h I__1770 (
            .O(N__8254),
            .I(N__8235));
    LocalMux I__1769 (
            .O(N__8251),
            .I(N__8235));
    LocalMux I__1768 (
            .O(N__8248),
            .I(N__8235));
    InMux I__1767 (
            .O(N__8247),
            .I(N__8232));
    LocalMux I__1766 (
            .O(N__8244),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1765 (
            .O(N__8235),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1764 (
            .O(N__8232),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__1763 (
            .O(N__8225),
            .I(N__8220));
    CascadeMux I__1762 (
            .O(N__8224),
            .I(N__8216));
    InMux I__1761 (
            .O(N__8223),
            .I(N__8213));
    InMux I__1760 (
            .O(N__8220),
            .I(N__8210));
    InMux I__1759 (
            .O(N__8219),
            .I(N__8205));
    InMux I__1758 (
            .O(N__8216),
            .I(N__8205));
    LocalMux I__1757 (
            .O(N__8213),
            .I(N__8201));
    LocalMux I__1756 (
            .O(N__8210),
            .I(N__8195));
    LocalMux I__1755 (
            .O(N__8205),
            .I(N__8195));
    InMux I__1754 (
            .O(N__8204),
            .I(N__8192));
    Span4Mux_h I__1753 (
            .O(N__8201),
            .I(N__8189));
    InMux I__1752 (
            .O(N__8200),
            .I(N__8186));
    Span4Mux_h I__1751 (
            .O(N__8195),
            .I(N__8181));
    LocalMux I__1750 (
            .O(N__8192),
            .I(N__8181));
    Odrv4 I__1749 (
            .O(N__8189),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1748 (
            .O(N__8186),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1747 (
            .O(N__8181),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1746 (
            .O(N__8174),
            .I(N__8170));
    InMux I__1745 (
            .O(N__8173),
            .I(N__8167));
    LocalMux I__1744 (
            .O(N__8170),
            .I(N__8162));
    LocalMux I__1743 (
            .O(N__8167),
            .I(N__8159));
    InMux I__1742 (
            .O(N__8166),
            .I(N__8156));
    CascadeMux I__1741 (
            .O(N__8165),
            .I(N__8153));
    Span4Mux_v I__1740 (
            .O(N__8162),
            .I(N__8146));
    Span4Mux_h I__1739 (
            .O(N__8159),
            .I(N__8146));
    LocalMux I__1738 (
            .O(N__8156),
            .I(N__8146));
    InMux I__1737 (
            .O(N__8153),
            .I(N__8143));
    Odrv4 I__1736 (
            .O(N__8146),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1735 (
            .O(N__8143),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1734 (
            .O(N__8138),
            .I(N__8135));
    LocalMux I__1733 (
            .O(N__8135),
            .I(N__8132));
    Span4Mux_s3_v I__1732 (
            .O(N__8132),
            .I(N__8129));
    Sp12to4 I__1731 (
            .O(N__8129),
            .I(N__8126));
    Span12Mux_h I__1730 (
            .O(N__8126),
            .I(N__8123));
    Odrv12 I__1729 (
            .O(N__8123),
            .I(CMA_c_10));
    InMux I__1728 (
            .O(N__8120),
            .I(N__8117));
    LocalMux I__1727 (
            .O(N__8117),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1726 (
            .O(N__8114),
            .I(N__8111));
    LocalMux I__1725 (
            .O(N__8111),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1724 (
            .O(N__8108),
            .I(N__8105));
    LocalMux I__1723 (
            .O(N__8105),
            .I(N__8102));
    Odrv4 I__1722 (
            .O(N__8102),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1721 (
            .O(N__8099),
            .I(N__8096));
    LocalMux I__1720 (
            .O(N__8096),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1719 (
            .O(N__8093),
            .I(N__8090));
    LocalMux I__1718 (
            .O(N__8090),
            .I(N__8087));
    Span12Mux_s11_v I__1717 (
            .O(N__8087),
            .I(N__8084));
    Odrv12 I__1716 (
            .O(N__8084),
            .I(CMA_c_2));
    IoInMux I__1715 (
            .O(N__8081),
            .I(N__8078));
    LocalMux I__1714 (
            .O(N__8078),
            .I(N__8075));
    Span4Mux_s3_h I__1713 (
            .O(N__8075),
            .I(N__8072));
    Sp12to4 I__1712 (
            .O(N__8072),
            .I(N__8069));
    Span12Mux_s6_v I__1711 (
            .O(N__8069),
            .I(N__8066));
    Span12Mux_h I__1710 (
            .O(N__8066),
            .I(N__8063));
    Odrv12 I__1709 (
            .O(N__8063),
            .I(CMA_c_3));
    InMux I__1708 (
            .O(N__8060),
            .I(N__8057));
    LocalMux I__1707 (
            .O(N__8057),
            .I(N__8054));
    Odrv4 I__1706 (
            .O(N__8054),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1705 (
            .O(N__8051),
            .I(N__8048));
    LocalMux I__1704 (
            .O(N__8048),
            .I(N__8045));
    Span4Mux_h I__1703 (
            .O(N__8045),
            .I(N__8042));
    Odrv4 I__1702 (
            .O(N__8042),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1701 (
            .O(N__8039),
            .I(N__8036));
    LocalMux I__1700 (
            .O(N__8036),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1699 (
            .O(N__8033),
            .I(N__8027));
    InMux I__1698 (
            .O(N__8032),
            .I(N__8027));
    LocalMux I__1697 (
            .O(N__8027),
            .I(N__8024));
    Span4Mux_h I__1696 (
            .O(N__8024),
            .I(N__8021));
    Odrv4 I__1695 (
            .O(N__8021),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1694 (
            .O(N__8018),
            .I(N__8015));
    LocalMux I__1693 (
            .O(N__8015),
            .I(N__8012));
    Span4Mux_v I__1692 (
            .O(N__8012),
            .I(N__8009));
    Odrv4 I__1691 (
            .O(N__8009),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1690 (
            .O(N__8006),
            .I(N__8003));
    LocalMux I__1689 (
            .O(N__8003),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1688 (
            .O(N__8000),
            .I(N__7996));
    InMux I__1687 (
            .O(N__7999),
            .I(N__7993));
    LocalMux I__1686 (
            .O(N__7996),
            .I(N__7990));
    LocalMux I__1685 (
            .O(N__7993),
            .I(N__7987));
    Odrv12 I__1684 (
            .O(N__7990),
            .I(DBRn_c_i));
    Odrv12 I__1683 (
            .O(N__7987),
            .I(DBRn_c_i));
    InMux I__1682 (
            .O(N__7982),
            .I(N__7979));
    LocalMux I__1681 (
            .O(N__7979),
            .I(N__7976));
    Span4Mux_h I__1680 (
            .O(N__7976),
            .I(N__7972));
    InMux I__1679 (
            .O(N__7975),
            .I(N__7969));
    Span4Mux_h I__1678 (
            .O(N__7972),
            .I(N__7966));
    LocalMux I__1677 (
            .O(N__7969),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__1676 (
            .O(N__7966),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__1675 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1674 (
            .O(N__7958),
            .I(N__7954));
    InMux I__1673 (
            .O(N__7957),
            .I(N__7951));
    Odrv4 I__1672 (
            .O(N__7954),
            .I(\U712_BYTE_ENABLE.N_370 ));
    LocalMux I__1671 (
            .O(N__7951),
            .I(\U712_BYTE_ENABLE.N_370 ));
    CascadeMux I__1670 (
            .O(N__7946),
            .I(\U712_BYTE_ENABLE.N_369_cascade_ ));
    IoInMux I__1669 (
            .O(N__7943),
            .I(N__7940));
    LocalMux I__1668 (
            .O(N__7940),
            .I(N__7937));
    Span4Mux_s0_h I__1667 (
            .O(N__7937),
            .I(N__7934));
    Span4Mux_h I__1666 (
            .O(N__7934),
            .I(N__7931));
    Sp12to4 I__1665 (
            .O(N__7931),
            .I(N__7928));
    Span12Mux_s11_v I__1664 (
            .O(N__7928),
            .I(N__7925));
    Span12Mux_h I__1663 (
            .O(N__7925),
            .I(N__7922));
    Odrv12 I__1662 (
            .O(N__7922),
            .I(N_55_i));
    IoInMux I__1661 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__1660 (
            .O(N__7916),
            .I(N__7913));
    Span4Mux_s3_h I__1659 (
            .O(N__7913),
            .I(N__7910));
    Sp12to4 I__1658 (
            .O(N__7910),
            .I(N__7907));
    Span12Mux_s6_v I__1657 (
            .O(N__7907),
            .I(N__7904));
    Odrv12 I__1656 (
            .O(N__7904),
            .I(WEn_c));
    IoInMux I__1655 (
            .O(N__7901),
            .I(N__7898));
    LocalMux I__1654 (
            .O(N__7898),
            .I(N__7895));
    Span4Mux_s3_v I__1653 (
            .O(N__7895),
            .I(N__7892));
    Span4Mux_v I__1652 (
            .O(N__7892),
            .I(N__7889));
    Span4Mux_h I__1651 (
            .O(N__7889),
            .I(N__7886));
    Odrv4 I__1650 (
            .O(N__7886),
            .I(CRCSn_c));
    IoInMux I__1649 (
            .O(N__7883),
            .I(N__7880));
    LocalMux I__1648 (
            .O(N__7880),
            .I(N__7877));
    Span4Mux_s2_v I__1647 (
            .O(N__7877),
            .I(N__7874));
    Sp12to4 I__1646 (
            .O(N__7874),
            .I(N__7871));
    Span12Mux_h I__1645 (
            .O(N__7871),
            .I(N__7868));
    Odrv12 I__1644 (
            .O(N__7868),
            .I(RASn_c));
    CascadeMux I__1643 (
            .O(N__7865),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ));
    InMux I__1642 (
            .O(N__7862),
            .I(N__7859));
    LocalMux I__1641 (
            .O(N__7859),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1640 (
            .O(N__7856),
            .I(N__7853));
    LocalMux I__1639 (
            .O(N__7853),
            .I(N__7850));
    Span4Mux_h I__1638 (
            .O(N__7850),
            .I(N__7847));
    Odrv4 I__1637 (
            .O(N__7847),
            .I(\U712_CHIP_RAM.N_392 ));
    InMux I__1636 (
            .O(N__7844),
            .I(N__7841));
    LocalMux I__1635 (
            .O(N__7841),
            .I(N__7838));
    Span12Mux_h I__1634 (
            .O(N__7838),
            .I(N__7835));
    Odrv12 I__1633 (
            .O(N__7835),
            .I(A_c_13));
    InMux I__1632 (
            .O(N__7832),
            .I(N__7829));
    LocalMux I__1631 (
            .O(N__7829),
            .I(N__7826));
    Span4Mux_v I__1630 (
            .O(N__7826),
            .I(N__7823));
    Span4Mux_v I__1629 (
            .O(N__7823),
            .I(N__7820));
    Sp12to4 I__1628 (
            .O(N__7820),
            .I(N__7817));
    Span12Mux_h I__1627 (
            .O(N__7817),
            .I(N__7814));
    Odrv12 I__1626 (
            .O(N__7814),
            .I(A_c_6));
    InMux I__1625 (
            .O(N__7811),
            .I(N__7805));
    InMux I__1624 (
            .O(N__7810),
            .I(N__7805));
    LocalMux I__1623 (
            .O(N__7805),
            .I(N__7802));
    Span4Mux_v I__1622 (
            .O(N__7802),
            .I(N__7799));
    Span4Mux_v I__1621 (
            .O(N__7799),
            .I(N__7796));
    Sp12to4 I__1620 (
            .O(N__7796),
            .I(N__7793));
    Span12Mux_h I__1619 (
            .O(N__7793),
            .I(N__7790));
    Odrv12 I__1618 (
            .O(N__7790),
            .I(A_c_14));
    InMux I__1617 (
            .O(N__7787),
            .I(N__7784));
    LocalMux I__1616 (
            .O(N__7784),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1615 (
            .O(N__7781),
            .I(N__7778));
    LocalMux I__1614 (
            .O(N__7778),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1613 (
            .O(N__7775),
            .I(N__7772));
    LocalMux I__1612 (
            .O(N__7772),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1611 (
            .O(N__7769),
            .I(N__7766));
    LocalMux I__1610 (
            .O(N__7766),
            .I(N__7763));
    IoSpan4Mux I__1609 (
            .O(N__7763),
            .I(N__7760));
    Span4Mux_s2_h I__1608 (
            .O(N__7760),
            .I(N__7757));
    Sp12to4 I__1607 (
            .O(N__7757),
            .I(N__7754));
    Span12Mux_h I__1606 (
            .O(N__7754),
            .I(N__7751));
    Odrv12 I__1605 (
            .O(N__7751),
            .I(CMA_c_5));
    InMux I__1604 (
            .O(N__7748),
            .I(N__7745));
    LocalMux I__1603 (
            .O(N__7745),
            .I(N__7742));
    Span12Mux_v I__1602 (
            .O(N__7742),
            .I(N__7739));
    Span12Mux_h I__1601 (
            .O(N__7739),
            .I(N__7736));
    Odrv12 I__1600 (
            .O(N__7736),
            .I(A_c_11));
    InMux I__1599 (
            .O(N__7733),
            .I(N__7730));
    LocalMux I__1598 (
            .O(N__7730),
            .I(N__7727));
    Span4Mux_v I__1597 (
            .O(N__7727),
            .I(N__7724));
    Span4Mux_v I__1596 (
            .O(N__7724),
            .I(N__7721));
    Sp12to4 I__1595 (
            .O(N__7721),
            .I(N__7718));
    Span12Mux_h I__1594 (
            .O(N__7718),
            .I(N__7715));
    Odrv12 I__1593 (
            .O(N__7715),
            .I(A_c_4));
    CascadeMux I__1592 (
            .O(N__7712),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__1591 (
            .O(N__7709),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1590 (
            .O(N__7706),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__1589 (
            .O(N__7703),
            .I(N__7699));
    InMux I__1588 (
            .O(N__7702),
            .I(N__7696));
    LocalMux I__1587 (
            .O(N__7699),
            .I(N__7684));
    LocalMux I__1586 (
            .O(N__7696),
            .I(N__7681));
    ClkMux I__1585 (
            .O(N__7695),
            .I(N__7658));
    ClkMux I__1584 (
            .O(N__7694),
            .I(N__7658));
    ClkMux I__1583 (
            .O(N__7693),
            .I(N__7658));
    ClkMux I__1582 (
            .O(N__7692),
            .I(N__7658));
    ClkMux I__1581 (
            .O(N__7691),
            .I(N__7658));
    ClkMux I__1580 (
            .O(N__7690),
            .I(N__7658));
    ClkMux I__1579 (
            .O(N__7689),
            .I(N__7658));
    ClkMux I__1578 (
            .O(N__7688),
            .I(N__7658));
    ClkMux I__1577 (
            .O(N__7687),
            .I(N__7658));
    Glb2LocalMux I__1576 (
            .O(N__7684),
            .I(N__7658));
    Glb2LocalMux I__1575 (
            .O(N__7681),
            .I(N__7658));
    GlobalMux I__1574 (
            .O(N__7658),
            .I(N__7655));
    gio2CtrlBuf I__1573 (
            .O(N__7655),
            .I(C1_c_g));
    SRMux I__1572 (
            .O(N__7652),
            .I(N__7649));
    LocalMux I__1571 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_v I__1570 (
            .O(N__7646),
            .I(N__7643));
    Odrv4 I__1569 (
            .O(N__7643),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1568 (
            .O(N__7640),
            .I(N__7636));
    InMux I__1567 (
            .O(N__7639),
            .I(N__7633));
    LocalMux I__1566 (
            .O(N__7636),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1565 (
            .O(N__7633),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1564 (
            .O(N__7628),
            .I(N__7624));
    InMux I__1563 (
            .O(N__7627),
            .I(N__7621));
    LocalMux I__1562 (
            .O(N__7624),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1561 (
            .O(N__7621),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1560 (
            .O(N__7616),
            .I(N__7612));
    InMux I__1559 (
            .O(N__7615),
            .I(N__7609));
    LocalMux I__1558 (
            .O(N__7612),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1557 (
            .O(N__7609),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1556 (
            .O(N__7604),
            .I(N__7601));
    LocalMux I__1555 (
            .O(N__7601),
            .I(N__7598));
    Odrv4 I__1554 (
            .O(N__7598),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__1553 (
            .O(N__7595),
            .I(N__7591));
    InMux I__1552 (
            .O(N__7594),
            .I(N__7588));
    LocalMux I__1551 (
            .O(N__7591),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1550 (
            .O(N__7588),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1549 (
            .O(N__7583),
            .I(N__7579));
    InMux I__1548 (
            .O(N__7582),
            .I(N__7576));
    LocalMux I__1547 (
            .O(N__7579),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__1546 (
            .O(N__7576),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    CascadeMux I__1545 (
            .O(N__7571),
            .I(N__7567));
    InMux I__1544 (
            .O(N__7570),
            .I(N__7564));
    InMux I__1543 (
            .O(N__7567),
            .I(N__7561));
    LocalMux I__1542 (
            .O(N__7564),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1541 (
            .O(N__7561),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1540 (
            .O(N__7556),
            .I(N__7552));
    InMux I__1539 (
            .O(N__7555),
            .I(N__7549));
    LocalMux I__1538 (
            .O(N__7552),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__1537 (
            .O(N__7549),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__1536 (
            .O(N__7544),
            .I(N__7541));
    LocalMux I__1535 (
            .O(N__7541),
            .I(N__7538));
    Odrv4 I__1534 (
            .O(N__7538),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    CascadeMux I__1533 (
            .O(N__7535),
            .I(N__7523));
    CascadeMux I__1532 (
            .O(N__7534),
            .I(N__7512));
    InMux I__1531 (
            .O(N__7533),
            .I(N__7509));
    InMux I__1530 (
            .O(N__7532),
            .I(N__7506));
    InMux I__1529 (
            .O(N__7531),
            .I(N__7499));
    InMux I__1528 (
            .O(N__7530),
            .I(N__7499));
    InMux I__1527 (
            .O(N__7529),
            .I(N__7499));
    InMux I__1526 (
            .O(N__7528),
            .I(N__7496));
    InMux I__1525 (
            .O(N__7527),
            .I(N__7492));
    InMux I__1524 (
            .O(N__7526),
            .I(N__7485));
    InMux I__1523 (
            .O(N__7523),
            .I(N__7485));
    InMux I__1522 (
            .O(N__7522),
            .I(N__7485));
    InMux I__1521 (
            .O(N__7521),
            .I(N__7482));
    CascadeMux I__1520 (
            .O(N__7520),
            .I(N__7478));
    InMux I__1519 (
            .O(N__7519),
            .I(N__7471));
    InMux I__1518 (
            .O(N__7518),
            .I(N__7471));
    InMux I__1517 (
            .O(N__7517),
            .I(N__7468));
    InMux I__1516 (
            .O(N__7516),
            .I(N__7463));
    InMux I__1515 (
            .O(N__7515),
            .I(N__7463));
    InMux I__1514 (
            .O(N__7512),
            .I(N__7460));
    LocalMux I__1513 (
            .O(N__7509),
            .I(N__7457));
    LocalMux I__1512 (
            .O(N__7506),
            .I(N__7450));
    LocalMux I__1511 (
            .O(N__7499),
            .I(N__7450));
    LocalMux I__1510 (
            .O(N__7496),
            .I(N__7450));
    InMux I__1509 (
            .O(N__7495),
            .I(N__7447));
    LocalMux I__1508 (
            .O(N__7492),
            .I(N__7442));
    LocalMux I__1507 (
            .O(N__7485),
            .I(N__7437));
    LocalMux I__1506 (
            .O(N__7482),
            .I(N__7437));
    InMux I__1505 (
            .O(N__7481),
            .I(N__7432));
    InMux I__1504 (
            .O(N__7478),
            .I(N__7432));
    InMux I__1503 (
            .O(N__7477),
            .I(N__7429));
    InMux I__1502 (
            .O(N__7476),
            .I(N__7426));
    LocalMux I__1501 (
            .O(N__7471),
            .I(N__7421));
    LocalMux I__1500 (
            .O(N__7468),
            .I(N__7421));
    LocalMux I__1499 (
            .O(N__7463),
            .I(N__7416));
    LocalMux I__1498 (
            .O(N__7460),
            .I(N__7416));
    Span4Mux_v I__1497 (
            .O(N__7457),
            .I(N__7409));
    Span4Mux_v I__1496 (
            .O(N__7450),
            .I(N__7409));
    LocalMux I__1495 (
            .O(N__7447),
            .I(N__7409));
    InMux I__1494 (
            .O(N__7446),
            .I(N__7404));
    InMux I__1493 (
            .O(N__7445),
            .I(N__7404));
    Span4Mux_v I__1492 (
            .O(N__7442),
            .I(N__7393));
    Span4Mux_v I__1491 (
            .O(N__7437),
            .I(N__7393));
    LocalMux I__1490 (
            .O(N__7432),
            .I(N__7393));
    LocalMux I__1489 (
            .O(N__7429),
            .I(N__7393));
    LocalMux I__1488 (
            .O(N__7426),
            .I(N__7393));
    Span4Mux_v I__1487 (
            .O(N__7421),
            .I(N__7384));
    Span4Mux_h I__1486 (
            .O(N__7416),
            .I(N__7384));
    Span4Mux_h I__1485 (
            .O(N__7409),
            .I(N__7384));
    LocalMux I__1484 (
            .O(N__7404),
            .I(N__7384));
    Span4Mux_v I__1483 (
            .O(N__7393),
            .I(N__7378));
    Span4Mux_v I__1482 (
            .O(N__7384),
            .I(N__7375));
    InMux I__1481 (
            .O(N__7383),
            .I(N__7372));
    InMux I__1480 (
            .O(N__7382),
            .I(N__7369));
    InMux I__1479 (
            .O(N__7381),
            .I(N__7366));
    Sp12to4 I__1478 (
            .O(N__7378),
            .I(N__7355));
    Sp12to4 I__1477 (
            .O(N__7375),
            .I(N__7355));
    LocalMux I__1476 (
            .O(N__7372),
            .I(N__7355));
    LocalMux I__1475 (
            .O(N__7369),
            .I(N__7355));
    LocalMux I__1474 (
            .O(N__7366),
            .I(N__7355));
    Span12Mux_h I__1473 (
            .O(N__7355),
            .I(N__7352));
    Odrv12 I__1472 (
            .O(N__7352),
            .I(RESETn_c));
    IoInMux I__1471 (
            .O(N__7349),
            .I(N__7346));
    LocalMux I__1470 (
            .O(N__7346),
            .I(N__7343));
    IoSpan4Mux I__1469 (
            .O(N__7343),
            .I(N__7340));
    Span4Mux_s3_v I__1468 (
            .O(N__7340),
            .I(N__7336));
    InMux I__1467 (
            .O(N__7339),
            .I(N__7333));
    Span4Mux_v I__1466 (
            .O(N__7336),
            .I(N__7330));
    LocalMux I__1465 (
            .O(N__7333),
            .I(N__7327));
    Span4Mux_v I__1464 (
            .O(N__7330),
            .I(N__7324));
    Span4Mux_h I__1463 (
            .O(N__7327),
            .I(N__7321));
    Span4Mux_v I__1462 (
            .O(N__7324),
            .I(N__7316));
    Span4Mux_v I__1461 (
            .O(N__7321),
            .I(N__7316));
    Odrv4 I__1460 (
            .O(N__7316),
            .I(RESETn_c_i));
    InMux I__1459 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__1458 (
            .O(N__7310),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__1457 (
            .O(N__7307),
            .I(N__7304));
    LocalMux I__1456 (
            .O(N__7304),
            .I(N__7301));
    Odrv12 I__1455 (
            .O(N__7301),
            .I(CMA_c_1));
    InMux I__1454 (
            .O(N__7298),
            .I(N__7295));
    LocalMux I__1453 (
            .O(N__7295),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1452 (
            .O(N__7292),
            .I(N__7289));
    LocalMux I__1451 (
            .O(N__7289),
            .I(N__7286));
    Span4Mux_v I__1450 (
            .O(N__7286),
            .I(N__7283));
    Span4Mux_v I__1449 (
            .O(N__7283),
            .I(N__7280));
    Sp12to4 I__1448 (
            .O(N__7280),
            .I(N__7277));
    Span12Mux_h I__1447 (
            .O(N__7277),
            .I(N__7274));
    Odrv12 I__1446 (
            .O(N__7274),
            .I(A_c_16));
    InMux I__1445 (
            .O(N__7271),
            .I(N__7268));
    LocalMux I__1444 (
            .O(N__7268),
            .I(N__7265));
    Span4Mux_v I__1443 (
            .O(N__7265),
            .I(N__7262));
    Span4Mux_v I__1442 (
            .O(N__7262),
            .I(N__7259));
    Sp12to4 I__1441 (
            .O(N__7259),
            .I(N__7256));
    Span12Mux_h I__1440 (
            .O(N__7256),
            .I(N__7253));
    Odrv12 I__1439 (
            .O(N__7253),
            .I(A_c_18));
    CascadeMux I__1438 (
            .O(N__7250),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ));
    InMux I__1437 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__1436 (
            .O(N__7244),
            .I(\U712_CHIP_RAM.CLK_EN_5_0_a2_0 ));
    CascadeMux I__1435 (
            .O(N__7241),
            .I(N__7238));
    InMux I__1434 (
            .O(N__7238),
            .I(N__7235));
    LocalMux I__1433 (
            .O(N__7235),
            .I(\U712_CHIP_RAM.N_112 ));
    IoInMux I__1432 (
            .O(N__7232),
            .I(N__7229));
    LocalMux I__1431 (
            .O(N__7229),
            .I(N__7226));
    IoSpan4Mux I__1430 (
            .O(N__7226),
            .I(N__7223));
    IoSpan4Mux I__1429 (
            .O(N__7223),
            .I(N__7220));
    Span4Mux_s2_h I__1428 (
            .O(N__7220),
            .I(N__7217));
    Sp12to4 I__1427 (
            .O(N__7217),
            .I(N__7214));
    Span12Mux_s9_h I__1426 (
            .O(N__7214),
            .I(N__7210));
    InMux I__1425 (
            .O(N__7213),
            .I(N__7207));
    Odrv12 I__1424 (
            .O(N__7210),
            .I(CLK_EN_c));
    LocalMux I__1423 (
            .O(N__7207),
            .I(CLK_EN_c));
    InMux I__1422 (
            .O(N__7202),
            .I(bfn_11_7_0_));
    InMux I__1421 (
            .O(N__7199),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1420 (
            .O(N__7196),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1419 (
            .O(N__7193),
            .I(N__7190));
    LocalMux I__1418 (
            .O(N__7190),
            .I(N__7186));
    InMux I__1417 (
            .O(N__7189),
            .I(N__7183));
    Span4Mux_h I__1416 (
            .O(N__7186),
            .I(N__7180));
    LocalMux I__1415 (
            .O(N__7183),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__1414 (
            .O(N__7180),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1413 (
            .O(N__7175),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__1412 (
            .O(N__7172),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1411 (
            .O(N__7169),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    CascadeMux I__1410 (
            .O(N__7166),
            .I(N__7161));
    CascadeMux I__1409 (
            .O(N__7165),
            .I(N__7156));
    InMux I__1408 (
            .O(N__7164),
            .I(N__7148));
    InMux I__1407 (
            .O(N__7161),
            .I(N__7148));
    InMux I__1406 (
            .O(N__7160),
            .I(N__7148));
    InMux I__1405 (
            .O(N__7159),
            .I(N__7141));
    InMux I__1404 (
            .O(N__7156),
            .I(N__7141));
    InMux I__1403 (
            .O(N__7155),
            .I(N__7141));
    LocalMux I__1402 (
            .O(N__7148),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1401 (
            .O(N__7141),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__1400 (
            .O(N__7136),
            .I(N__7133));
    LocalMux I__1399 (
            .O(N__7133),
            .I(\U712_REG_SM.m17_i_0_o2_1 ));
    CascadeMux I__1398 (
            .O(N__7130),
            .I(N__7127));
    InMux I__1397 (
            .O(N__7127),
            .I(N__7124));
    LocalMux I__1396 (
            .O(N__7124),
            .I(\U712_REG_SM.N_435 ));
    CascadeMux I__1395 (
            .O(N__7121),
            .I(\U712_REG_SM.N_435_cascade_ ));
    InMux I__1394 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__1393 (
            .O(N__7115),
            .I(\U712_REG_SM.N_363 ));
    IoInMux I__1392 (
            .O(N__7112),
            .I(N__7108));
    IoInMux I__1391 (
            .O(N__7111),
            .I(N__7105));
    LocalMux I__1390 (
            .O(N__7108),
            .I(N__7102));
    LocalMux I__1389 (
            .O(N__7105),
            .I(N__7099));
    Span4Mux_s0_v I__1388 (
            .O(N__7102),
            .I(N__7096));
    Span4Mux_s0_v I__1387 (
            .O(N__7099),
            .I(N__7093));
    Span4Mux_v I__1386 (
            .O(N__7096),
            .I(N__7090));
    Span4Mux_v I__1385 (
            .O(N__7093),
            .I(N__7087));
    Sp12to4 I__1384 (
            .O(N__7090),
            .I(N__7084));
    Sp12to4 I__1383 (
            .O(N__7087),
            .I(N__7081));
    Span12Mux_s10_h I__1382 (
            .O(N__7084),
            .I(N__7078));
    Span12Mux_s9_h I__1381 (
            .O(N__7081),
            .I(N__7075));
    Span12Mux_v I__1380 (
            .O(N__7078),
            .I(N__7069));
    Span12Mux_v I__1379 (
            .O(N__7075),
            .I(N__7069));
    InMux I__1378 (
            .O(N__7074),
            .I(N__7066));
    Odrv12 I__1377 (
            .O(N__7069),
            .I(ASn_c));
    LocalMux I__1376 (
            .O(N__7066),
            .I(ASn_c));
    InMux I__1375 (
            .O(N__7061),
            .I(N__7055));
    InMux I__1374 (
            .O(N__7060),
            .I(N__7055));
    LocalMux I__1373 (
            .O(N__7055),
            .I(\U712_REG_SM.ASn_0_sqmuxa ));
    CascadeMux I__1372 (
            .O(N__7052),
            .I(N__7048));
    CascadeMux I__1371 (
            .O(N__7051),
            .I(N__7045));
    InMux I__1370 (
            .O(N__7048),
            .I(N__7031));
    InMux I__1369 (
            .O(N__7045),
            .I(N__7031));
    InMux I__1368 (
            .O(N__7044),
            .I(N__7022));
    InMux I__1367 (
            .O(N__7043),
            .I(N__7022));
    InMux I__1366 (
            .O(N__7042),
            .I(N__7022));
    InMux I__1365 (
            .O(N__7041),
            .I(N__7022));
    InMux I__1364 (
            .O(N__7040),
            .I(N__7013));
    InMux I__1363 (
            .O(N__7039),
            .I(N__7013));
    InMux I__1362 (
            .O(N__7038),
            .I(N__7013));
    InMux I__1361 (
            .O(N__7037),
            .I(N__7013));
    InMux I__1360 (
            .O(N__7036),
            .I(N__7010));
    LocalMux I__1359 (
            .O(N__7031),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1358 (
            .O(N__7022),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1357 (
            .O(N__7013),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1356 (
            .O(N__7010),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__1355 (
            .O(N__7001),
            .I(N__6993));
    InMux I__1354 (
            .O(N__7000),
            .I(N__6993));
    InMux I__1353 (
            .O(N__6999),
            .I(N__6990));
    InMux I__1352 (
            .O(N__6998),
            .I(N__6987));
    LocalMux I__1351 (
            .O(N__6993),
            .I(\U712_REG_SM.m17_i_0_o2 ));
    LocalMux I__1350 (
            .O(N__6990),
            .I(\U712_REG_SM.m17_i_0_o2 ));
    LocalMux I__1349 (
            .O(N__6987),
            .I(\U712_REG_SM.m17_i_0_o2 ));
    InMux I__1348 (
            .O(N__6980),
            .I(N__6973));
    InMux I__1347 (
            .O(N__6979),
            .I(N__6968));
    InMux I__1346 (
            .O(N__6978),
            .I(N__6968));
    InMux I__1345 (
            .O(N__6977),
            .I(N__6963));
    InMux I__1344 (
            .O(N__6976),
            .I(N__6963));
    LocalMux I__1343 (
            .O(N__6973),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1342 (
            .O(N__6968),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1341 (
            .O(N__6963),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__1340 (
            .O(N__6956),
            .I(N__6953));
    InMux I__1339 (
            .O(N__6953),
            .I(N__6945));
    InMux I__1338 (
            .O(N__6952),
            .I(N__6945));
    InMux I__1337 (
            .O(N__6951),
            .I(N__6940));
    InMux I__1336 (
            .O(N__6950),
            .I(N__6940));
    LocalMux I__1335 (
            .O(N__6945),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1334 (
            .O(N__6940),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__1333 (
            .O(N__6935),
            .I(N__6931));
    InMux I__1332 (
            .O(N__6934),
            .I(N__6927));
    LocalMux I__1331 (
            .O(N__6931),
            .I(N__6924));
    InMux I__1330 (
            .O(N__6930),
            .I(N__6921));
    LocalMux I__1329 (
            .O(N__6927),
            .I(N__6916));
    Span4Mux_v I__1328 (
            .O(N__6924),
            .I(N__6916));
    LocalMux I__1327 (
            .O(N__6921),
            .I(N__6913));
    Sp12to4 I__1326 (
            .O(N__6916),
            .I(N__6910));
    Span4Mux_v I__1325 (
            .O(N__6913),
            .I(N__6907));
    Span12Mux_h I__1324 (
            .O(N__6910),
            .I(N__6904));
    Sp12to4 I__1323 (
            .O(N__6907),
            .I(N__6901));
    Span12Mux_v I__1322 (
            .O(N__6904),
            .I(N__6896));
    Span12Mux_h I__1321 (
            .O(N__6901),
            .I(N__6896));
    Odrv12 I__1320 (
            .O(N__6896),
            .I(RnW_c));
    InMux I__1319 (
            .O(N__6893),
            .I(N__6888));
    InMux I__1318 (
            .O(N__6892),
            .I(N__6885));
    CascadeMux I__1317 (
            .O(N__6891),
            .I(N__6879));
    LocalMux I__1316 (
            .O(N__6888),
            .I(N__6874));
    LocalMux I__1315 (
            .O(N__6885),
            .I(N__6874));
    InMux I__1314 (
            .O(N__6884),
            .I(N__6871));
    InMux I__1313 (
            .O(N__6883),
            .I(N__6868));
    CascadeMux I__1312 (
            .O(N__6882),
            .I(N__6864));
    InMux I__1311 (
            .O(N__6879),
            .I(N__6861));
    Span12Mux_h I__1310 (
            .O(N__6874),
            .I(N__6858));
    LocalMux I__1309 (
            .O(N__6871),
            .I(N__6852));
    LocalMux I__1308 (
            .O(N__6868),
            .I(N__6852));
    InMux I__1307 (
            .O(N__6867),
            .I(N__6849));
    InMux I__1306 (
            .O(N__6864),
            .I(N__6843));
    LocalMux I__1305 (
            .O(N__6861),
            .I(N__6840));
    Span12Mux_v I__1304 (
            .O(N__6858),
            .I(N__6837));
    InMux I__1303 (
            .O(N__6857),
            .I(N__6834));
    Span4Mux_v I__1302 (
            .O(N__6852),
            .I(N__6829));
    LocalMux I__1301 (
            .O(N__6849),
            .I(N__6829));
    InMux I__1300 (
            .O(N__6848),
            .I(N__6826));
    InMux I__1299 (
            .O(N__6847),
            .I(N__6821));
    InMux I__1298 (
            .O(N__6846),
            .I(N__6821));
    LocalMux I__1297 (
            .O(N__6843),
            .I(N__6816));
    Span4Mux_v I__1296 (
            .O(N__6840),
            .I(N__6816));
    Odrv12 I__1295 (
            .O(N__6837),
            .I(WRITE_CYCLEm));
    LocalMux I__1294 (
            .O(N__6834),
            .I(WRITE_CYCLEm));
    Odrv4 I__1293 (
            .O(N__6829),
            .I(WRITE_CYCLEm));
    LocalMux I__1292 (
            .O(N__6826),
            .I(WRITE_CYCLEm));
    LocalMux I__1291 (
            .O(N__6821),
            .I(WRITE_CYCLEm));
    Odrv4 I__1290 (
            .O(N__6816),
            .I(WRITE_CYCLEm));
    IoInMux I__1289 (
            .O(N__6803),
            .I(N__6800));
    LocalMux I__1288 (
            .O(N__6800),
            .I(N__6797));
    IoSpan4Mux I__1287 (
            .O(N__6797),
            .I(N__6794));
    IoSpan4Mux I__1286 (
            .O(N__6794),
            .I(N__6791));
    Sp12to4 I__1285 (
            .O(N__6791),
            .I(N__6788));
    Span12Mux_s7_h I__1284 (
            .O(N__6788),
            .I(N__6785));
    Odrv12 I__1283 (
            .O(N__6785),
            .I(N_276));
    InMux I__1282 (
            .O(N__6782),
            .I(N__6779));
    LocalMux I__1281 (
            .O(N__6779),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1280 (
            .O(N__6776),
            .I(N__6770));
    InMux I__1279 (
            .O(N__6775),
            .I(N__6767));
    InMux I__1278 (
            .O(N__6774),
            .I(N__6758));
    InMux I__1277 (
            .O(N__6773),
            .I(N__6755));
    LocalMux I__1276 (
            .O(N__6770),
            .I(N__6749));
    LocalMux I__1275 (
            .O(N__6767),
            .I(N__6746));
    InMux I__1274 (
            .O(N__6766),
            .I(N__6743));
    InMux I__1273 (
            .O(N__6765),
            .I(N__6738));
    InMux I__1272 (
            .O(N__6764),
            .I(N__6738));
    InMux I__1271 (
            .O(N__6763),
            .I(N__6731));
    InMux I__1270 (
            .O(N__6762),
            .I(N__6731));
    InMux I__1269 (
            .O(N__6761),
            .I(N__6728));
    LocalMux I__1268 (
            .O(N__6758),
            .I(N__6725));
    LocalMux I__1267 (
            .O(N__6755),
            .I(N__6715));
    InMux I__1266 (
            .O(N__6754),
            .I(N__6712));
    InMux I__1265 (
            .O(N__6753),
            .I(N__6709));
    InMux I__1264 (
            .O(N__6752),
            .I(N__6706));
    Span4Mux_v I__1263 (
            .O(N__6749),
            .I(N__6699));
    Span4Mux_v I__1262 (
            .O(N__6746),
            .I(N__6699));
    LocalMux I__1261 (
            .O(N__6743),
            .I(N__6699));
    LocalMux I__1260 (
            .O(N__6738),
            .I(N__6696));
    InMux I__1259 (
            .O(N__6737),
            .I(N__6691));
    InMux I__1258 (
            .O(N__6736),
            .I(N__6691));
    LocalMux I__1257 (
            .O(N__6731),
            .I(N__6684));
    LocalMux I__1256 (
            .O(N__6728),
            .I(N__6684));
    Span4Mux_h I__1255 (
            .O(N__6725),
            .I(N__6684));
    InMux I__1254 (
            .O(N__6724),
            .I(N__6681));
    InMux I__1253 (
            .O(N__6723),
            .I(N__6678));
    InMux I__1252 (
            .O(N__6722),
            .I(N__6673));
    InMux I__1251 (
            .O(N__6721),
            .I(N__6673));
    InMux I__1250 (
            .O(N__6720),
            .I(N__6666));
    InMux I__1249 (
            .O(N__6719),
            .I(N__6666));
    InMux I__1248 (
            .O(N__6718),
            .I(N__6666));
    Odrv4 I__1247 (
            .O(N__6715),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1246 (
            .O(N__6712),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1245 (
            .O(N__6709),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1244 (
            .O(N__6706),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1243 (
            .O(N__6699),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1242 (
            .O(N__6696),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1241 (
            .O(N__6691),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1240 (
            .O(N__6684),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1239 (
            .O(N__6681),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1238 (
            .O(N__6678),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1237 (
            .O(N__6673),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1236 (
            .O(N__6666),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1235 (
            .O(N__6641),
            .I(N__6638));
    LocalMux I__1234 (
            .O(N__6638),
            .I(N__6635));
    Span4Mux_h I__1233 (
            .O(N__6635),
            .I(N__6632));
    Odrv4 I__1232 (
            .O(N__6632),
            .I(\U712_CHIP_RAM.N_300 ));
    CascadeMux I__1231 (
            .O(N__6629),
            .I(N__6625));
    CascadeMux I__1230 (
            .O(N__6628),
            .I(N__6622));
    InMux I__1229 (
            .O(N__6625),
            .I(N__6615));
    InMux I__1228 (
            .O(N__6622),
            .I(N__6610));
    InMux I__1227 (
            .O(N__6621),
            .I(N__6610));
    CascadeMux I__1226 (
            .O(N__6620),
            .I(N__6605));
    CascadeMux I__1225 (
            .O(N__6619),
            .I(N__6597));
    InMux I__1224 (
            .O(N__6618),
            .I(N__6593));
    LocalMux I__1223 (
            .O(N__6615),
            .I(N__6589));
    LocalMux I__1222 (
            .O(N__6610),
            .I(N__6586));
    InMux I__1221 (
            .O(N__6609),
            .I(N__6581));
    InMux I__1220 (
            .O(N__6608),
            .I(N__6576));
    InMux I__1219 (
            .O(N__6605),
            .I(N__6576));
    InMux I__1218 (
            .O(N__6604),
            .I(N__6571));
    InMux I__1217 (
            .O(N__6603),
            .I(N__6571));
    CascadeMux I__1216 (
            .O(N__6602),
            .I(N__6568));
    CascadeMux I__1215 (
            .O(N__6601),
            .I(N__6564));
    InMux I__1214 (
            .O(N__6600),
            .I(N__6561));
    InMux I__1213 (
            .O(N__6597),
            .I(N__6558));
    InMux I__1212 (
            .O(N__6596),
            .I(N__6555));
    LocalMux I__1211 (
            .O(N__6593),
            .I(N__6552));
    CascadeMux I__1210 (
            .O(N__6592),
            .I(N__6545));
    Span4Mux_v I__1209 (
            .O(N__6589),
            .I(N__6539));
    Span4Mux_v I__1208 (
            .O(N__6586),
            .I(N__6539));
    InMux I__1207 (
            .O(N__6585),
            .I(N__6536));
    InMux I__1206 (
            .O(N__6584),
            .I(N__6533));
    LocalMux I__1205 (
            .O(N__6581),
            .I(N__6528));
    LocalMux I__1204 (
            .O(N__6576),
            .I(N__6528));
    LocalMux I__1203 (
            .O(N__6571),
            .I(N__6525));
    InMux I__1202 (
            .O(N__6568),
            .I(N__6522));
    InMux I__1201 (
            .O(N__6567),
            .I(N__6517));
    InMux I__1200 (
            .O(N__6564),
            .I(N__6517));
    LocalMux I__1199 (
            .O(N__6561),
            .I(N__6508));
    LocalMux I__1198 (
            .O(N__6558),
            .I(N__6508));
    LocalMux I__1197 (
            .O(N__6555),
            .I(N__6508));
    Span4Mux_h I__1196 (
            .O(N__6552),
            .I(N__6508));
    InMux I__1195 (
            .O(N__6551),
            .I(N__6505));
    InMux I__1194 (
            .O(N__6550),
            .I(N__6500));
    InMux I__1193 (
            .O(N__6549),
            .I(N__6500));
    InMux I__1192 (
            .O(N__6548),
            .I(N__6493));
    InMux I__1191 (
            .O(N__6545),
            .I(N__6493));
    InMux I__1190 (
            .O(N__6544),
            .I(N__6493));
    Odrv4 I__1189 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1188 (
            .O(N__6536),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1187 (
            .O(N__6533),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1186 (
            .O(N__6528),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1185 (
            .O(N__6525),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1184 (
            .O(N__6522),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1183 (
            .O(N__6517),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1182 (
            .O(N__6508),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1181 (
            .O(N__6505),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1180 (
            .O(N__6500),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1179 (
            .O(N__6493),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1178 (
            .O(N__6470),
            .I(N__6461));
    InMux I__1177 (
            .O(N__6469),
            .I(N__6457));
    CascadeMux I__1176 (
            .O(N__6468),
            .I(N__6454));
    CascadeMux I__1175 (
            .O(N__6467),
            .I(N__6450));
    InMux I__1174 (
            .O(N__6466),
            .I(N__6447));
    InMux I__1173 (
            .O(N__6465),
            .I(N__6444));
    InMux I__1172 (
            .O(N__6464),
            .I(N__6439));
    LocalMux I__1171 (
            .O(N__6461),
            .I(N__6436));
    InMux I__1170 (
            .O(N__6460),
            .I(N__6432));
    LocalMux I__1169 (
            .O(N__6457),
            .I(N__6429));
    InMux I__1168 (
            .O(N__6454),
            .I(N__6426));
    InMux I__1167 (
            .O(N__6453),
            .I(N__6422));
    InMux I__1166 (
            .O(N__6450),
            .I(N__6419));
    LocalMux I__1165 (
            .O(N__6447),
            .I(N__6414));
    LocalMux I__1164 (
            .O(N__6444),
            .I(N__6414));
    InMux I__1163 (
            .O(N__6443),
            .I(N__6411));
    InMux I__1162 (
            .O(N__6442),
            .I(N__6408));
    LocalMux I__1161 (
            .O(N__6439),
            .I(N__6403));
    Span4Mux_v I__1160 (
            .O(N__6436),
            .I(N__6403));
    InMux I__1159 (
            .O(N__6435),
            .I(N__6400));
    LocalMux I__1158 (
            .O(N__6432),
            .I(N__6393));
    Span4Mux_h I__1157 (
            .O(N__6429),
            .I(N__6393));
    LocalMux I__1156 (
            .O(N__6426),
            .I(N__6393));
    InMux I__1155 (
            .O(N__6425),
            .I(N__6390));
    LocalMux I__1154 (
            .O(N__6422),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1153 (
            .O(N__6419),
            .I(\U712_CHIP_RAM.N_241 ));
    Odrv4 I__1152 (
            .O(N__6414),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1151 (
            .O(N__6411),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1150 (
            .O(N__6408),
            .I(\U712_CHIP_RAM.N_241 ));
    Odrv4 I__1149 (
            .O(N__6403),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1148 (
            .O(N__6400),
            .I(\U712_CHIP_RAM.N_241 ));
    Odrv4 I__1147 (
            .O(N__6393),
            .I(\U712_CHIP_RAM.N_241 ));
    LocalMux I__1146 (
            .O(N__6390),
            .I(\U712_CHIP_RAM.N_241 ));
    CascadeMux I__1145 (
            .O(N__6371),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    InMux I__1144 (
            .O(N__6368),
            .I(N__6356));
    InMux I__1143 (
            .O(N__6367),
            .I(N__6353));
    InMux I__1142 (
            .O(N__6366),
            .I(N__6350));
    InMux I__1141 (
            .O(N__6365),
            .I(N__6345));
    InMux I__1140 (
            .O(N__6364),
            .I(N__6342));
    InMux I__1139 (
            .O(N__6363),
            .I(N__6339));
    InMux I__1138 (
            .O(N__6362),
            .I(N__6334));
    InMux I__1137 (
            .O(N__6361),
            .I(N__6334));
    InMux I__1136 (
            .O(N__6360),
            .I(N__6331));
    InMux I__1135 (
            .O(N__6359),
            .I(N__6328));
    LocalMux I__1134 (
            .O(N__6356),
            .I(N__6323));
    LocalMux I__1133 (
            .O(N__6353),
            .I(N__6318));
    LocalMux I__1132 (
            .O(N__6350),
            .I(N__6318));
    InMux I__1131 (
            .O(N__6349),
            .I(N__6315));
    InMux I__1130 (
            .O(N__6348),
            .I(N__6312));
    LocalMux I__1129 (
            .O(N__6345),
            .I(N__6305));
    LocalMux I__1128 (
            .O(N__6342),
            .I(N__6305));
    LocalMux I__1127 (
            .O(N__6339),
            .I(N__6300));
    LocalMux I__1126 (
            .O(N__6334),
            .I(N__6300));
    LocalMux I__1125 (
            .O(N__6331),
            .I(N__6295));
    LocalMux I__1124 (
            .O(N__6328),
            .I(N__6295));
    InMux I__1123 (
            .O(N__6327),
            .I(N__6290));
    InMux I__1122 (
            .O(N__6326),
            .I(N__6287));
    Span4Mux_v I__1121 (
            .O(N__6323),
            .I(N__6284));
    Span4Mux_h I__1120 (
            .O(N__6318),
            .I(N__6281));
    LocalMux I__1119 (
            .O(N__6315),
            .I(N__6276));
    LocalMux I__1118 (
            .O(N__6312),
            .I(N__6276));
    InMux I__1117 (
            .O(N__6311),
            .I(N__6271));
    InMux I__1116 (
            .O(N__6310),
            .I(N__6271));
    Span4Mux_v I__1115 (
            .O(N__6305),
            .I(N__6264));
    Span4Mux_h I__1114 (
            .O(N__6300),
            .I(N__6264));
    Span4Mux_v I__1113 (
            .O(N__6295),
            .I(N__6264));
    InMux I__1112 (
            .O(N__6294),
            .I(N__6259));
    InMux I__1111 (
            .O(N__6293),
            .I(N__6259));
    LocalMux I__1110 (
            .O(N__6290),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1109 (
            .O(N__6287),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1108 (
            .O(N__6284),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1107 (
            .O(N__6281),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1106 (
            .O(N__6276),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1105 (
            .O(N__6271),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1104 (
            .O(N__6264),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1103 (
            .O(N__6259),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1102 (
            .O(N__6242),
            .I(N__6239));
    LocalMux I__1101 (
            .O(N__6239),
            .I(N__6236));
    Span4Mux_v I__1100 (
            .O(N__6236),
            .I(N__6233));
    Sp12to4 I__1099 (
            .O(N__6233),
            .I(N__6230));
    Span12Mux_h I__1098 (
            .O(N__6230),
            .I(N__6227));
    Odrv12 I__1097 (
            .O(N__6227),
            .I(A_c_9));
    InMux I__1096 (
            .O(N__6224),
            .I(N__6221));
    LocalMux I__1095 (
            .O(N__6221),
            .I(N__6218));
    Span4Mux_h I__1094 (
            .O(N__6218),
            .I(N__6215));
    Sp12to4 I__1093 (
            .O(N__6215),
            .I(N__6212));
    Span12Mux_v I__1092 (
            .O(N__6212),
            .I(N__6209));
    Odrv12 I__1091 (
            .O(N__6209),
            .I(A_c_2));
    InMux I__1090 (
            .O(N__6206),
            .I(N__6202));
    InMux I__1089 (
            .O(N__6205),
            .I(N__6198));
    LocalMux I__1088 (
            .O(N__6202),
            .I(N__6195));
    InMux I__1087 (
            .O(N__6201),
            .I(N__6192));
    LocalMux I__1086 (
            .O(N__6198),
            .I(N__6189));
    Odrv4 I__1085 (
            .O(N__6195),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1084 (
            .O(N__6192),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__1083 (
            .O(N__6189),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__1082 (
            .O(N__6182),
            .I(\U712_REG_SM.N_360_1_cascade_ ));
    CascadeMux I__1081 (
            .O(N__6179),
            .I(N__6175));
    InMux I__1080 (
            .O(N__6178),
            .I(N__6170));
    InMux I__1079 (
            .O(N__6175),
            .I(N__6170));
    LocalMux I__1078 (
            .O(N__6170),
            .I(\U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1 ));
    CascadeMux I__1077 (
            .O(N__6167),
            .I(\U712_REG_SM.m17_i_0_o2_cascade_ ));
    CascadeMux I__1076 (
            .O(N__6164),
            .I(\U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_ ));
    InMux I__1075 (
            .O(N__6161),
            .I(N__6158));
    LocalMux I__1074 (
            .O(N__6158),
            .I(N__6152));
    InMux I__1073 (
            .O(N__6157),
            .I(N__6149));
    InMux I__1072 (
            .O(N__6156),
            .I(N__6146));
    InMux I__1071 (
            .O(N__6155),
            .I(N__6143));
    Odrv12 I__1070 (
            .O(N__6152),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1069 (
            .O(N__6149),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1068 (
            .O(N__6146),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1067 (
            .O(N__6143),
            .I(\U712_CHIP_RAM.N_388 ));
    CascadeMux I__1066 (
            .O(N__6134),
            .I(N__6129));
    InMux I__1065 (
            .O(N__6133),
            .I(N__6125));
    InMux I__1064 (
            .O(N__6132),
            .I(N__6122));
    InMux I__1063 (
            .O(N__6129),
            .I(N__6119));
    CascadeMux I__1062 (
            .O(N__6128),
            .I(N__6116));
    LocalMux I__1061 (
            .O(N__6125),
            .I(N__6112));
    LocalMux I__1060 (
            .O(N__6122),
            .I(N__6107));
    LocalMux I__1059 (
            .O(N__6119),
            .I(N__6107));
    InMux I__1058 (
            .O(N__6116),
            .I(N__6102));
    InMux I__1057 (
            .O(N__6115),
            .I(N__6102));
    Odrv4 I__1056 (
            .O(N__6112),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1055 (
            .O(N__6107),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1054 (
            .O(N__6102),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1053 (
            .O(N__6095),
            .I(N__6089));
    InMux I__1052 (
            .O(N__6094),
            .I(N__6086));
    InMux I__1051 (
            .O(N__6093),
            .I(N__6083));
    CascadeMux I__1050 (
            .O(N__6092),
            .I(N__6080));
    LocalMux I__1049 (
            .O(N__6089),
            .I(N__6073));
    LocalMux I__1048 (
            .O(N__6086),
            .I(N__6073));
    LocalMux I__1047 (
            .O(N__6083),
            .I(N__6070));
    InMux I__1046 (
            .O(N__6080),
            .I(N__6063));
    InMux I__1045 (
            .O(N__6079),
            .I(N__6063));
    InMux I__1044 (
            .O(N__6078),
            .I(N__6060));
    Span4Mux_h I__1043 (
            .O(N__6073),
            .I(N__6055));
    Span4Mux_h I__1042 (
            .O(N__6070),
            .I(N__6055));
    InMux I__1041 (
            .O(N__6069),
            .I(N__6050));
    InMux I__1040 (
            .O(N__6068),
            .I(N__6050));
    LocalMux I__1039 (
            .O(N__6063),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1038 (
            .O(N__6060),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1037 (
            .O(N__6055),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1036 (
            .O(N__6050),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1035 (
            .O(N__6041),
            .I(\U712_CHIP_RAM.N_271_cascade_ ));
    InMux I__1034 (
            .O(N__6038),
            .I(N__6035));
    LocalMux I__1033 (
            .O(N__6035),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ));
    CascadeMux I__1032 (
            .O(N__6032),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ));
    InMux I__1031 (
            .O(N__6029),
            .I(N__6026));
    LocalMux I__1030 (
            .O(N__6026),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1 ));
    InMux I__1029 (
            .O(N__6023),
            .I(N__6020));
    LocalMux I__1028 (
            .O(N__6020),
            .I(\U712_CHIP_RAM.N_317 ));
    CascadeMux I__1027 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ));
    InMux I__1026 (
            .O(N__6014),
            .I(N__6010));
    InMux I__1025 (
            .O(N__6013),
            .I(N__6007));
    LocalMux I__1024 (
            .O(N__6010),
            .I(\U712_CHIP_RAM.N_434 ));
    LocalMux I__1023 (
            .O(N__6007),
            .I(\U712_CHIP_RAM.N_434 ));
    InMux I__1022 (
            .O(N__6002),
            .I(N__5999));
    LocalMux I__1021 (
            .O(N__5999),
            .I(\U712_CHIP_RAM.N_13 ));
    InMux I__1020 (
            .O(N__5996),
            .I(N__5993));
    LocalMux I__1019 (
            .O(N__5993),
            .I(N__5990));
    Span4Mux_v I__1018 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_v I__1017 (
            .O(N__5987),
            .I(N__5984));
    Sp12to4 I__1016 (
            .O(N__5984),
            .I(N__5981));
    Span12Mux_h I__1015 (
            .O(N__5981),
            .I(N__5978));
    Odrv12 I__1014 (
            .O(N__5978),
            .I(A_c_15));
    InMux I__1013 (
            .O(N__5975),
            .I(N__5972));
    LocalMux I__1012 (
            .O(N__5972),
            .I(N__5969));
    Span12Mux_v I__1011 (
            .O(N__5969),
            .I(N__5966));
    Span12Mux_h I__1010 (
            .O(N__5966),
            .I(N__5963));
    Odrv12 I__1009 (
            .O(N__5963),
            .I(A_c_8));
    InMux I__1008 (
            .O(N__5960),
            .I(N__5949));
    InMux I__1007 (
            .O(N__5959),
            .I(N__5946));
    InMux I__1006 (
            .O(N__5958),
            .I(N__5943));
    InMux I__1005 (
            .O(N__5957),
            .I(N__5940));
    InMux I__1004 (
            .O(N__5956),
            .I(N__5934));
    InMux I__1003 (
            .O(N__5955),
            .I(N__5931));
    CascadeMux I__1002 (
            .O(N__5954),
            .I(N__5927));
    InMux I__1001 (
            .O(N__5953),
            .I(N__5922));
    InMux I__1000 (
            .O(N__5952),
            .I(N__5922));
    LocalMux I__999 (
            .O(N__5949),
            .I(N__5917));
    LocalMux I__998 (
            .O(N__5946),
            .I(N__5917));
    LocalMux I__997 (
            .O(N__5943),
            .I(N__5914));
    LocalMux I__996 (
            .O(N__5940),
            .I(N__5911));
    InMux I__995 (
            .O(N__5939),
            .I(N__5904));
    InMux I__994 (
            .O(N__5938),
            .I(N__5904));
    InMux I__993 (
            .O(N__5937),
            .I(N__5904));
    LocalMux I__992 (
            .O(N__5934),
            .I(N__5897));
    LocalMux I__991 (
            .O(N__5931),
            .I(N__5897));
    InMux I__990 (
            .O(N__5930),
            .I(N__5891));
    InMux I__989 (
            .O(N__5927),
            .I(N__5888));
    LocalMux I__988 (
            .O(N__5922),
            .I(N__5885));
    Span4Mux_v I__987 (
            .O(N__5917),
            .I(N__5876));
    Span4Mux_v I__986 (
            .O(N__5914),
            .I(N__5876));
    Span4Mux_h I__985 (
            .O(N__5911),
            .I(N__5876));
    LocalMux I__984 (
            .O(N__5904),
            .I(N__5876));
    InMux I__983 (
            .O(N__5903),
            .I(N__5873));
    InMux I__982 (
            .O(N__5902),
            .I(N__5870));
    Span4Mux_h I__981 (
            .O(N__5897),
            .I(N__5867));
    InMux I__980 (
            .O(N__5896),
            .I(N__5860));
    InMux I__979 (
            .O(N__5895),
            .I(N__5860));
    InMux I__978 (
            .O(N__5894),
            .I(N__5860));
    LocalMux I__977 (
            .O(N__5891),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__976 (
            .O(N__5888),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__975 (
            .O(N__5885),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__974 (
            .O(N__5876),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__973 (
            .O(N__5873),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__972 (
            .O(N__5870),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__971 (
            .O(N__5867),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__970 (
            .O(N__5860),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__969 (
            .O(N__5843),
            .I(N__5835));
    InMux I__968 (
            .O(N__5842),
            .I(N__5830));
    InMux I__967 (
            .O(N__5841),
            .I(N__5830));
    InMux I__966 (
            .O(N__5840),
            .I(N__5827));
    InMux I__965 (
            .O(N__5839),
            .I(N__5824));
    InMux I__964 (
            .O(N__5838),
            .I(N__5819));
    LocalMux I__963 (
            .O(N__5835),
            .I(N__5814));
    LocalMux I__962 (
            .O(N__5830),
            .I(N__5811));
    LocalMux I__961 (
            .O(N__5827),
            .I(N__5808));
    LocalMux I__960 (
            .O(N__5824),
            .I(N__5805));
    InMux I__959 (
            .O(N__5823),
            .I(N__5800));
    InMux I__958 (
            .O(N__5822),
            .I(N__5800));
    LocalMux I__957 (
            .O(N__5819),
            .I(N__5793));
    InMux I__956 (
            .O(N__5818),
            .I(N__5788));
    InMux I__955 (
            .O(N__5817),
            .I(N__5788));
    Span4Mux_v I__954 (
            .O(N__5814),
            .I(N__5777));
    Span4Mux_v I__953 (
            .O(N__5811),
            .I(N__5777));
    Span4Mux_v I__952 (
            .O(N__5808),
            .I(N__5777));
    Span4Mux_h I__951 (
            .O(N__5805),
            .I(N__5777));
    LocalMux I__950 (
            .O(N__5800),
            .I(N__5777));
    InMux I__949 (
            .O(N__5799),
            .I(N__5774));
    InMux I__948 (
            .O(N__5798),
            .I(N__5767));
    InMux I__947 (
            .O(N__5797),
            .I(N__5767));
    InMux I__946 (
            .O(N__5796),
            .I(N__5767));
    Odrv4 I__945 (
            .O(N__5793),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__944 (
            .O(N__5788),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__943 (
            .O(N__5777),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__942 (
            .O(N__5774),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__941 (
            .O(N__5767),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__940 (
            .O(N__5756),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_ ));
    CascadeMux I__939 (
            .O(N__5753),
            .I(\U712_BYTE_ENABLE.N_374_cascade_ ));
    IoInMux I__938 (
            .O(N__5750),
            .I(N__5747));
    LocalMux I__937 (
            .O(N__5747),
            .I(N__5744));
    Span4Mux_s0_v I__936 (
            .O(N__5744),
            .I(N__5741));
    Sp12to4 I__935 (
            .O(N__5741),
            .I(N__5738));
    Span12Mux_h I__934 (
            .O(N__5738),
            .I(N__5735));
    Span12Mux_v I__933 (
            .O(N__5735),
            .I(N__5732));
    Odrv12 I__932 (
            .O(N__5732),
            .I(N_51_i));
    IoInMux I__931 (
            .O(N__5729),
            .I(N__5726));
    LocalMux I__930 (
            .O(N__5726),
            .I(N__5723));
    IoSpan4Mux I__929 (
            .O(N__5723),
            .I(N__5719));
    InMux I__928 (
            .O(N__5722),
            .I(N__5716));
    Span4Mux_s2_v I__927 (
            .O(N__5719),
            .I(N__5713));
    LocalMux I__926 (
            .O(N__5716),
            .I(N__5710));
    Span4Mux_v I__925 (
            .O(N__5713),
            .I(N__5705));
    Span4Mux_v I__924 (
            .O(N__5710),
            .I(N__5705));
    Odrv4 I__923 (
            .O(N__5705),
            .I(CONSTANT_ONE_NET));
    InMux I__922 (
            .O(N__5702),
            .I(N__5699));
    LocalMux I__921 (
            .O(N__5699),
            .I(N__5696));
    Span12Mux_s11_v I__920 (
            .O(N__5696),
            .I(N__5693));
    Span12Mux_h I__919 (
            .O(N__5693),
            .I(N__5690));
    Odrv12 I__918 (
            .O(N__5690),
            .I(A_c_10));
    InMux I__917 (
            .O(N__5687),
            .I(N__5684));
    LocalMux I__916 (
            .O(N__5684),
            .I(N__5681));
    Span12Mux_v I__915 (
            .O(N__5681),
            .I(N__5678));
    Span12Mux_h I__914 (
            .O(N__5678),
            .I(N__5675));
    Span12Mux_v I__913 (
            .O(N__5675),
            .I(N__5672));
    Odrv12 I__912 (
            .O(N__5672),
            .I(A_c_3));
    CascadeMux I__911 (
            .O(N__5669),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_ ));
    CascadeMux I__910 (
            .O(N__5666),
            .I(\U712_CHIP_RAM.N_322_cascade_ ));
    InMux I__909 (
            .O(N__5663),
            .I(N__5660));
    LocalMux I__908 (
            .O(N__5660),
            .I(N__5657));
    Odrv4 I__907 (
            .O(N__5657),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ));
    CEMux I__906 (
            .O(N__5654),
            .I(N__5651));
    LocalMux I__905 (
            .O(N__5651),
            .I(N__5647));
    CEMux I__904 (
            .O(N__5650),
            .I(N__5644));
    Span4Mux_v I__903 (
            .O(N__5647),
            .I(N__5641));
    LocalMux I__902 (
            .O(N__5644),
            .I(N__5638));
    Span4Mux_h I__901 (
            .O(N__5641),
            .I(N__5635));
    Span4Mux_v I__900 (
            .O(N__5638),
            .I(N__5632));
    Odrv4 I__899 (
            .O(N__5635),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    Odrv4 I__898 (
            .O(N__5632),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    InMux I__897 (
            .O(N__5627),
            .I(N__5624));
    LocalMux I__896 (
            .O(N__5624),
            .I(\U712_REG_SM.N_289 ));
    CascadeMux I__895 (
            .O(N__5621),
            .I(\U712_REG_SM.N_358_cascade_ ));
    InMux I__894 (
            .O(N__5618),
            .I(N__5615));
    LocalMux I__893 (
            .O(N__5615),
            .I(\U712_REG_SM.N_360 ));
    InMux I__892 (
            .O(N__5612),
            .I(N__5608));
    InMux I__891 (
            .O(N__5611),
            .I(N__5605));
    LocalMux I__890 (
            .O(N__5608),
            .I(\U712_REG_SM.N_359 ));
    LocalMux I__889 (
            .O(N__5605),
            .I(\U712_REG_SM.N_359 ));
    InMux I__888 (
            .O(N__5600),
            .I(N__5597));
    LocalMux I__887 (
            .O(N__5597),
            .I(\U712_REG_SM.N_270_i ));
    InMux I__886 (
            .O(N__5594),
            .I(N__5591));
    LocalMux I__885 (
            .O(N__5591),
            .I(\U712_REG_SM.REG_TACK_7 ));
    CascadeMux I__884 (
            .O(N__5588),
            .I(N__5584));
    InMux I__883 (
            .O(N__5587),
            .I(N__5581));
    InMux I__882 (
            .O(N__5584),
            .I(N__5577));
    LocalMux I__881 (
            .O(N__5581),
            .I(N__5574));
    InMux I__880 (
            .O(N__5580),
            .I(N__5571));
    LocalMux I__879 (
            .O(N__5577),
            .I(REG_TACK));
    Odrv4 I__878 (
            .O(N__5574),
            .I(REG_TACK));
    LocalMux I__877 (
            .O(N__5571),
            .I(REG_TACK));
    InMux I__876 (
            .O(N__5564),
            .I(N__5561));
    LocalMux I__875 (
            .O(N__5561),
            .I(N__5557));
    IoInMux I__874 (
            .O(N__5560),
            .I(N__5554));
    Span4Mux_v I__873 (
            .O(N__5557),
            .I(N__5551));
    LocalMux I__872 (
            .O(N__5554),
            .I(N__5548));
    Sp12to4 I__871 (
            .O(N__5551),
            .I(N__5545));
    IoSpan4Mux I__870 (
            .O(N__5548),
            .I(N__5542));
    Span12Mux_h I__869 (
            .O(N__5545),
            .I(N__5539));
    IoSpan4Mux I__868 (
            .O(N__5542),
            .I(N__5536));
    Span12Mux_v I__867 (
            .O(N__5539),
            .I(N__5533));
    IoSpan4Mux I__866 (
            .O(N__5536),
            .I(N__5530));
    Odrv12 I__865 (
            .O(N__5533),
            .I(C1_c));
    Odrv4 I__864 (
            .O(N__5530),
            .I(C1_c));
    CascadeMux I__863 (
            .O(N__5525),
            .I(\U712_REG_SM.N_340_cascade_ ));
    InMux I__862 (
            .O(N__5522),
            .I(N__5519));
    LocalMux I__861 (
            .O(N__5519),
            .I(N__5516));
    Span4Mux_h I__860 (
            .O(N__5516),
            .I(N__5513));
    Span4Mux_h I__859 (
            .O(N__5513),
            .I(N__5510));
    Sp12to4 I__858 (
            .O(N__5510),
            .I(N__5507));
    Span12Mux_v I__857 (
            .O(N__5507),
            .I(N__5504));
    Odrv12 I__856 (
            .O(N__5504),
            .I(REGSPACEn_c));
    IoInMux I__855 (
            .O(N__5501),
            .I(N__5498));
    LocalMux I__854 (
            .O(N__5498),
            .I(N__5493));
    InMux I__853 (
            .O(N__5497),
            .I(N__5490));
    InMux I__852 (
            .O(N__5496),
            .I(N__5487));
    Span4Mux_s3_v I__851 (
            .O(N__5493),
            .I(N__5484));
    LocalMux I__850 (
            .O(N__5490),
            .I(N__5479));
    LocalMux I__849 (
            .O(N__5487),
            .I(N__5479));
    Span4Mux_v I__848 (
            .O(N__5484),
            .I(N__5476));
    Span4Mux_v I__847 (
            .O(N__5479),
            .I(N__5473));
    Span4Mux_v I__846 (
            .O(N__5476),
            .I(N__5469));
    Span4Mux_v I__845 (
            .O(N__5473),
            .I(N__5466));
    InMux I__844 (
            .O(N__5472),
            .I(N__5463));
    Odrv4 I__843 (
            .O(N__5469),
            .I(DBENn_c));
    Odrv4 I__842 (
            .O(N__5466),
            .I(DBENn_c));
    LocalMux I__841 (
            .O(N__5463),
            .I(DBENn_c));
    InMux I__840 (
            .O(N__5456),
            .I(N__5452));
    InMux I__839 (
            .O(N__5455),
            .I(N__5449));
    LocalMux I__838 (
            .O(N__5452),
            .I(N__5443));
    LocalMux I__837 (
            .O(N__5449),
            .I(N__5443));
    InMux I__836 (
            .O(N__5448),
            .I(N__5439));
    Span4Mux_v I__835 (
            .O(N__5443),
            .I(N__5436));
    InMux I__834 (
            .O(N__5442),
            .I(N__5432));
    LocalMux I__833 (
            .O(N__5439),
            .I(N__5428));
    Span4Mux_v I__832 (
            .O(N__5436),
            .I(N__5425));
    InMux I__831 (
            .O(N__5435),
            .I(N__5422));
    LocalMux I__830 (
            .O(N__5432),
            .I(N__5419));
    InMux I__829 (
            .O(N__5431),
            .I(N__5416));
    Span4Mux_h I__828 (
            .O(N__5428),
            .I(N__5413));
    Odrv4 I__827 (
            .O(N__5425),
            .I(DMA_CYCLEm));
    LocalMux I__826 (
            .O(N__5422),
            .I(DMA_CYCLEm));
    Odrv12 I__825 (
            .O(N__5419),
            .I(DMA_CYCLEm));
    LocalMux I__824 (
            .O(N__5416),
            .I(DMA_CYCLEm));
    Odrv4 I__823 (
            .O(N__5413),
            .I(DMA_CYCLEm));
    InMux I__822 (
            .O(N__5402),
            .I(N__5398));
    InMux I__821 (
            .O(N__5401),
            .I(N__5395));
    LocalMux I__820 (
            .O(N__5398),
            .I(N__5390));
    LocalMux I__819 (
            .O(N__5395),
            .I(N__5390));
    Span4Mux_v I__818 (
            .O(N__5390),
            .I(N__5387));
    Sp12to4 I__817 (
            .O(N__5387),
            .I(N__5384));
    Span12Mux_h I__816 (
            .O(N__5384),
            .I(N__5381));
    Span12Mux_v I__815 (
            .O(N__5381),
            .I(N__5378));
    Odrv12 I__814 (
            .O(N__5378),
            .I(TSn_c));
    InMux I__813 (
            .O(N__5375),
            .I(N__5372));
    LocalMux I__812 (
            .O(N__5372),
            .I(N__5369));
    Span4Mux_h I__811 (
            .O(N__5369),
            .I(N__5366));
    Span4Mux_v I__810 (
            .O(N__5366),
            .I(N__5363));
    Span4Mux_v I__809 (
            .O(N__5363),
            .I(N__5360));
    Span4Mux_v I__808 (
            .O(N__5360),
            .I(N__5357));
    Odrv4 I__807 (
            .O(N__5357),
            .I(RAMSPACEn_c));
    InMux I__806 (
            .O(N__5354),
            .I(N__5351));
    LocalMux I__805 (
            .O(N__5351),
            .I(N__5348));
    Odrv12 I__804 (
            .O(N__5348),
            .I(\U712_CHIP_RAM.N_345 ));
    InMux I__803 (
            .O(N__5345),
            .I(N__5341));
    InMux I__802 (
            .O(N__5344),
            .I(N__5338));
    LocalMux I__801 (
            .O(N__5341),
            .I(DBR_SYNCZ0Z_0));
    LocalMux I__800 (
            .O(N__5338),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__799 (
            .O(N__5333),
            .I(N__5329));
    InMux I__798 (
            .O(N__5332),
            .I(N__5326));
    InMux I__797 (
            .O(N__5329),
            .I(N__5322));
    LocalMux I__796 (
            .O(N__5326),
            .I(N__5319));
    InMux I__795 (
            .O(N__5325),
            .I(N__5316));
    LocalMux I__794 (
            .O(N__5322),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__793 (
            .O(N__5319),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__792 (
            .O(N__5316),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__791 (
            .O(N__5309),
            .I(\U712_REG_SM.m17_i_0_o2_1_cascade_ ));
    InMux I__790 (
            .O(N__5306),
            .I(N__5303));
    LocalMux I__789 (
            .O(N__5303),
            .I(N__5300));
    Span4Mux_h I__788 (
            .O(N__5300),
            .I(N__5297));
    Span4Mux_v I__787 (
            .O(N__5297),
            .I(N__5294));
    Sp12to4 I__786 (
            .O(N__5294),
            .I(N__5291));
    Odrv12 I__785 (
            .O(N__5291),
            .I(A_c_7));
    CascadeMux I__784 (
            .O(N__5288),
            .I(\U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_ ));
    InMux I__783 (
            .O(N__5285),
            .I(N__5279));
    InMux I__782 (
            .O(N__5284),
            .I(N__5274));
    InMux I__781 (
            .O(N__5283),
            .I(N__5274));
    InMux I__780 (
            .O(N__5282),
            .I(N__5271));
    LocalMux I__779 (
            .O(N__5279),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__778 (
            .O(N__5274),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__777 (
            .O(N__5271),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__776 (
            .O(N__5264),
            .I(N__5257));
    InMux I__775 (
            .O(N__5263),
            .I(N__5252));
    InMux I__774 (
            .O(N__5262),
            .I(N__5252));
    InMux I__773 (
            .O(N__5261),
            .I(N__5247));
    InMux I__772 (
            .O(N__5260),
            .I(N__5247));
    LocalMux I__771 (
            .O(N__5257),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__770 (
            .O(N__5252),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__769 (
            .O(N__5247),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__768 (
            .O(N__5240),
            .I(\U712_REG_SM.m15_i_0_a2_0_0_cascade_ ));
    InMux I__767 (
            .O(N__5237),
            .I(N__5234));
    LocalMux I__766 (
            .O(N__5234),
            .I(\U712_CHIP_RAM.N_386 ));
    CascadeMux I__765 (
            .O(N__5231),
            .I(\U712_CHIP_RAM.N_434_cascade_ ));
    InMux I__764 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__763 (
            .O(N__5225),
            .I(N__5222));
    Span4Mux_h I__762 (
            .O(N__5222),
            .I(N__5217));
    InMux I__761 (
            .O(N__5221),
            .I(N__5212));
    InMux I__760 (
            .O(N__5220),
            .I(N__5212));
    Odrv4 I__759 (
            .O(N__5217),
            .I(\U712_CHIP_RAM.N_439 ));
    LocalMux I__758 (
            .O(N__5212),
            .I(\U712_CHIP_RAM.N_439 ));
    InMux I__757 (
            .O(N__5207),
            .I(N__5204));
    LocalMux I__756 (
            .O(N__5204),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0 ));
    InMux I__755 (
            .O(N__5201),
            .I(N__5198));
    LocalMux I__754 (
            .O(N__5198),
            .I(\U712_CHIP_RAM.N_335 ));
    InMux I__753 (
            .O(N__5195),
            .I(N__5192));
    LocalMux I__752 (
            .O(N__5192),
            .I(N__5189));
    Span4Mux_v I__751 (
            .O(N__5189),
            .I(N__5186));
    Span4Mux_h I__750 (
            .O(N__5186),
            .I(N__5183));
    Sp12to4 I__749 (
            .O(N__5183),
            .I(N__5180));
    Odrv12 I__748 (
            .O(N__5180),
            .I(A_c_12));
    InMux I__747 (
            .O(N__5177),
            .I(N__5174));
    LocalMux I__746 (
            .O(N__5174),
            .I(N__5171));
    Span4Mux_h I__745 (
            .O(N__5171),
            .I(N__5168));
    Sp12to4 I__744 (
            .O(N__5168),
            .I(N__5165));
    Span12Mux_v I__743 (
            .O(N__5165),
            .I(N__5162));
    Odrv12 I__742 (
            .O(N__5162),
            .I(A_c_5));
    CascadeMux I__741 (
            .O(N__5159),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_ ));
    InMux I__740 (
            .O(N__5156),
            .I(N__5153));
    LocalMux I__739 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1 ));
    InMux I__738 (
            .O(N__5150),
            .I(N__5146));
    InMux I__737 (
            .O(N__5149),
            .I(N__5142));
    LocalMux I__736 (
            .O(N__5146),
            .I(N__5139));
    InMux I__735 (
            .O(N__5145),
            .I(N__5136));
    LocalMux I__734 (
            .O(N__5142),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__733 (
            .O(N__5139),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__732 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__731 (
            .O(N__5129),
            .I(N__5124));
    InMux I__730 (
            .O(N__5128),
            .I(N__5121));
    InMux I__729 (
            .O(N__5127),
            .I(N__5118));
    LocalMux I__728 (
            .O(N__5124),
            .I(N__5115));
    LocalMux I__727 (
            .O(N__5121),
            .I(CPU_TACKm));
    LocalMux I__726 (
            .O(N__5118),
            .I(CPU_TACKm));
    Odrv12 I__725 (
            .O(N__5115),
            .I(CPU_TACKm));
    CascadeMux I__724 (
            .O(N__5108),
            .I(N__5103));
    InMux I__723 (
            .O(N__5107),
            .I(N__5099));
    InMux I__722 (
            .O(N__5106),
            .I(N__5096));
    InMux I__721 (
            .O(N__5103),
            .I(N__5093));
    InMux I__720 (
            .O(N__5102),
            .I(N__5090));
    LocalMux I__719 (
            .O(N__5099),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__718 (
            .O(N__5096),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__717 (
            .O(N__5093),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__716 (
            .O(N__5090),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__715 (
            .O(N__5081),
            .I(\U712_CYCLE_TERM.N_351_cascade_ ));
    InMux I__714 (
            .O(N__5078),
            .I(N__5073));
    InMux I__713 (
            .O(N__5077),
            .I(N__5069));
    InMux I__712 (
            .O(N__5076),
            .I(N__5066));
    LocalMux I__711 (
            .O(N__5073),
            .I(N__5063));
    InMux I__710 (
            .O(N__5072),
            .I(N__5060));
    LocalMux I__709 (
            .O(N__5069),
            .I(N__5055));
    LocalMux I__708 (
            .O(N__5066),
            .I(N__5055));
    Span4Mux_v I__707 (
            .O(N__5063),
            .I(N__5050));
    LocalMux I__706 (
            .O(N__5060),
            .I(N__5050));
    Span4Mux_v I__705 (
            .O(N__5055),
            .I(N__5047));
    Span4Mux_h I__704 (
            .O(N__5050),
            .I(N__5044));
    Sp12to4 I__703 (
            .O(N__5047),
            .I(N__5041));
    Span4Mux_h I__702 (
            .O(N__5044),
            .I(N__5038));
    Span12Mux_h I__701 (
            .O(N__5041),
            .I(N__5033));
    Sp12to4 I__700 (
            .O(N__5038),
            .I(N__5033));
    Span12Mux_v I__699 (
            .O(N__5033),
            .I(N__5030));
    Odrv12 I__698 (
            .O(N__5030),
            .I(CLK40_PLL_i));
    InMux I__697 (
            .O(N__5027),
            .I(N__5024));
    LocalMux I__696 (
            .O(N__5024),
            .I(N__5020));
    InMux I__695 (
            .O(N__5023),
            .I(N__5017));
    Span4Mux_v I__694 (
            .O(N__5020),
            .I(N__5012));
    LocalMux I__693 (
            .O(N__5017),
            .I(N__5009));
    InMux I__692 (
            .O(N__5016),
            .I(N__5006));
    InMux I__691 (
            .O(N__5015),
            .I(N__5003));
    Odrv4 I__690 (
            .O(N__5012),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__689 (
            .O(N__5009),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__688 (
            .O(N__5006),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__687 (
            .O(N__5003),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__686 (
            .O(N__4994),
            .I(N__4990));
    InMux I__685 (
            .O(N__4993),
            .I(N__4987));
    LocalMux I__684 (
            .O(N__4990),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ));
    LocalMux I__683 (
            .O(N__4987),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ));
    InMux I__682 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__681 (
            .O(N__4979),
            .I(N__4976));
    Odrv4 I__680 (
            .O(N__4976),
            .I(\U712_CHIP_RAM.N_325 ));
    CascadeMux I__679 (
            .O(N__4973),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ));
    InMux I__678 (
            .O(N__4970),
            .I(N__4967));
    LocalMux I__677 (
            .O(N__4967),
            .I(N__4964));
    Odrv4 I__676 (
            .O(N__4964),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__675 (
            .O(N__4961),
            .I(N__4957));
    InMux I__674 (
            .O(N__4960),
            .I(N__4954));
    LocalMux I__673 (
            .O(N__4957),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__672 (
            .O(N__4954),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__671 (
            .O(N__4949),
            .I(N__4945));
    InMux I__670 (
            .O(N__4948),
            .I(N__4942));
    LocalMux I__669 (
            .O(N__4945),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__668 (
            .O(N__4942),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__667 (
            .O(N__4937),
            .I(N__4933));
    InMux I__666 (
            .O(N__4936),
            .I(N__4930));
    InMux I__665 (
            .O(N__4933),
            .I(N__4927));
    LocalMux I__664 (
            .O(N__4930),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__663 (
            .O(N__4927),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__662 (
            .O(N__4922),
            .I(N__4918));
    InMux I__661 (
            .O(N__4921),
            .I(N__4915));
    LocalMux I__660 (
            .O(N__4918),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__659 (
            .O(N__4915),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__658 (
            .O(N__4910),
            .I(\U712_CHIP_RAM.N_241_cascade_ ));
    CascadeMux I__657 (
            .O(N__4907),
            .I(\U712_CHIP_RAM.N_388_cascade_ ));
    InMux I__656 (
            .O(N__4904),
            .I(N__4900));
    InMux I__655 (
            .O(N__4903),
            .I(N__4897));
    LocalMux I__654 (
            .O(N__4900),
            .I(\U712_CHIP_RAM.N_325_1 ));
    LocalMux I__653 (
            .O(N__4897),
            .I(\U712_CHIP_RAM.N_325_1 ));
    CascadeMux I__652 (
            .O(N__4892),
            .I(N__4888));
    CascadeMux I__651 (
            .O(N__4891),
            .I(N__4884));
    InMux I__650 (
            .O(N__4888),
            .I(N__4879));
    InMux I__649 (
            .O(N__4887),
            .I(N__4875));
    InMux I__648 (
            .O(N__4884),
            .I(N__4872));
    InMux I__647 (
            .O(N__4883),
            .I(N__4867));
    InMux I__646 (
            .O(N__4882),
            .I(N__4867));
    LocalMux I__645 (
            .O(N__4879),
            .I(N__4864));
    InMux I__644 (
            .O(N__4878),
            .I(N__4861));
    LocalMux I__643 (
            .O(N__4875),
            .I(\U712_CHIP_RAM.N_381 ));
    LocalMux I__642 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.N_381 ));
    LocalMux I__641 (
            .O(N__4867),
            .I(\U712_CHIP_RAM.N_381 ));
    Odrv4 I__640 (
            .O(N__4864),
            .I(\U712_CHIP_RAM.N_381 ));
    LocalMux I__639 (
            .O(N__4861),
            .I(\U712_CHIP_RAM.N_381 ));
    InMux I__638 (
            .O(N__4850),
            .I(N__4844));
    InMux I__637 (
            .O(N__4849),
            .I(N__4844));
    LocalMux I__636 (
            .O(N__4844),
            .I(N__4841));
    Odrv4 I__635 (
            .O(N__4841),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    IoInMux I__634 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__633 (
            .O(N__4835),
            .I(N__4832));
    IoSpan4Mux I__632 (
            .O(N__4832),
            .I(N__4829));
    Span4Mux_s3_v I__631 (
            .O(N__4829),
            .I(N__4826));
    Span4Mux_v I__630 (
            .O(N__4826),
            .I(N__4823));
    Odrv4 I__629 (
            .O(N__4823),
            .I(N_249_i));
    InMux I__628 (
            .O(N__4820),
            .I(N__4817));
    LocalMux I__627 (
            .O(N__4817),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0 ));
    CascadeMux I__626 (
            .O(N__4814),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_ ));
    CascadeMux I__625 (
            .O(N__4811),
            .I(\U712_CHIP_RAM.N_325_cascade_ ));
    IoInMux I__624 (
            .O(N__4808),
            .I(N__4805));
    LocalMux I__623 (
            .O(N__4805),
            .I(N__4802));
    IoSpan4Mux I__622 (
            .O(N__4802),
            .I(N__4799));
    Span4Mux_s3_h I__621 (
            .O(N__4799),
            .I(N__4795));
    InMux I__620 (
            .O(N__4798),
            .I(N__4792));
    Span4Mux_h I__619 (
            .O(N__4795),
            .I(N__4789));
    LocalMux I__618 (
            .O(N__4792),
            .I(N__4786));
    Sp12to4 I__617 (
            .O(N__4789),
            .I(N__4783));
    Span4Mux_v I__616 (
            .O(N__4786),
            .I(N__4780));
    Span12Mux_h I__615 (
            .O(N__4783),
            .I(N__4775));
    Sp12to4 I__614 (
            .O(N__4780),
            .I(N__4775));
    Span12Mux_h I__613 (
            .O(N__4775),
            .I(N__4772));
    Span12Mux_v I__612 (
            .O(N__4772),
            .I(N__4769));
    Odrv12 I__611 (
            .O(N__4769),
            .I(C3_c));
    InMux I__610 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__609 (
            .O(N__4763),
            .I(N__4759));
    InMux I__608 (
            .O(N__4762),
            .I(N__4756));
    Span4Mux_h I__607 (
            .O(N__4759),
            .I(N__4751));
    LocalMux I__606 (
            .O(N__4756),
            .I(N__4751));
    Span4Mux_v I__605 (
            .O(N__4751),
            .I(N__4748));
    Span4Mux_h I__604 (
            .O(N__4748),
            .I(N__4745));
    Sp12to4 I__603 (
            .O(N__4745),
            .I(N__4742));
    Span12Mux_v I__602 (
            .O(N__4742),
            .I(N__4739));
    Odrv12 I__601 (
            .O(N__4739),
            .I(DBRn_c));
    InMux I__600 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__599 (
            .O(N__4733),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    InMux I__598 (
            .O(N__4730),
            .I(N__4727));
    LocalMux I__597 (
            .O(N__4727),
            .I(N__4724));
    Span4Mux_h I__596 (
            .O(N__4724),
            .I(N__4721));
    Sp12to4 I__595 (
            .O(N__4721),
            .I(N__4718));
    Span12Mux_v I__594 (
            .O(N__4718),
            .I(N__4715));
    Odrv12 I__593 (
            .O(N__4715),
            .I(A_c_20));
    InMux I__592 (
            .O(N__4712),
            .I(N__4709));
    LocalMux I__591 (
            .O(N__4709),
            .I(N__4706));
    Span4Mux_v I__590 (
            .O(N__4706),
            .I(N__4703));
    Odrv4 I__589 (
            .O(N__4703),
            .I(\U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0 ));
    InMux I__588 (
            .O(N__4700),
            .I(N__4696));
    InMux I__587 (
            .O(N__4699),
            .I(N__4693));
    LocalMux I__586 (
            .O(N__4696),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__585 (
            .O(N__4693),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__584 (
            .O(N__4688),
            .I(N__4685));
    InMux I__583 (
            .O(N__4685),
            .I(N__4681));
    InMux I__582 (
            .O(N__4684),
            .I(N__4678));
    LocalMux I__581 (
            .O(N__4681),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__580 (
            .O(N__4678),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__579 (
            .O(N__4673),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    CascadeMux I__578 (
            .O(N__4670),
            .I(\U712_CYCLE_TERM.N_269_i_0_en_cascade_ ));
    CEMux I__577 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__576 (
            .O(N__4664),
            .I(N__4661));
    Odrv4 I__575 (
            .O(N__4661),
            .I(\U712_CYCLE_TERM.N_269_i_0_en_0 ));
    CascadeMux I__574 (
            .O(N__4658),
            .I(\U712_CHIP_RAM.N_76_cascade_ ));
    InMux I__573 (
            .O(N__4655),
            .I(N__4651));
    InMux I__572 (
            .O(N__4654),
            .I(N__4648));
    LocalMux I__571 (
            .O(N__4651),
            .I(\U712_CHIP_RAM.N_328 ));
    LocalMux I__570 (
            .O(N__4648),
            .I(\U712_CHIP_RAM.N_328 ));
    IoInMux I__569 (
            .O(N__4643),
            .I(N__4640));
    LocalMux I__568 (
            .O(N__4640),
            .I(N__4637));
    Span4Mux_s3_v I__567 (
            .O(N__4637),
            .I(N__4634));
    Sp12to4 I__566 (
            .O(N__4634),
            .I(N__4631));
    Span12Mux_s11_h I__565 (
            .O(N__4631),
            .I(N__4628));
    Span12Mux_v I__564 (
            .O(N__4628),
            .I(N__4624));
    InMux I__563 (
            .O(N__4627),
            .I(N__4621));
    Odrv12 I__562 (
            .O(N__4624),
            .I(LATCH_CLK_c));
    LocalMux I__561 (
            .O(N__4621),
            .I(LATCH_CLK_c));
    CascadeMux I__560 (
            .O(N__4616),
            .I(\U712_CHIP_RAM.N_438_cascade_ ));
    InMux I__559 (
            .O(N__4613),
            .I(N__4607));
    InMux I__558 (
            .O(N__4612),
            .I(N__4607));
    LocalMux I__557 (
            .O(N__4607),
            .I(\U712_CHIP_RAM.N_336 ));
    CascadeMux I__556 (
            .O(N__4604),
            .I(N__4600));
    CascadeMux I__555 (
            .O(N__4603),
            .I(N__4595));
    InMux I__554 (
            .O(N__4600),
            .I(N__4592));
    InMux I__553 (
            .O(N__4599),
            .I(N__4589));
    InMux I__552 (
            .O(N__4598),
            .I(N__4585));
    InMux I__551 (
            .O(N__4595),
            .I(N__4582));
    LocalMux I__550 (
            .O(N__4592),
            .I(N__4577));
    LocalMux I__549 (
            .O(N__4589),
            .I(N__4577));
    InMux I__548 (
            .O(N__4588),
            .I(N__4574));
    LocalMux I__547 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__546 (
            .O(N__4582),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__545 (
            .O(N__4577),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__544 (
            .O(N__4574),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    InMux I__543 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__542 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_h I__541 (
            .O(N__4559),
            .I(N__4556));
    Odrv4 I__540 (
            .O(N__4556),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    CascadeMux I__539 (
            .O(N__4553),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ));
    InMux I__538 (
            .O(N__4550),
            .I(N__4546));
    InMux I__537 (
            .O(N__4549),
            .I(N__4543));
    LocalMux I__536 (
            .O(N__4546),
            .I(\U712_CHIP_RAM.N_438 ));
    LocalMux I__535 (
            .O(N__4543),
            .I(\U712_CHIP_RAM.N_438 ));
    InMux I__534 (
            .O(N__4538),
            .I(N__4535));
    LocalMux I__533 (
            .O(N__4535),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0 ));
    InMux I__532 (
            .O(N__4532),
            .I(N__4529));
    LocalMux I__531 (
            .O(N__4529),
            .I(\U712_CHIP_RAM.N_247 ));
    CascadeMux I__530 (
            .O(N__4526),
            .I(\U712_CHIP_RAM.N_247_cascade_ ));
    InMux I__529 (
            .O(N__4523),
            .I(N__4520));
    LocalMux I__528 (
            .O(N__4520),
            .I(N__4517));
    Span4Mux_h I__527 (
            .O(N__4517),
            .I(N__4513));
    InMux I__526 (
            .O(N__4516),
            .I(N__4510));
    Odrv4 I__525 (
            .O(N__4513),
            .I(\U712_CHIP_RAM.N_244 ));
    LocalMux I__524 (
            .O(N__4510),
            .I(\U712_CHIP_RAM.N_244 ));
    InMux I__523 (
            .O(N__4505),
            .I(N__4502));
    LocalMux I__522 (
            .O(N__4502),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0 ));
    InMux I__521 (
            .O(N__4499),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__520 (
            .O(N__4496),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__519 (
            .O(N__4493),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__518 (
            .O(N__4490),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__517 (
            .O(N__4487),
            .I(N__4474));
    InMux I__516 (
            .O(N__4486),
            .I(N__4474));
    InMux I__515 (
            .O(N__4485),
            .I(N__4474));
    InMux I__514 (
            .O(N__4484),
            .I(N__4471));
    InMux I__513 (
            .O(N__4483),
            .I(N__4464));
    InMux I__512 (
            .O(N__4482),
            .I(N__4464));
    InMux I__511 (
            .O(N__4481),
            .I(N__4464));
    LocalMux I__510 (
            .O(N__4474),
            .I(\U712_CHIP_RAM.N_236 ));
    LocalMux I__509 (
            .O(N__4471),
            .I(\U712_CHIP_RAM.N_236 ));
    LocalMux I__508 (
            .O(N__4464),
            .I(\U712_CHIP_RAM.N_236 ));
    InMux I__507 (
            .O(N__4457),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__506 (
            .O(N__4454),
            .I(N__4451));
    LocalMux I__505 (
            .O(N__4451),
            .I(N__4447));
    CEMux I__504 (
            .O(N__4450),
            .I(N__4444));
    Span4Mux_v I__503 (
            .O(N__4447),
            .I(N__4441));
    LocalMux I__502 (
            .O(N__4444),
            .I(N__4438));
    Span4Mux_h I__501 (
            .O(N__4441),
            .I(N__4435));
    Span4Mux_h I__500 (
            .O(N__4438),
            .I(N__4432));
    Odrv4 I__499 (
            .O(N__4435),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__498 (
            .O(N__4432),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__497 (
            .O(N__4427),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_ ));
    InMux I__496 (
            .O(N__4424),
            .I(N__4421));
    LocalMux I__495 (
            .O(N__4421),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1 ));
    InMux I__494 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__493 (
            .O(N__4415),
            .I(\U712_CHIP_RAM.N_348 ));
    InMux I__492 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__491 (
            .O(N__4409),
            .I(N__4405));
    InMux I__490 (
            .O(N__4408),
            .I(N__4402));
    Odrv4 I__489 (
            .O(N__4405),
            .I(\U712_CHIP_RAM.N_437 ));
    LocalMux I__488 (
            .O(N__4402),
            .I(\U712_CHIP_RAM.N_437 ));
    CascadeMux I__487 (
            .O(N__4397),
            .I(N__4393));
    InMux I__486 (
            .O(N__4396),
            .I(N__4388));
    InMux I__485 (
            .O(N__4393),
            .I(N__4385));
    InMux I__484 (
            .O(N__4392),
            .I(N__4382));
    InMux I__483 (
            .O(N__4391),
            .I(N__4379));
    LocalMux I__482 (
            .O(N__4388),
            .I(\U712_CHIP_RAM.N_426 ));
    LocalMux I__481 (
            .O(N__4385),
            .I(\U712_CHIP_RAM.N_426 ));
    LocalMux I__480 (
            .O(N__4382),
            .I(\U712_CHIP_RAM.N_426 ));
    LocalMux I__479 (
            .O(N__4379),
            .I(\U712_CHIP_RAM.N_426 ));
    CascadeMux I__478 (
            .O(N__4370),
            .I(\U712_CHIP_RAM.N_300_cascade_ ));
    InMux I__477 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__476 (
            .O(N__4364),
            .I(\U712_CHIP_RAM.N_301 ));
    InMux I__475 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__474 (
            .O(N__4358),
            .I(\U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431 ));
    InMux I__473 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__472 (
            .O(N__4352),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1 ));
    InMux I__471 (
            .O(N__4349),
            .I(N__4346));
    LocalMux I__470 (
            .O(N__4346),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ));
    InMux I__469 (
            .O(N__4343),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__468 (
            .O(N__4340),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__467 (
            .O(N__4337),
            .I(N__4334));
    InMux I__466 (
            .O(N__4334),
            .I(N__4329));
    InMux I__465 (
            .O(N__4333),
            .I(N__4324));
    InMux I__464 (
            .O(N__4332),
            .I(N__4324));
    LocalMux I__463 (
            .O(N__4329),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__462 (
            .O(N__4324),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__461 (
            .O(N__4319),
            .I(N__4316));
    InMux I__460 (
            .O(N__4316),
            .I(N__4310));
    InMux I__459 (
            .O(N__4315),
            .I(N__4310));
    LocalMux I__458 (
            .O(N__4310),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__457 (
            .O(N__4307),
            .I(N__4304));
    LocalMux I__456 (
            .O(N__4304),
            .I(N__4301));
    Span4Mux_v I__455 (
            .O(N__4301),
            .I(N__4298));
    Odrv4 I__454 (
            .O(N__4298),
            .I(TACK_EN_i_ess));
    IoInMux I__453 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__452 (
            .O(N__4292),
            .I(N__4289));
    Odrv12 I__451 (
            .O(N__4289),
            .I(VBENn_c));
    CascadeMux I__450 (
            .O(N__4286),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_ ));
    CascadeMux I__449 (
            .O(N__4283),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_ ));
    CEMux I__448 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__447 (
            .O(N__4277),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0 ));
    InMux I__446 (
            .O(N__4274),
            .I(N__4271));
    LocalMux I__445 (
            .O(N__4271),
            .I(N__4268));
    Odrv4 I__444 (
            .O(N__4268),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0 ));
    CascadeMux I__443 (
            .O(N__4265),
            .I(\U712_CHIP_RAM.N_350_cascade_ ));
    CascadeMux I__442 (
            .O(N__4262),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ));
    CEMux I__441 (
            .O(N__4259),
            .I(N__4256));
    LocalMux I__440 (
            .O(N__4256),
            .I(N__4253));
    Span4Mux_h I__439 (
            .O(N__4253),
            .I(N__4250));
    Odrv4 I__438 (
            .O(N__4250),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ));
    InMux I__437 (
            .O(N__4247),
            .I(N__4244));
    LocalMux I__436 (
            .O(N__4244),
            .I(\U712_CHIP_RAM.N_350 ));
    InMux I__435 (
            .O(N__4241),
            .I(N__4237));
    InMux I__434 (
            .O(N__4240),
            .I(N__4234));
    LocalMux I__433 (
            .O(N__4237),
            .I(N__4231));
    LocalMux I__432 (
            .O(N__4234),
            .I(N__4228));
    Span4Mux_h I__431 (
            .O(N__4231),
            .I(N__4223));
    Span4Mux_v I__430 (
            .O(N__4228),
            .I(N__4223));
    Sp12to4 I__429 (
            .O(N__4223),
            .I(N__4220));
    Span12Mux_h I__428 (
            .O(N__4220),
            .I(N__4217));
    Span12Mux_v I__427 (
            .O(N__4217),
            .I(N__4214));
    Odrv12 I__426 (
            .O(N__4214),
            .I(AWEn_c));
    InMux I__425 (
            .O(N__4211),
            .I(N__4208));
    LocalMux I__424 (
            .O(N__4208),
            .I(\U712_CHIP_RAM.N_287 ));
    InMux I__423 (
            .O(N__4205),
            .I(N__4202));
    LocalMux I__422 (
            .O(N__4202),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__421 (
            .O(N__4199),
            .I(N__4196));
    LocalMux I__420 (
            .O(N__4196),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__419 (
            .O(N__4193),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_ ));
    CascadeMux I__418 (
            .O(N__4190),
            .I(\U712_CHIP_RAM.N_265_cascade_ ));
    InMux I__417 (
            .O(N__4187),
            .I(N__4184));
    LocalMux I__416 (
            .O(N__4184),
            .I(\U712_CHIP_RAM.N_265 ));
    CascadeMux I__415 (
            .O(N__4181),
            .I(\U712_CHIP_RAM.N_236_cascade_ ));
    CascadeMux I__414 (
            .O(N__4178),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    CascadeMux I__413 (
            .O(N__4175),
            .I(\U712_CHIP_RAM.N_426_cascade_ ));
    IoInMux I__412 (
            .O(N__4172),
            .I(N__4169));
    LocalMux I__411 (
            .O(N__4169),
            .I(N__4166));
    IoSpan4Mux I__410 (
            .O(N__4166),
            .I(N__4163));
    Span4Mux_s3_v I__409 (
            .O(N__4163),
            .I(N__4160));
    Span4Mux_v I__408 (
            .O(N__4160),
            .I(N__4157));
    Span4Mux_v I__407 (
            .O(N__4157),
            .I(N__4154));
    Odrv4 I__406 (
            .O(N__4154),
            .I(BANK0_c));
    InMux I__405 (
            .O(N__4151),
            .I(N__4148));
    LocalMux I__404 (
            .O(N__4148),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ));
    CascadeMux I__403 (
            .O(N__4145),
            .I(\U712_CHIP_RAM.N_186_cascade_ ));
    IoInMux I__402 (
            .O(N__4142),
            .I(N__4139));
    LocalMux I__401 (
            .O(N__4139),
            .I(N__4136));
    Span4Mux_s3_v I__400 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_v I__399 (
            .O(N__4133),
            .I(N__4129));
    InMux I__398 (
            .O(N__4132),
            .I(N__4126));
    Odrv4 I__397 (
            .O(N__4129),
            .I(DBDIR_c));
    LocalMux I__396 (
            .O(N__4126),
            .I(DBDIR_c));
    IoInMux I__395 (
            .O(N__4121),
            .I(N__4118));
    LocalMux I__394 (
            .O(N__4118),
            .I(N__4115));
    Span4Mux_s2_h I__393 (
            .O(N__4115),
            .I(N__4112));
    Sp12to4 I__392 (
            .O(N__4112),
            .I(N__4109));
    Span12Mux_v I__391 (
            .O(N__4109),
            .I(N__4105));
    InMux I__390 (
            .O(N__4108),
            .I(N__4102));
    Odrv12 I__389 (
            .O(N__4105),
            .I(TACK_OUTn));
    LocalMux I__388 (
            .O(N__4102),
            .I(TACK_OUTn));
    IoInMux I__387 (
            .O(N__4097),
            .I(N__4094));
    LocalMux I__386 (
            .O(N__4094),
            .I(N__4090));
    IoInMux I__385 (
            .O(N__4093),
            .I(N__4087));
    IoSpan4Mux I__384 (
            .O(N__4090),
            .I(N__4082));
    LocalMux I__383 (
            .O(N__4087),
            .I(N__4082));
    IoSpan4Mux I__382 (
            .O(N__4082),
            .I(N__4078));
    IoInMux I__381 (
            .O(N__4081),
            .I(N__4075));
    IoSpan4Mux I__380 (
            .O(N__4078),
            .I(N__4072));
    LocalMux I__379 (
            .O(N__4075),
            .I(N__4069));
    Sp12to4 I__378 (
            .O(N__4072),
            .I(N__4066));
    IoSpan4Mux I__377 (
            .O(N__4069),
            .I(N__4063));
    Span12Mux_s6_v I__376 (
            .O(N__4066),
            .I(N__4060));
    Span4Mux_s2_h I__375 (
            .O(N__4063),
            .I(N__4057));
    Span12Mux_h I__374 (
            .O(N__4060),
            .I(N__4054));
    Span4Mux_h I__373 (
            .O(N__4057),
            .I(N__4051));
    Odrv12 I__372 (
            .O(N__4054),
            .I(CLK40_PLL_i_i));
    Odrv4 I__371 (
            .O(N__4051),
            .I(CLK40_PLL_i_i));
    CascadeMux I__370 (
            .O(N__4046),
            .I(N__4043));
    InMux I__369 (
            .O(N__4043),
            .I(N__4040));
    LocalMux I__368 (
            .O(N__4040),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0 ));
    IoInMux I__367 (
            .O(N__4037),
            .I(N__4034));
    LocalMux I__366 (
            .O(N__4034),
            .I(N__4031));
    IoSpan4Mux I__365 (
            .O(N__4031),
            .I(N__4028));
    Span4Mux_s3_h I__364 (
            .O(N__4028),
            .I(N__4025));
    Odrv4 I__363 (
            .O(N__4025),
            .I(DBRn_c_i_0));
    IoInMux I__362 (
            .O(N__4022),
            .I(N__4019));
    LocalMux I__361 (
            .O(N__4019),
            .I(N__4016));
    Span4Mux_s2_h I__360 (
            .O(N__4016),
            .I(N__4013));
    Span4Mux_h I__359 (
            .O(N__4013),
            .I(N__4010));
    Span4Mux_v I__358 (
            .O(N__4010),
            .I(N__4007));
    Odrv4 I__357 (
            .O(N__4007),
            .I(N_996_i));
    IoInMux I__356 (
            .O(N__4004),
            .I(N__4001));
    LocalMux I__355 (
            .O(N__4001),
            .I(N__3998));
    Span4Mux_s2_v I__354 (
            .O(N__3998),
            .I(N__3995));
    Span4Mux_v I__353 (
            .O(N__3995),
            .I(N__3992));
    Span4Mux_h I__352 (
            .O(N__3992),
            .I(N__3989));
    Odrv4 I__351 (
            .O(N__3989),
            .I(CLK80_PLL_i_i));
    IoInMux I__350 (
            .O(N__3986),
            .I(N__3983));
    LocalMux I__349 (
            .O(N__3983),
            .I(N__3980));
    Span4Mux_s0_v I__348 (
            .O(N__3980),
            .I(N__3977));
    Span4Mux_v I__347 (
            .O(N__3977),
            .I(N__3974));
    Sp12to4 I__346 (
            .O(N__3974),
            .I(N__3971));
    Span12Mux_h I__345 (
            .O(N__3971),
            .I(N__3968));
    Span12Mux_v I__344 (
            .O(N__3968),
            .I(N__3965));
    Odrv12 I__343 (
            .O(N__3965),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__7693));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__7695));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__7690));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__7692));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__7687));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__7688));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__7689));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__7691));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7349),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5560),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4037),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4808),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__10997),
            .in2(_gnd_net_),
            .in3(N__7999),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_3_14_2.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_3_14_2.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_3_14_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_3_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4307),
            .lcout(N_996_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_10_7.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4762),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_6_1_7.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_6_1_7.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_6_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_6_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8696),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_6_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_6_6_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_6_6_0 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_6_6_0  (
            .in0(N__5472),
            .in1(N__4151),
            .in2(N__4603),
            .in3(N__10316),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8679),
            .ce(),
            .sr(N__10976));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNICLGI4_LC_6_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNICLGI4_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNICLGI4_LC_6_6_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNICLGI4_LC_6_6_2  (
            .in0(N__4391),
            .in1(N__6367),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_6_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_6_6_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_6_6_3 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_6_6_3  (
            .in0(N__4240),
            .in1(_gnd_net_),
            .in2(N__4145),
            .in3(N__4132),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8679),
            .ce(),
            .sr(N__10976));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_6_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_6_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__6161),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_6_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_6_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__4396),
            .in2(_gnd_net_),
            .in3(N__6363),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8684),
            .ce(N__4280),
            .sr(N__10972));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_6_8_3 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_6_8_3  (
            .in0(N__4108),
            .in1(N__5076),
            .in2(N__4337),
            .in3(N__5023),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8688),
            .ce(),
            .sr(N__10967));
    defparam pll_RNI8MQ3_LC_6_9_3.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_6_9_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_6_9_3 (
            .in0(N__5077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_5_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_5_2  (
            .in0(N__4349),
            .in1(N__4484),
            .in2(N__4046),
            .in3(N__4598),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8672),
            .ce(N__4450),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5012_1_LC_7_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5012_1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5012_1_LC_7_5_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5012_1_LC_7_5_3  (
            .in0(N__4361),
            .in1(N__6723),
            .in2(_gnd_net_),
            .in3(N__5902),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINE0O4_LC_7_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINE0O4_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINE0O4_LC_7_5_4 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINE0O4_LC_7_5_4  (
            .in0(N__7533),
            .in1(N__6368),
            .in2(N__4193),
            .in3(N__6470),
            .lcout(\U712_CHIP_RAM.N_265 ),
            .ltout(\U712_CHIP_RAM.N_265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMBRQ8_3_LC_7_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMBRQ8_3_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMBRQ8_3_LC_7_5_5 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMBRQ8_3_LC_7_5_5  (
            .in0(N__4367),
            .in1(_gnd_net_),
            .in2(N__4190),
            .in3(N__4887),
            .lcout(\U712_CHIP_RAM.N_236 ),
            .ltout(\U712_CHIP_RAM.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_5_6 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_5_6  (
            .in0(N__4970),
            .in1(N__4187),
            .in2(N__4181),
            .in3(N__5228),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8672),
            .ce(N__4450),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_7_6_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_7_6_0  (
            .in0(N__6551),
            .in1(N__5903),
            .in2(N__4892),
            .in3(N__6724),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_7_6_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__6078),
            .in2(N__4178),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_426 ),
            .ltout(\U712_CHIP_RAM.N_426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIQ2RS7_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIQ2RS7_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIQ2RS7_LC_7_6_2 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIQ2RS7_LC_7_6_2  (
            .in0(N__5431),
            .in1(N__6366),
            .in2(N__4175),
            .in3(N__4408),
            .lcout(\U712_CHIP_RAM.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_LC_7_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_7_6_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_LC_7_6_5  (
            .in0(N__4565),
            .in1(N__4712),
            .in2(N__4397),
            .in3(N__7982),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8675),
            .ce(N__4259),
            .sr(N__10973));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_0 .LUT_INIT=16'b1011100011111000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_0  (
            .in0(N__4205),
            .in1(N__7515),
            .in2(N__6092),
            .in3(N__5435),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIIE53C_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIIE53C_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIIE53C_LC_7_7_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIIE53C_LC_7_7_1  (
            .in0(N__4505),
            .in1(N__4549),
            .in2(_gnd_net_),
            .in3(N__4654),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2  (
            .in0(N__7339),
            .in1(_gnd_net_),
            .in2(N__4283),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ6QH5_LC_7_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ6QH5_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ6QH5_LC_7_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ6QH5_LC_7_7_3  (
            .in0(N__6361),
            .in1(N__4588),
            .in2(_gnd_net_),
            .in3(N__4516),
            .lcout(\U712_CHIP_RAM.N_350 ),
            .ltout(\U712_CHIP_RAM.N_350_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_7_7_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_7_7_4  (
            .in0(N__4274),
            .in1(N__6362),
            .in2(N__4265),
            .in3(N__6469),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_7_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_7_5  (
            .in0(N__10996),
            .in1(_gnd_net_),
            .in2(N__4262),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_7_6 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_7_7_6  (
            .in0(N__4211),
            .in1(N__7516),
            .in2(N__6882),
            .in3(N__4247),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_7_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_7_7  (
            .in0(N__4241),
            .in1(N__6935),
            .in2(_gnd_net_),
            .in3(N__6079),
            .lcout(\U712_CHIP_RAM.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_7_8_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_7_8_0  (
            .in0(N__6761),
            .in1(N__9321),
            .in2(N__6619),
            .in3(N__6848),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_8_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__4199),
            .in2(_gnd_net_),
            .in3(N__4849),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_4  (
            .in0(N__4850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7532),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8685),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__7531),
            .in2(_gnd_net_),
            .in3(N__4333),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8689),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_1  (
            .in0(N__7529),
            .in1(N__5072),
            .in2(_gnd_net_),
            .in3(N__5027),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8689),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_3  (
            .in0(N__7530),
            .in1(_gnd_net_),
            .in2(N__4319),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8689),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__4332),
            .in2(_gnd_net_),
            .in3(N__4315),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_3  (
            .in0(N__7528),
            .in1(N__4700),
            .in2(_gnd_net_),
            .in3(N__5107),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8691),
            .ce(N__4667),
            .sr(N__10949));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_3_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_3_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_3_3  (
            .in0(N__10843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9385),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_4_0 .LUT_INIT=16'b0000111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_4_0  (
            .in0(N__6764),
            .in1(N__5817),
            .in2(N__6620),
            .in3(N__6364),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_4_1 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_4_1  (
            .in0(N__6460),
            .in1(_gnd_net_),
            .in2(N__4286),
            .in3(N__7527),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_4_5 .LUT_INIT=16'b1111100011101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_4_5  (
            .in0(N__5818),
            .in1(N__6765),
            .in2(N__5954),
            .in3(N__6608),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_5_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_5_0  (
            .in0(N__6435),
            .in1(N__4355),
            .in2(_gnd_net_),
            .in3(N__6155),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_5_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_5_1  (
            .in0(N__6359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5896),
            .lcout(\U712_CHIP_RAM.N_300 ),
            .ltout(\U712_CHIP_RAM.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_5_2 .LUT_INIT=16'b1111111110100101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_5_2  (
            .in0(N__6720),
            .in1(_gnd_net_),
            .in2(N__4370),
            .in3(N__6548),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_8_5_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_8_5_4  (
            .in0(N__6095),
            .in1(N__6132),
            .in2(N__4604),
            .in3(N__4904),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_8_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_8_5_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_8_5_5  (
            .in0(N__5798),
            .in1(N__5895),
            .in2(N__6468),
            .in3(N__6719),
            .lcout(\U712_CHIP_RAM.N_437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIUL431_LC_8_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIUL431_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIUL431_LC_8_5_6 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIUL431_LC_8_5_6  (
            .in0(N__5448),
            .in1(N__6544),
            .in2(N__6891),
            .in3(N__5796),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_5_7 .LUT_INIT=16'b0010100011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_5_7  (
            .in0(N__5797),
            .in1(N__6718),
            .in2(N__6592),
            .in3(N__5894),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__5799),
            .in2(_gnd_net_),
            .in3(N__6425),
            .lcout(\U712_CHIP_RAM.N_381 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_1_LC_8_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_1_LC_8_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__5930),
            .in2(_gnd_net_),
            .in3(N__4343),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_2  (
            .in0(N__4485),
            .in1(N__6585),
            .in2(_gnd_net_),
            .in3(N__4340),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_6_3  (
            .in0(N__4481),
            .in1(N__6754),
            .in2(_gnd_net_),
            .in3(N__4499),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_4  (
            .in0(N__4486),
            .in1(N__4922),
            .in2(_gnd_net_),
            .in3(N__4496),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_5  (
            .in0(N__4482),
            .in1(N__4949),
            .in2(_gnd_net_),
            .in3(N__4493),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_6  (
            .in0(N__4487),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__4490),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_7  (
            .in0(N__4483),
            .in1(N__4936),
            .in2(_gnd_net_),
            .in3(N__4457),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8673),
            .ce(N__4454),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_0 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_0  (
            .in0(N__5156),
            .in1(N__4418),
            .in2(N__6467),
            .in3(N__5838),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_7_1  (
            .in0(N__5201),
            .in1(N__5128),
            .in2(N__4427),
            .in3(N__4612),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8676),
            .ce(),
            .sr(N__10963));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2  (
            .in0(N__5953),
            .in1(N__4424),
            .in2(_gnd_net_),
            .in3(N__4883),
            .lcout(\U712_CHIP_RAM.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_7_3 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_7_3  (
            .in0(N__5442),
            .in1(N__4412),
            .in2(_gnd_net_),
            .in3(N__4392),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_76_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_8_7_4 .LUT_INIT=16'b0000111101001110;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_8_7_4  (
            .in0(N__4613),
            .in1(N__4627),
            .in2(N__4658),
            .in3(N__4655),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8676),
            .ce(),
            .sr(N__10963));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_8_7_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_8_7_6  (
            .in0(N__5952),
            .in1(N__6360),
            .in2(_gnd_net_),
            .in3(N__4882),
            .lcout(\U712_CHIP_RAM.N_438 ),
            .ltout(\U712_CHIP_RAM.N_438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_7_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_7_7  (
            .in0(N__6609),
            .in1(N__6857),
            .in2(N__4616),
            .in3(N__6753),
            .lcout(\U712_CHIP_RAM.N_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_8_8_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_8_8_0  (
            .in0(N__6069),
            .in1(N__4599),
            .in2(N__6128),
            .in3(N__4532),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_1 .LUT_INIT=16'b1111010011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_1  (
            .in0(N__4538),
            .in1(N__9341),
            .in2(N__4553),
            .in3(N__4550),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8681),
            .ce(),
            .sr(N__10955));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_3  (
            .in0(N__6763),
            .in1(N__6600),
            .in2(_gnd_net_),
            .in3(N__6847),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_8_8_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__5145),
            .in2(_gnd_net_),
            .in3(N__5325),
            .lcout(\U712_CHIP_RAM.N_247 ),
            .ltout(\U712_CHIP_RAM.N_247_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_8_5 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__6115),
            .in2(N__4526),
            .in3(N__6068),
            .lcout(\U712_CHIP_RAM.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOVA11_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOVA11_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOVA11_LC_8_8_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIOVA11_LC_8_8_6  (
            .in0(N__6846),
            .in1(N__6762),
            .in2(_gnd_net_),
            .in3(N__6596),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_1_LC_8_8_7.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_8_8_7.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_8_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_8_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5345),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8681),
            .ce(),
            .sr(N__10955));
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_9_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5264),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8686),
            .ce(),
            .sr(N__10950));
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_9_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_8_9_1  (
            .in0(N__4798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8686),
            .ce(),
            .sr(N__10950));
    defparam DBR_SYNC_0_LC_8_9_2.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_8_9_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_8_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4766),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8686),
            .ce(),
            .sr(N__10950));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_9_4 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_9_4  (
            .in0(N__5016),
            .in1(N__4699),
            .in2(N__4688),
            .in3(N__4736),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8686),
            .ce(),
            .sr(N__10950));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__9965),
            .in2(_gnd_net_),
            .in3(N__4730),
            .lcout(\U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_8_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__5580),
            .in2(_gnd_net_),
            .in3(N__5129),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_10_4 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_10_4  (
            .in0(N__7476),
            .in1(N__4684),
            .in2(N__4673),
            .in3(N__5102),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_269_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_10_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_10_5  (
            .in0(N__10994),
            .in1(_gnd_net_),
            .in2(N__4670),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_269_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_11_3 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_8_11_3  (
            .in0(N__10776),
            .in1(N__7383),
            .in2(_gnd_net_),
            .in3(N__10715),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8692),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_0_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_0_LC_8_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_0_LC_8_12_3  (
            .in0(N__5496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5455),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_249_i_LC_8_19_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_249_i_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_249_i_LC_8_19_3 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.N_249_i_LC_8_19_3  (
            .in0(N__10787),
            .in1(N__10701),
            .in2(_gnd_net_),
            .in3(N__6892),
            .lcout(N_249_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_4_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_4_0  (
            .in0(N__6365),
            .in1(N__6773),
            .in2(_gnd_net_),
            .in3(N__5843),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_4_1 .LUT_INIT=16'b1111101010111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_4_1  (
            .in0(N__4820),
            .in1(N__6884),
            .in2(N__4814),
            .in3(N__5960),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8665),
            .ce(N__5650),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIIPOI5_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIIPOI5_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIIPOI5_LC_9_5_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIIPOI5_LC_9_5_0  (
            .in0(N__6093),
            .in1(N__4903),
            .in2(N__6134),
            .in3(N__6013),
            .lcout(\U712_CHIP_RAM.N_325 ),
            .ltout(\U712_CHIP_RAM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI0N6TH_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI0N6TH_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI0N6TH_LC_9_5_1 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI0N6TH_LC_9_5_1  (
            .in0(N__7522),
            .in1(N__4993),
            .in2(N__4811),
            .in3(N__5221),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_5_2 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_5_2  (
            .in0(N__6736),
            .in1(N__7526),
            .in2(N__6601),
            .in3(N__5937),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_5_3 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_5_3  (
            .in0(N__5938),
            .in1(N__5822),
            .in2(N__6602),
            .in3(N__6737),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_4  (
            .in0(N__6567),
            .in1(N__5939),
            .in2(N__4891),
            .in3(N__6157),
            .lcout(\U712_CHIP_RAM.N_317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_5 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_5  (
            .in0(N__4994),
            .in1(N__5220),
            .in2(N__7535),
            .in3(N__4982),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_6 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_6  (
            .in0(N__6002),
            .in1(_gnd_net_),
            .in2(N__4973),
            .in3(N__9034),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8669),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_7  (
            .in0(N__5722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5823),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_6_0  (
            .in0(N__4960),
            .in1(N__4948),
            .in2(N__4937),
            .in3(N__4921),
            .lcout(\U712_CHIP_RAM.N_241 ),
            .ltout(\U712_CHIP_RAM.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4GV43_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4GV43_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4GV43_LC_9_6_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4GV43_LC_9_6_1  (
            .in0(N__6721),
            .in1(N__6549),
            .in2(N__4910),
            .in3(N__6310),
            .lcout(\U712_CHIP_RAM.N_386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__7521),
            .in2(_gnd_net_),
            .in3(N__6293),
            .lcout(\U712_CHIP_RAM.N_388 ),
            .ltout(\U712_CHIP_RAM.N_388_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_9_6_3 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__5150),
            .in2(N__4907),
            .in3(N__5332),
            .lcout(\U712_CHIP_RAM.N_325_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_9_6_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_9_6_4  (
            .in0(N__6550),
            .in1(N__6722),
            .in2(_gnd_net_),
            .in3(N__4878),
            .lcout(\U712_CHIP_RAM.N_434 ),
            .ltout(\U712_CHIP_RAM.N_434_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3DQ77_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3DQ77_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3DQ77_LC_9_6_5 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3DQ77_LC_9_6_5  (
            .in0(N__5955),
            .in1(N__5237),
            .in2(N__5231),
            .in3(N__6311),
            .lcout(\U712_CHIP_RAM.N_439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_6_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_6_6  (
            .in0(N__5207),
            .in1(N__6294),
            .in2(_gnd_net_),
            .in3(N__6443),
            .lcout(\U712_CHIP_RAM.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_7  (
            .in0(N__5195),
            .in1(N__5177),
            .in2(_gnd_net_),
            .in3(N__9054),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_9_7_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__9339),
            .in2(_gnd_net_),
            .in3(N__6867),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_2  (
            .in0(N__6752),
            .in1(N__6584),
            .in2(N__5159),
            .in3(N__5958),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_3 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_3  (
            .in0(N__5354),
            .in1(N__9340),
            .in2(N__7534),
            .in3(N__5149),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8674),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_8_1 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_8_1  (
            .in0(N__7193),
            .in1(N__7604),
            .in2(N__7520),
            .in3(N__7544),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8677),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_8_3 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_8_3  (
            .in0(N__5587),
            .in1(N__5127),
            .in2(N__5108),
            .in3(N__5015),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_8_4 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_8_4  (
            .in0(N__5106),
            .in1(N__7481),
            .in2(N__5081),
            .in3(N__5078),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8677),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_1_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_1_LC_9_8_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_1_LC_9_8_5  (
            .in0(N__5262),
            .in1(N__5344),
            .in2(N__5333),
            .in3(N__5283),
            .lcout(\U712_REG_SM.m17_i_0_o2_1 ),
            .ltout(\U712_REG_SM.m17_i_0_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_m2_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_m2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_m2_LC_9_8_6 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_m2_LC_9_8_6  (
            .in0(N__5284),
            .in1(N__7036),
            .in2(N__5309),
            .in3(N__5263),
            .lcout(\U712_REG_SM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_8_7  (
            .in0(N__5306),
            .in1(N__9320),
            .in2(_gnd_net_),
            .in3(N__9512),
            .lcout(\U712_CHIP_RAM.N_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_9_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__5260),
            .in2(_gnd_net_),
            .in3(N__5282),
            .lcout(\U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1 ),
            .ltout(\U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_1_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_1_LC_9_9_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_1_LC_9_9_1  (
            .in0(N__7043),
            .in1(N__6206),
            .in2(N__5288),
            .in3(N__7703),
            .lcout(\U712_REG_SM.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__7160),
            .in2(_gnd_net_),
            .in3(N__7041),
            .lcout(\U712_REG_SM.N_270_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_0_LC_9_9_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_0_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__6952),
            .in2(_gnd_net_),
            .in3(N__6978),
            .lcout(),
            .ltout(\U712_REG_SM.m15_i_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_LC_9_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_LC_9_9_4  (
            .in0(N__5285),
            .in1(N__5261),
            .in2(N__5240),
            .in3(N__7042),
            .lcout(\U712_REG_SM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_9_5 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_9_9_5  (
            .in0(N__7044),
            .in1(N__6934),
            .in2(N__7166),
            .in3(N__6998),
            .lcout(\U712_REG_SM.REG_TACK_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_LC_9_9_6 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_LC_9_9_6  (
            .in0(N__6979),
            .in1(N__7164),
            .in2(N__6956),
            .in3(N__5627),
            .lcout(),
            .ltout(\U712_REG_SM.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_9_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_9_7  (
            .in0(N__7477),
            .in1(N__5611),
            .in2(N__5621),
            .in3(N__5618),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_9_10_0 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_9_10_0  (
            .in0(N__5612),
            .in1(N__5600),
            .in2(N__5588),
            .in3(N__5594),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8687),
            .ce(),
            .sr(N__10940));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_10_5  (
            .in0(N__5564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8687),
            .ce(),
            .sr(N__10940));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_11_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__10826),
            .in2(_gnd_net_),
            .in3(N__6201),
            .lcout(),
            .ltout(\U712_REG_SM.N_340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_11_1 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_11_1  (
            .in0(N__7382),
            .in1(N__5402),
            .in2(N__5525),
            .in3(N__5522),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8690),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_0_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_0_LC_9_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5497),
            .in2(_gnd_net_),
            .in3(N__5456),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__5401),
            .in2(_gnd_net_),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_9_13_3 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_9_13_3  (
            .in0(N__9441),
            .in1(N__10540),
            .in2(_gnd_net_),
            .in3(N__10460),
            .lcout(\U712_BYTE_ENABLE.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_9_13_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_9_13_5  (
            .in0(N__10632),
            .in1(N__10459),
            .in2(N__10170),
            .in3(N__9440),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_374_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_51_i_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_51_i_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_51_i_LC_9_13_6 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_51_i_LC_9_13_6  (
            .in0(N__8341),
            .in1(N__7957),
            .in2(N__5753),
            .in3(N__10714),
            .lcout(N_51_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_1_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_1_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_1_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_3_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_3_4  (
            .in0(N__5702),
            .in1(N__5687),
            .in2(_gnd_net_),
            .in3(N__9069),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_4_2 .LUT_INIT=16'b1111111011011010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_4_2  (
            .in0(N__5841),
            .in1(N__6776),
            .in2(N__6628),
            .in3(N__5959),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_4_3 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(N__6465),
            .in2(N__5669),
            .in3(N__7518),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8660),
            .ce(N__5654),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_4_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_4_5  (
            .in0(N__6349),
            .in1(N__6621),
            .in2(_gnd_net_),
            .in3(N__5842),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6  (
            .in0(N__7519),
            .in1(N__6466),
            .in2(N__5666),
            .in3(N__5663),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8660),
            .ce(N__5654),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_5_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_5_0  (
            .in0(N__8260),
            .in1(N__9008),
            .in2(_gnd_net_),
            .in3(N__8200),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_5_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_5_2  (
            .in0(N__6156),
            .in1(N__6133),
            .in2(_gnd_net_),
            .in3(N__6094),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_10_5_3 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_10_5_3  (
            .in0(N__6774),
            .in1(N__6618),
            .in2(_gnd_net_),
            .in3(N__5957),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_5_4 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__7517),
            .in2(N__6041),
            .in3(N__6348),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_5_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_5_5  (
            .in0(N__6038),
            .in1(N__5839),
            .in2(N__6032),
            .in3(N__6442),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_6  (
            .in0(N__6029),
            .in1(N__6023),
            .in2(N__6017),
            .in3(N__6014),
            .lcout(\U712_CHIP_RAM.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_5_7  (
            .in0(N__9009),
            .in1(N__5996),
            .in2(_gnd_net_),
            .in3(N__5975),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__6883),
            .in2(_gnd_net_),
            .in3(N__6604),
            .lcout(\U712_CHIP_RAM.CLK_EN_5_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_10_6_4 .LUT_INIT=16'b1001100111111111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_10_6_4  (
            .in0(N__6766),
            .in1(N__6603),
            .in2(_gnd_net_),
            .in3(N__5956),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_6_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_6_5  (
            .in0(N__6326),
            .in1(N__5840),
            .in2(N__5756),
            .in3(N__6464),
            .lcout(\U712_CHIP_RAM.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_7_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_7_1  (
            .in0(N__6775),
            .in1(N__6641),
            .in2(N__6629),
            .in3(N__6453),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_2  (
            .in0(N__7495),
            .in1(_gnd_net_),
            .in2(N__6371),
            .in3(N__6327),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8671),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_7_3  (
            .in0(N__6242),
            .in1(N__6224),
            .in2(_gnd_net_),
            .in3(N__9053),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIC74N_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIC74N_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIC74N_LC_10_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIC74N_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__6205),
            .in2(_gnd_net_),
            .in3(N__7702),
            .lcout(),
            .ltout(\U712_REG_SM.N_360_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI8VBS1_0_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI8VBS1_0_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI8VBS1_0_LC_10_9_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI8VBS1_0_LC_10_9_1  (
            .in0(N__6178),
            .in1(N__7159),
            .in2(N__6182),
            .in3(N__7037),
            .lcout(\U712_REG_SM.ASn_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_9_2 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_10_9_2  (
            .in0(N__7040),
            .in1(N__7446),
            .in2(N__7130),
            .in3(N__6999),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_LC_10_9_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_LC_10_9_3  (
            .in0(N__6950),
            .in1(N__7155),
            .in2(N__6179),
            .in3(N__6977),
            .lcout(\U712_REG_SM.m17_i_0_o2 ),
            .ltout(\U712_REG_SM.m17_i_0_o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_9_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_9_4  (
            .in0(N__7039),
            .in1(_gnd_net_),
            .in2(N__6167),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_9_5 .LUT_INIT=16'b1110111011000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_10_9_5  (
            .in0(N__7445),
            .in1(N__10816),
            .in2(N__6164),
            .in3(N__7118),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_a2_0_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_a2_0_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_a2_0_LC_10_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_a2_0_LC_10_9_6  (
            .in0(N__6976),
            .in1(N__6951),
            .in2(N__7165),
            .in3(N__7136),
            .lcout(\U712_REG_SM.N_435 ),
            .ltout(\U712_REG_SM.N_435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_9_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7121),
            .in3(N__7038),
            .lcout(\U712_REG_SM.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_10_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_10_10_0 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \U712_REG_SM.ASn_LC_10_10_0  (
            .in0(N__7074),
            .in1(N__7060),
            .in2(N__7051),
            .in3(N__7000),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8683),
            .ce(),
            .sr(N__10938));
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_10_10_4 .LUT_INIT=16'b1110111011001110;
    LogicCell40 \U712_REG_SM.DS_EN_LC_10_10_4  (
            .in0(N__10192),
            .in1(N__7061),
            .in2(N__7052),
            .in3(N__7001),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8683),
            .ce(),
            .sr(N__10938));
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6980),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8683),
            .ce(),
            .sr(N__10938));
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_10_19_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_LC_10_19_5 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_LC_10_19_5  (
            .in0(N__6930),
            .in1(N__10839),
            .in2(_gnd_net_),
            .in3(N__6893),
            .lcout(N_276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_3_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_3_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_3_1  (
            .in0(N__9454),
            .in1(N__6782),
            .in2(N__9114),
            .in3(N__8018),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_0  (
            .in0(N__8247),
            .in1(N__8204),
            .in2(N__8165),
            .in3(N__9073),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_5_6  (
            .in0(N__7292),
            .in1(N__7271),
            .in2(_gnd_net_),
            .in3(N__9060),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_7  (
            .in0(N__9061),
            .in1(N__9413),
            .in2(N__7250),
            .in3(N__10328),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_6_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_6_0 .LUT_INIT=16'b1111011100000111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_11_6_0  (
            .in0(N__7247),
            .in1(N__9456),
            .in2(N__7241),
            .in3(N__7213),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8666),
            .ce(),
            .sr(N__10951));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__7583),
            .in2(_gnd_net_),
            .in3(N__7202),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__7556),
            .in2(_gnd_net_),
            .in3(N__7199),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__7595),
            .in2(_gnd_net_),
            .in3(N__7196),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__7189),
            .in2(_gnd_net_),
            .in3(N__7175),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__7570),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__7616),
            .in2(_gnd_net_),
            .in3(N__7169),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__7628),
            .in2(_gnd_net_),
            .in3(N__7709),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__7640),
            .in2(_gnd_net_),
            .in3(N__7706),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7694),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_0  (
            .in0(N__7639),
            .in1(N__7627),
            .in2(_gnd_net_),
            .in3(N__7615),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_3 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_3  (
            .in0(N__7594),
            .in1(N__7582),
            .in2(N__7571),
            .in3(N__7555),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_11_11_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_11_11_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_11_11_6 (
            .in0(N__7381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3  (
            .in0(N__7298),
            .in1(N__7862),
            .in2(_gnd_net_),
            .in3(N__7313),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8655),
            .ce(N__8546),
            .sr(N__10962));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_4_2 .LUT_INIT=16'b0011111100101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_4_2  (
            .in0(N__8033),
            .in1(N__8825),
            .in2(N__9102),
            .in3(N__9443),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_4_3 .LUT_INIT=16'b0001000101000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_4_3  (
            .in0(N__8166),
            .in1(N__8262),
            .in2(N__8224),
            .in3(N__9074),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_4_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(N__8261),
            .in2(_gnd_net_),
            .in3(N__8219),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_7 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_7  (
            .in0(N__9442),
            .in1(N__8032),
            .in2(N__7865),
            .in3(N__9078),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_3  (
            .in0(N__9059),
            .in1(N__8826),
            .in2(_gnd_net_),
            .in3(N__7856),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_4  (
            .in0(N__7844),
            .in1(N__7832),
            .in2(_gnd_net_),
            .in3(N__9058),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_5 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_5  (
            .in0(N__8762),
            .in1(N__7810),
            .in2(N__8501),
            .in3(N__9452),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6 .LUT_INIT=16'b1010110011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6  (
            .in0(N__7811),
            .in1(N__8497),
            .in2(N__9470),
            .in3(N__8763),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_12_6_7  (
            .in0(N__7787),
            .in1(N__7781),
            .in2(_gnd_net_),
            .in3(N__7775),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8659),
            .ce(N__8576),
            .sr(N__10943));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_4  (
            .in0(N__7748),
            .in1(N__7733),
            .in2(_gnd_net_),
            .in3(N__9103),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5  (
            .in0(N__9104),
            .in1(N__9455),
            .in2(N__7712),
            .in3(N__8006),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_8_4  (
            .in0(N__9958),
            .in1(N__8414),
            .in2(_gnd_net_),
            .in3(N__8482),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9675),
            .sr(N__10937));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_5  (
            .in0(N__8483),
            .in1(N__9959),
            .in2(_gnd_net_),
            .in3(N__9584),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9675),
            .sr(N__10937));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_9_4  (
            .in0(N__8480),
            .in1(N__9957),
            .in2(_gnd_net_),
            .in3(N__8413),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9711),
            .ce(N__9673),
            .sr(N__10935));
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_10_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_12_10_5  (
            .in0(N__8000),
            .in1(N__9947),
            .in2(N__9783),
            .in3(N__7975),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10934));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_12_13_4 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_12_13_4  (
            .in0(N__10619),
            .in1(N__10161),
            .in2(N__9476),
            .in3(N__10468),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_55_i_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_55_i_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_55_i_LC_12_13_5 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_55_i_LC_12_13_5  (
            .in0(N__9496),
            .in1(N__7961),
            .in2(N__7946),
            .in3(N__10700),
            .lcout(N_55_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_13_1_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_13_1_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_13_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_13_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8223),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8654),
            .ce(),
            .sr(N__10977));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8174),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8656),
            .ce(),
            .sr(N__10974));
    defparam \U712_CHIP_RAM.RASn_LC_13_2_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8270),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8656),
            .ce(),
            .sr(N__10974));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_13_4_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_13_4_6  (
            .in0(N__8269),
            .in1(N__9111),
            .in2(N__8225),
            .in3(N__8173),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8658),
            .ce(N__8547),
            .sr(N__10964));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__10995),
            .in2(_gnd_net_),
            .in3(N__8120),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_5_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_5_2  (
            .in0(N__9448),
            .in1(N__8114),
            .in2(N__9095),
            .in3(N__8435),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__9447),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_13_6_6  (
            .in0(N__8895),
            .in1(N__8108),
            .in2(N__8867),
            .in3(N__8099),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8667),
            .ce(N__8563),
            .sr(N__10952));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_6_7  (
            .in0(N__8856),
            .in1(N__8896),
            .in2(N__8447),
            .in3(N__8039),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8667),
            .ce(N__8563),
            .sr(N__10952));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_4  (
            .in0(N__9460),
            .in1(N__8060),
            .in2(N__9115),
            .in3(N__8357),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_7_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_7_6  (
            .in0(N__9461),
            .in1(N__8051),
            .in2(N__9116),
            .in3(N__8423),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_1  (
            .in0(N__9950),
            .in1(N__8412),
            .in2(_gnd_net_),
            .in3(N__10304),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9712),
            .ce(N__9677),
            .sr(N__10941));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_5  (
            .in0(N__9620),
            .in1(_gnd_net_),
            .in2(N__9964),
            .in3(N__10064),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9712),
            .ce(N__9677),
            .sr(N__10941));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_7  (
            .in0(N__9583),
            .in1(_gnd_net_),
            .in2(N__9963),
            .in3(N__8481),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9712),
            .ce(N__9677),
            .sr(N__10941));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0  (
            .in0(N__9949),
            .in1(N__10057),
            .in2(_gnd_net_),
            .in3(N__9616),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9676),
            .sr(N__10939));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_9_5  (
            .in0(N__9615),
            .in1(N__9948),
            .in2(_gnd_net_),
            .in3(N__9581),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9676),
            .sr(N__10939));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_2  (
            .in0(N__8402),
            .in1(N__10300),
            .in2(_gnd_net_),
            .in3(N__9946),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9674),
            .sr(N__10936));
    defparam \U712_BYTE_ENABLE.N_53_i_LC_13_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_53_i_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_53_i_LC_13_12_2 .LUT_INIT=16'b0010101000111111;
    LogicCell40 \U712_BYTE_ENABLE.N_53_i_LC_13_12_2  (
            .in0(N__10780),
            .in1(N__8309),
            .in2(N__9475),
            .in3(N__8348),
            .lcout(N_53_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_0_o2_i_o2_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_0_o2_i_o2_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_0_o2_i_o2_LC_13_13_1 .LUT_INIT=16'b1111001000101111;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_0_o2_i_o2_LC_13_13_1  (
            .in0(N__10633),
            .in1(N__10178),
            .in2(N__10472),
            .in3(N__10544),
            .lcout(\U712_BYTE_ENABLE.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_0_o2_i_LC_13_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_o2_i_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_o2_i_LC_13_20_2 .LUT_INIT=16'b0000101110100000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_o2_i_LC_13_20_2  (
            .in0(N__10620),
            .in1(N__10179),
            .in2(N__10461),
            .in3(N__10524),
            .lcout(UMBE_0_o2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_13_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_13_20_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_LC_13_20_4  (
            .in0(N__10621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10180),
            .lcout(U712_BYTE_ENABLE_UUBE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_14_1_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_1_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9112),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8657),
            .ce(),
            .sr(N__10978));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_4_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_4_0  (
            .in0(N__8900),
            .in1(N__9521),
            .in2(N__8868),
            .in3(N__9188),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8661),
            .ce(N__8570),
            .sr(N__10968));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_4_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_4_7  (
            .in0(N__8770),
            .in1(N__9161),
            .in2(N__9469),
            .in3(N__10373),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8661),
            .ce(N__8570),
            .sr(N__10968));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_5_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_5_4  (
            .in0(N__9453),
            .in1(N__9125),
            .in2(N__9113),
            .in3(N__9638),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_5_5  (
            .in0(N__8863),
            .in1(N__8897),
            .in2(N__8942),
            .in3(N__9977),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8668),
            .ce(N__8572),
            .sr(N__10965));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_14_5_6  (
            .in0(N__8898),
            .in1(N__9629),
            .in2(N__8869),
            .in3(N__8924),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8668),
            .ce(N__8572),
            .sr(N__10965));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_6_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_6_0  (
            .in0(N__10223),
            .in1(N__8899),
            .in2(N__8870),
            .in3(N__8795),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8670),
            .ce(N__8571),
            .sr(N__10956));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1  (
            .in0(N__8771),
            .in1(N__8738),
            .in2(N__9474),
            .in3(N__9722),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8670),
            .ce(N__8571),
            .sr(N__10956));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_4  (
            .in0(N__9863),
            .in1(_gnd_net_),
            .in2(N__10019),
            .in3(N__10363),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__9681),
            .sr(N__10953));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1  (
            .in0(N__10362),
            .in1(N__10015),
            .in2(_gnd_net_),
            .in3(N__9907),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9710),
            .ce(N__9679),
            .sr(N__10944));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_7  (
            .in0(N__9614),
            .in1(N__9906),
            .in2(_gnd_net_),
            .in3(N__9582),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9710),
            .ce(N__9679),
            .sr(N__10944));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_9_4  (
            .in0(N__10014),
            .in1(N__9905),
            .in2(_gnd_net_),
            .in3(N__10056),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9678),
            .sr(N__10942));
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_12_5 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_57_i_LC_14_12_5  (
            .in0(N__10772),
            .in1(N__9497),
            .in2(N__9251),
            .in3(N__9468),
            .lcout(N_57_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_14_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_14_13_3 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_14_13_3  (
            .in0(N__10177),
            .in1(N__10634),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_BYTE_ENABLE.UUBE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_o2_i_LC_14_19_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_o2_i_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_o2_i_LC_14_19_0 .LUT_INIT=16'b0001000100101010;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_o2_i_LC_14_19_0  (
            .in0(N__10539),
            .in1(N__10583),
            .in2(N__10181),
            .in3(N__10453),
            .lcout(N_185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_3 .LUT_INIT=16'b0001111100001111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_3  (
            .in0(N__10452),
            .in1(N__10175),
            .in2(N__10210),
            .in3(N__10528),
            .lcout(N_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_303_i_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_303_i_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_303_i_LC_14_20_4 .LUT_INIT=16'b0000101110110000;
    LogicCell40 \U712_BYTE_ENABLE.N_303_i_LC_14_20_4  (
            .in0(N__10174),
            .in1(N__10628),
            .in2(N__10538),
            .in3(N__10451),
            .lcout(N_303_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_1  (
            .in0(N__9785),
            .in1(N__9944),
            .in2(_gnd_net_),
            .in3(N__10364),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9713),
            .ce(N__9685),
            .sr(N__10966));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_7_0  (
            .in0(N__9862),
            .in1(N__9784),
            .in2(_gnd_net_),
            .in3(N__10361),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__9683),
            .sr(N__10957));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_5  (
            .in0(N__10250),
            .in1(N__9904),
            .in2(_gnd_net_),
            .in3(N__10299),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__9682),
            .sr(N__10954));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_5  (
            .in0(N__9903),
            .in1(N__10281),
            .in2(_gnd_net_),
            .in3(N__10246),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9707),
            .ce(N__9680),
            .sr(N__10945));
    defparam \U712_BYTE_ENABLE.N_337_i_LC_15_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_337_i_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_337_i_LC_15_20_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_BYTE_ENABLE.N_337_i_LC_15_20_2  (
            .in0(N__10214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10176),
            .lcout(N_337_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_0  (
            .in0(N__10055),
            .in1(N__9911),
            .in2(_gnd_net_),
            .in3(N__10004),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9708),
            .ce(N__9684),
            .sr(N__10958));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_6_2  (
            .in0(N__9945),
            .in1(N__9800),
            .in2(_gnd_net_),
            .in3(N__9765),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9709),
            .ce(N__9686),
            .sr(N__10975));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_6  (
            .in0(N__10847),
            .in1(N__10768),
            .in2(_gnd_net_),
            .in3(N__10688),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

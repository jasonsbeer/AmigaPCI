-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Nov 28 2024 19:11:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    A : in std_logic_vector(31 downto 1);
    RnW : in std_logic;
    TT1 : in std_logic;
    TICK50 : out std_logic;
    nROMEN : out std_logic;
    nCIACS1 : out std_logic;
    TT0 : in std_logic;
    TICK60 : out std_logic;
    LBENn : in std_logic;
    CLKCIA : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    TSn : in std_logic;
    nBUFEN : out std_logic;
    nREGSPACE : out std_logic;
    nRAMSPACE : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    nCIACS0 : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2505\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_CIA.g0Z0Z_11_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.N_58\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\ : std_logic;
signal \U409_CIA.g0Z0Z_2_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_10\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\ : std_logic;
signal \nBUFEN_c\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nREGSPACE_i\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.N_23\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS1_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS0_i\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \ROMENm\ : std_logic;
signal \U409_TRANSFER_ACK.N_24_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_22\ : std_logic;
signal \bfn_10_5_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_22_0_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_24\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_49\ : std_logic;
signal \U409_TRANSFER_ACK.N_29_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_53\ : std_logic;
signal \U409_TRANSFER_ACK.N_52_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_29\ : std_logic;
signal \U409_TRANSFER_ACK.m9_i_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_54\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_60\ : std_logic;
signal \U409_TRANSFER_ACK.N_55\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_41\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_41_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_44_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_41_4\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_41_i\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5\ : std_logic;
signal \U409_TRANSFER_ACK.N_35\ : std_logic;
signal \U409_TRANSFER_ACK.N_44\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_391_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \nCIACS0_wire\ : std_logic;
signal \nCIACS1_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \nRAMSPACE_wire\ : std_logic;
signal \nROMEN_wire\ : std_logic;
signal \nBUFEN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \nREGSPACE_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    nCIACS0 <= \nCIACS0_wire\;
    nCIACS1 <= \nCIACS1_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    nRAMSPACE <= \nRAMSPACE_wire\;
    nROMEN <= \nROMEN_wire\;
    nBUFEN <= \nBUFEN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    nREGSPACE <= \nREGSPACE_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__5445\,
            RESETB => \N__5250\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6365\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6367\,
            DIN => \N__6366\,
            DOUT => \N__6365\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6367\,
            PADOUT => \N__6366\,
            PADIN => \N__6365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6355\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6357\,
            DIN => \N__6356\,
            DOUT => \N__6355\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6357\,
            PADOUT => \N__6356\,
            PADIN => \N__6355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6346\,
            DIN => \N__6345\,
            DOUT => \N__6344\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6346\,
            PADOUT => \N__6345\,
            PADIN => \N__6344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6337\,
            DIN => \N__6336\,
            DOUT => \N__6335\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6337\,
            PADOUT => \N__6336\,
            PADIN => \N__6335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6328\,
            DIN => \N__6327\,
            DOUT => \N__6326\,
            PACKAGEPIN => \nCIACS0_wire\
        );

    \nCIACS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6328\,
            PADOUT => \N__6327\,
            PADIN => \N__6326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3912\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6319\,
            DIN => \N__6318\,
            DOUT => \N__6317\,
            PACKAGEPIN => \nCIACS1_wire\
        );

    \nCIACS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6319\,
            PADOUT => \N__6318\,
            PADIN => \N__6317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6310\,
            DIN => \N__6309\,
            DOUT => \N__6308\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6310\,
            PADOUT => \N__6309\,
            PADIN => \N__6308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6301\,
            DIN => \N__6300\,
            DOUT => \N__6299\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6301\,
            PADOUT => \N__6300\,
            PADIN => \N__6299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6292\,
            DIN => \N__6291\,
            DOUT => \N__6290\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6292\,
            PADOUT => \N__6291\,
            PADIN => \N__6290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6283\,
            DIN => \N__6282\,
            DOUT => \N__6281\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6283\,
            PADOUT => \N__6282\,
            PADIN => \N__6281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5700\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__5301\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6274\,
            DIN => \N__6273\,
            DOUT => \N__6272\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6274\,
            PADOUT => \N__6273\,
            PADIN => \N__6272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6265\,
            DIN => \N__6264\,
            DOUT => \N__6263\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6265\,
            PADOUT => \N__6264\,
            PADIN => \N__6263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6256\,
            DIN => \N__6255\,
            DOUT => \N__6254\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6256\,
            PADOUT => \N__6255\,
            PADIN => \N__6254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2991\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nRAMSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6247\,
            DIN => \N__6246\,
            DOUT => \N__6245\,
            PACKAGEPIN => \nRAMSPACE_wire\
        );

    \nRAMSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6247\,
            PADOUT => \N__6246\,
            PADIN => \N__6245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3396\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nROMEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6238\,
            DIN => \N__6237\,
            DOUT => \N__6236\,
            PACKAGEPIN => \nROMEN_wire\
        );

    \nROMEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6238\,
            PADOUT => \N__6237\,
            PADIN => \N__6236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6229\,
            DIN => \N__6228\,
            DOUT => \N__6227\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6229\,
            PADOUT => \N__6228\,
            PADIN => \N__6227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6220\,
            DIN => \N__6219\,
            DOUT => \N__6218\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6220\,
            PADOUT => \N__6219\,
            PADIN => \N__6218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nBUFEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6211\,
            DIN => \N__6210\,
            DOUT => \N__6209\,
            PACKAGEPIN => \nBUFEN_wire\
        );

    \nBUFEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6211\,
            PADOUT => \N__6210\,
            PADIN => \N__6209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3294\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6202\,
            DIN => \N__6201\,
            DOUT => \N__6200\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6202\,
            PADOUT => \N__6201\,
            PADIN => \N__6200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6193\,
            DIN => \N__6192\,
            DOUT => \N__6191\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6193\,
            PADOUT => \N__6192\,
            PADIN => \N__6191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6184\,
            DIN => \N__6183\,
            DOUT => \N__6182\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6184\,
            PADOUT => \N__6183\,
            PADIN => \N__6182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6175\,
            DIN => \N__6174\,
            DOUT => \N__6173\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6175\,
            PADOUT => \N__6174\,
            PADIN => \N__6173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6166\,
            DIN => \N__6165\,
            DOUT => \N__6164\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6166\,
            PADOUT => \N__6165\,
            PADIN => \N__6164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6157\,
            DIN => \N__6156\,
            DOUT => \N__6155\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6157\,
            PADOUT => \N__6156\,
            PADIN => \N__6155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6148\,
            DIN => \N__6147\,
            DOUT => \N__6146\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6148\,
            PADOUT => \N__6147\,
            PADIN => \N__6146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nREGSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6139\,
            DIN => \N__6138\,
            DOUT => \N__6137\,
            PACKAGEPIN => \nREGSPACE_wire\
        );

    \nREGSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6139\,
            PADOUT => \N__6138\,
            PADIN => \N__6137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6130\,
            DIN => \N__6129\,
            DOUT => \N__6128\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6130\,
            PADOUT => \N__6129\,
            PADIN => \N__6128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4710\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6121\,
            DIN => \N__6120\,
            DOUT => \N__6119\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6121\,
            PADOUT => \N__6120\,
            PADIN => \N__6119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6112\,
            DIN => \N__6111\,
            DOUT => \N__6110\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6112\,
            PADOUT => \N__6111\,
            PADIN => \N__6110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6103\,
            DIN => \N__6102\,
            DOUT => \N__6101\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6103\,
            PADOUT => \N__6102\,
            PADIN => \N__6101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6094\,
            DIN => \N__6093\,
            DOUT => \N__6092\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6094\,
            PADOUT => \N__6093\,
            PADIN => \N__6092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6085\,
            DIN => \N__6084\,
            DOUT => \N__6083\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6085\,
            PADOUT => \N__6084\,
            PADIN => \N__6083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6076\,
            DIN => \N__6075\,
            DOUT => \N__6074\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6076\,
            PADOUT => \N__6075\,
            PADIN => \N__6074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6067\,
            DIN => \N__6066\,
            DOUT => \N__6065\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6067\,
            PADOUT => \N__6066\,
            PADIN => \N__6065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6058\,
            DIN => \N__6057\,
            DOUT => \N__6056\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6058\,
            PADOUT => \N__6057\,
            PADIN => \N__6056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__6039\,
            I => \N__6036\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6030\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6027\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6024\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6021\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6030\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6027\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6024\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6021\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6006\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__6003\,
            I => \N__5994\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5990\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5987\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5982\
        );

    \I__1381\ : InMux
    port map (
            O => \N__5999\,
            I => \N__5982\
        );

    \I__1380\ : InMux
    port map (
            O => \N__5998\,
            I => \N__5975\
        );

    \I__1379\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5975\
        );

    \I__1378\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5975\
        );

    \I__1377\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5972\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__5990\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__5987\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__5982\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__5975\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__5972\,
            I => \U409_TRANSFER_ACK.N_35\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__5961\,
            I => \N__5957\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__5960\,
            I => \N__5952\
        );

    \I__1369\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5945\
        );

    \I__1368\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5945\
        );

    \I__1367\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5938\
        );

    \I__1366\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5938\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5938\
        );

    \I__1364\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5935\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5945\,
            I => \U409_TRANSFER_ACK.N_44\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5938\,
            I => \U409_TRANSFER_ACK.N_44\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5935\,
            I => \U409_TRANSFER_ACK.N_44\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5928\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__5925\,
            I => \N__5920\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__5924\,
            I => \N__5917\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5914\
        );

    \I__1356\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5911\
        );

    \I__1355\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5908\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5905\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5900\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5900\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__5905\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__5900\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1349\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__1345\ : Span12Mux_h
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1344\ : Span12Mux_v
    port map (
            O => \N__5880\,
            I => \N__5877\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__5877\,
            I => \TACKn_in\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5870\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__5873\,
            I => \N__5867\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5870\,
            I => \N__5862\
        );

    \I__1339\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5859\
        );

    \I__1338\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5856\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__5865\,
            I => \N__5852\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__5862\,
            I => \N__5849\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__5859\,
            I => \N__5846\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5843\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5835\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5829\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__5849\,
            I => \N__5824\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__5846\,
            I => \N__5824\
        );

    \I__1329\ : Span4Mux_h
    port map (
            O => \N__5843\,
            I => \N__5821\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5818\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5809\
        );

    \I__1326\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5809\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5809\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5809\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5806\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5803\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5800\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5797\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5829\,
            I => \N__5792\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__5824\,
            I => \N__5792\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__5821\,
            I => \N__5785\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5818\,
            I => \N__5785\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__5809\,
            I => \N__5785\
        );

    \I__1314\ : Span4Mux_h
    port map (
            O => \N__5806\,
            I => \N__5778\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5778\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5800\,
            I => \N__5778\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5797\,
            I => \N__5775\
        );

    \I__1310\ : Span12Mux_h
    port map (
            O => \N__5792\,
            I => \N__5768\
        );

    \I__1309\ : Sp12to4
    port map (
            O => \N__5785\,
            I => \N__5768\
        );

    \I__1308\ : Sp12to4
    port map (
            O => \N__5778\,
            I => \N__5768\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__5775\,
            I => \N__5765\
        );

    \I__1306\ : Span12Mux_v
    port map (
            O => \N__5768\,
            I => \N__5762\
        );

    \I__1305\ : Span12Mux_v
    port map (
            O => \N__5765\,
            I => \N__5757\
        );

    \I__1304\ : Span12Mux_h
    port map (
            O => \N__5762\,
            I => \N__5757\
        );

    \I__1303\ : Odrv12
    port map (
            O => \N__5757\,
            I => \RESETn_c\
        );

    \I__1302\ : SRMux
    port map (
            O => \N__5754\,
            I => \N__5751\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5751\,
            I => \N__5746\
        );

    \I__1300\ : SRMux
    port map (
            O => \N__5750\,
            I => \N__5742\
        );

    \I__1299\ : SRMux
    port map (
            O => \N__5749\,
            I => \N__5739\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__5746\,
            I => \N__5736\
        );

    \I__1297\ : SRMux
    port map (
            O => \N__5745\,
            I => \N__5733\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5742\,
            I => \N__5730\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5727\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__5736\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__5733\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__5730\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__5727\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__1287\ : Span4Mux_h
    port map (
            O => \N__5709\,
            I => \N__5706\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__5706\,
            I => \N__5703\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__5703\,
            I => \TACK_EN_i\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__1282\ : Span4Mux_s3_v
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__1280\ : Sp12to4
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__5685\,
            I => \N_391_i\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5677\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5672\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5672\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5677\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5672\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__5667\,
            I => \N__5663\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5660\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5657\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5660\,
            I => \U409_TRANSFER_ACK.N_41_i\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5657\,
            I => \U409_TRANSFER_ACK.N_41_i\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5646\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5643\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5638\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5638\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5646\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5643\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5625\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5622\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__5619\,
            I => \N__5614\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5609\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5606\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5603\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5600\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5597\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5609\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5606\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5603\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5600\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5597\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5586\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5574\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5569\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5569\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5577\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5574\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5569\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5556\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5553\,
            I => \N__5547\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5544\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5541\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5538\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5547\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5544\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__5541\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5538\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5526\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5526\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5523\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5509\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5504\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5504\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5499\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5499\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5496\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5509\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5499\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5496\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5484\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5481\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__5472\,
            I => \N__5468\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5465\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__5468\,
            I => \N__5460\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5465\,
            I => \N__5460\
        );

    \I__1204\ : Span12Mux_h
    port map (
            O => \N__5460\,
            I => \N__5457\
        );

    \I__1203\ : Span12Mux_v
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__5454\,
            I => \TSn_c\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__5451\,
            I => \U409_TRANSFER_ACK.N_41_4_cascade_\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__5448\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_\
        );

    \I__1199\ : IoInMux
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5438\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5434\
        );

    \I__1196\ : IoSpan4Mux
    port map (
            O => \N__5438\,
            I => \N__5429\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5426\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5434\,
            I => \N__5423\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5420\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5417\
        );

    \I__1191\ : Span4Mux_s0_v
    port map (
            O => \N__5429\,
            I => \N__5414\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5426\,
            I => \N__5411\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__5423\,
            I => \N__5406\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5406\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5417\,
            I => \N__5403\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__5414\,
            I => \N__5400\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__5411\,
            I => \N__5397\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__5406\,
            I => \N__5392\
        );

    \I__1183\ : Span4Mux_h
    port map (
            O => \N__5403\,
            I => \N__5392\
        );

    \I__1182\ : Span12Mux_v
    port map (
            O => \N__5400\,
            I => \N__5389\
        );

    \I__1181\ : Sp12to4
    port map (
            O => \N__5397\,
            I => \N__5386\
        );

    \I__1180\ : Sp12to4
    port map (
            O => \N__5392\,
            I => \N__5383\
        );

    \I__1179\ : Span12Mux_v
    port map (
            O => \N__5389\,
            I => \N__5380\
        );

    \I__1178\ : Span12Mux_h
    port map (
            O => \N__5386\,
            I => \N__5377\
        );

    \I__1177\ : Span12Mux_v
    port map (
            O => \N__5383\,
            I => \N__5374\
        );

    \I__1176\ : Odrv12
    port map (
            O => \N__5380\,
            I => \CLK40_IN_c\
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__5377\,
            I => \CLK40_IN_c\
        );

    \I__1174\ : Odrv12
    port map (
            O => \N__5374\,
            I => \CLK40_IN_c\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__5367\,
            I => \U409_TRANSFER_ACK.N_44_cascade_\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__5364\,
            I => \N__5360\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5357\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5354\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5357\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5354\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__5349\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5342\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5339\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5342\,
            I => \U409_TRANSFER_ACK.N_41_4\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U409_TRANSFER_ACK.N_41_4\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5334\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5322\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5322\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5322\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5322\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5311\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5306\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5306\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5311\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5306\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1151\ : IoInMux
    port map (
            O => \N__5301\,
            I => \N__5298\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5298\,
            I => \N__5295\
        );

    \I__1149\ : IoSpan4Mux
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__1148\ : Span4Mux_s2_v
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__1147\ : Sp12to4
    port map (
            O => \N__5289\,
            I => \N__5286\
        );

    \I__1146\ : Span12Mux_v
    port map (
            O => \N__5286\,
            I => \N__5282\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__1144\ : Odrv12
    port map (
            O => \N__5282\,
            I => \TACK_OUTn\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5279\,
            I => \TACK_OUTn\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5270\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5267\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1138\ : CEMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__1136\ : Span4Mux_v
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__5253\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__1134\ : IoInMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__1132\ : Span4Mux_s3_v
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__1131\ : Span4Mux_h
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__5238\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5231\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5231\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5220\,
            I => \U409_TRANSFER_ACK.N_41\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5217\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5207\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5204\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5201\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5196\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5196\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5207\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5201\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__5187\,
            I => \N__5180\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5172\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5172\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5172\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5165\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5165\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5165\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5172\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5165\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5154\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__5159\,
            I => \N__5151\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__5158\,
            I => \N__5148\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__5157\,
            I => \N__5145\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5142\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5139\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5134\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5134\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__5142\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5139\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5134\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5124\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5124\,
            I => \U409_TRANSFER_ACK.N_53\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__5121\,
            I => \U409_TRANSFER_ACK.N_52_cascade_\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U409_TRANSFER_ACK.N_29\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__5112\,
            I => \U409_TRANSFER_ACK.m9_i_1_cascade_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5106\,
            I => \U409_TRANSFER_ACK.N_54\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5094\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5094\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5087\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5087\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5087\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5094\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5087\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5079\,
            I => \N__5074\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5071\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5068\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__5074\,
            I => \U409_TRANSFER_ACK.N_60\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U409_TRANSFER_ACK.N_60\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5068\,
            I => \U409_TRANSFER_ACK.N_60\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5058\,
            I => \U409_TRANSFER_ACK.N_55\
        );

    \I__1069\ : SRMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5052\,
            I => \N__5048\
        );

    \I__1067\ : SRMux
    port map (
            O => \N__5051\,
            I => \N__5045\
        );

    \I__1066\ : Span4Mux_v
    port map (
            O => \N__5048\,
            I => \N__5038\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__5038\
        );

    \I__1064\ : SRMux
    port map (
            O => \N__5044\,
            I => \N__5035\
        );

    \I__1063\ : SRMux
    port map (
            O => \N__5043\,
            I => \N__5032\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__5038\,
            I => \N__5027\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5035\,
            I => \N__5027\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__5024\
        );

    \I__1059\ : Span4Mux_v
    port map (
            O => \N__5027\,
            I => \N__5020\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__5024\,
            I => \N__5017\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5014\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__5020\,
            I => \RESETn_c_i\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__5017\,
            I => \RESETn_c_i\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5014\,
            I => \RESETn_c_i\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4997\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4994\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4997\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4994\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__4989\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4983\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4976\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4973\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4976\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4973\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4952\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4952\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4952\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4952\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4949\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4942\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4942\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4942\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4942\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4925\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4925\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__4933\,
            I => \N__4920\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__4932\,
            I => \N__4917\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4912\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4912\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4925\,
            I => \N__4909\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4900\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4900\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4900\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4900\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4912\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__4909\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4900\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__4893\,
            I => \N__4890\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__4884\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4863\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4863\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4863\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4863\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4863\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4856\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4856\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4856\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4856\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4847\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4844\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4844\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__997\ : ClkMux
    port map (
            O => \N__4839\,
            I => \N__4815\
        );

    \I__996\ : ClkMux
    port map (
            O => \N__4838\,
            I => \N__4815\
        );

    \I__995\ : ClkMux
    port map (
            O => \N__4837\,
            I => \N__4815\
        );

    \I__994\ : ClkMux
    port map (
            O => \N__4836\,
            I => \N__4815\
        );

    \I__993\ : ClkMux
    port map (
            O => \N__4835\,
            I => \N__4815\
        );

    \I__992\ : ClkMux
    port map (
            O => \N__4834\,
            I => \N__4815\
        );

    \I__991\ : ClkMux
    port map (
            O => \N__4833\,
            I => \N__4815\
        );

    \I__990\ : ClkMux
    port map (
            O => \N__4832\,
            I => \N__4815\
        );

    \I__989\ : GlobalMux
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__988\ : gio2CtrlBuf
    port map (
            O => \N__4812\,
            I => \CLK6_c_g\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__4809\,
            I => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\
        );

    \I__986\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4801\
        );

    \I__985\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4798\
        );

    \I__984\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4795\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4801\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4798\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4795\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__980\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4784\
        );

    \I__979\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4781\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4784\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4781\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__976\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U409_TRANSFER_ACK.N_49\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \U409_TRANSFER_ACK.N_29_cascade_\
        );

    \I__973\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4763\
        );

    \I__972\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4763\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__969\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4751\
        );

    \I__968\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4751\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4748\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__965\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4739\
        );

    \I__964\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4736\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4739\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__4731\,
            I => \N__4726\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__4730\,
            I => \N__4723\
        );

    \I__959\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4718\
        );

    \I__958\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4718\
        );

    \I__957\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4715\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__954\ : IoInMux
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4703\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__951\ : Span12Mux_s10_v
    port map (
            O => \N__4703\,
            I => \N__4697\
        );

    \I__950\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4694\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__4697\,
            I => \TICK50_c\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4694\,
            I => \TICK50_c\
        );

    \I__947\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4685\
        );

    \I__946\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4682\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__943\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4673\
        );

    \I__942\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4670\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4670\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__4665\,
            I => \N__4661\
        );

    \I__938\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4654\
        );

    \I__937\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4654\
        );

    \I__936\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4651\
        );

    \I__935\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4648\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4654\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4651\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4648\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__931\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U409_TICK.TICK503_11\
        );

    \I__929\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4631\
        );

    \I__928\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4628\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4631\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4628\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4616\
        );

    \I__923\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__920\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4605\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4602\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__916\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4592\
        );

    \I__915\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4592\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__912\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4581\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__909\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4571\
        );

    \I__908\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4568\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__904\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__4554\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__901\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4547\
        );

    \I__900\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4544\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__897\ : CEMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__4533\,
            I => \U409_TRANSFER_ACK.N_22_0_0\
        );

    \I__894\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4523\
        );

    \I__893\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4518\
        );

    \I__892\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4518\
        );

    \I__891\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4513\
        );

    \I__890\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4513\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4523\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4513\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__886\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4496\
        );

    \I__885\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4496\
        );

    \I__884\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4496\
        );

    \I__883\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4493\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4496\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4493\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__880\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4485\,
            I => \U409_TRANSFER_ACK.N_24\
        );

    \I__878\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4472\
        );

    \I__877\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4472\
        );

    \I__876\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4472\
        );

    \I__875\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4469\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4469\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__4464\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__871\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4458\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__869\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4451\
        );

    \I__868\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4448\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4448\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__865\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4439\
        );

    \I__864\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4436\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4439\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4436\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__861\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4427\
        );

    \I__860\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4427\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4424\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4419\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__856\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4413\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__854\ : InMux
    port map (
            O => \N__4410\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__853\ : InMux
    port map (
            O => \N__4407\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__852\ : InMux
    port map (
            O => \N__4404\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__851\ : InMux
    port map (
            O => \N__4401\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__850\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4395\,
            I => \N__4391\
        );

    \I__848\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4388\
        );

    \I__847\ : Span4Mux_h
    port map (
            O => \N__4391\,
            I => \N__4383\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4388\,
            I => \N__4383\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__4383\,
            I => \CIA_ENABLEm\
        );

    \I__844\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4377\,
            I => \N__4374\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__4374\,
            I => \N__4369\
        );

    \I__841\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4366\
        );

    \I__840\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4363\
        );

    \I__839\ : Sp12to4
    port map (
            O => \N__4369\,
            I => \N__4358\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4366\,
            I => \N__4358\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4363\,
            I => \N__4355\
        );

    \I__836\ : Span12Mux_h
    port map (
            O => \N__4358\,
            I => \N__4350\
        );

    \I__835\ : Span12Mux_v
    port map (
            O => \N__4355\,
            I => \N__4350\
        );

    \I__834\ : Odrv12
    port map (
            O => \N__4350\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__832\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4337\
        );

    \I__830\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4334\
        );

    \I__829\ : Span4Mux_h
    port map (
            O => \N__4337\,
            I => \N__4328\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4334\,
            I => \N__4328\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__4333\,
            I => \N__4325\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__4328\,
            I => \N__4322\
        );

    \I__825\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4319\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__4322\,
            I => \N__4316\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4319\,
            I => \N__4313\
        );

    \I__822\ : Span4Mux_h
    port map (
            O => \N__4316\,
            I => \N__4310\
        );

    \I__821\ : Span12Mux_v
    port map (
            O => \N__4313\,
            I => \N__4307\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__4310\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__819\ : Odrv12
    port map (
            O => \N__4307\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__817\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4295\
        );

    \I__816\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4292\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4295\,
            I => \N__4286\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4286\
        );

    \I__813\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4282\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__4286\,
            I => \N__4279\
        );

    \I__811\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4276\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4273\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__4279\,
            I => \U409_CIA.VMAZ0\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4276\,
            I => \U409_CIA.VMAZ0\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__4273\,
            I => \U409_CIA.VMAZ0\
        );

    \I__806\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4263\,
            I => \N__4259\
        );

    \I__804\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4256\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4259\,
            I => \N__4250\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__801\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4247\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__4250\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4247\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__796\ : Span4Mux_s1_v
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__4233\,
            I => \N__4229\
        );

    \I__794\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4226\
        );

    \I__793\ : Span12Mux_h
    port map (
            O => \N__4229\,
            I => \N__4223\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4226\,
            I => \N__4220\
        );

    \I__791\ : Span12Mux_v
    port map (
            O => \N__4223\,
            I => \N__4216\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__4220\,
            I => \N__4213\
        );

    \I__789\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4210\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4216\,
            I => \CLKCIA_c\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4213\,
            I => \CLKCIA_c\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4210\,
            I => \CLKCIA_c\
        );

    \I__785\ : InMux
    port map (
            O => \N__4203\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__784\ : InMux
    port map (
            O => \N__4200\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__783\ : InMux
    port map (
            O => \N__4197\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__782\ : InMux
    port map (
            O => \N__4194\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__781\ : InMux
    port map (
            O => \N__4191\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__780\ : InMux
    port map (
            O => \N__4188\,
            I => \bfn_10_6_0_\
        );

    \I__779\ : InMux
    port map (
            O => \N__4185\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__778\ : InMux
    port map (
            O => \N__4182\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__777\ : InMux
    port map (
            O => \N__4179\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__776\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4172\
        );

    \I__775\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4169\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4172\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4169\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__772\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4161\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__770\ : InMux
    port map (
            O => \N__4158\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__769\ : InMux
    port map (
            O => \N__4155\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__768\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4148\
        );

    \I__767\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4145\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4148\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4145\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__763\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__4131\,
            I => \ROMENm\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__4128\,
            I => \U409_TRANSFER_ACK.N_24_cascade_\
        );

    \I__759\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4122\,
            I => \U409_TRANSFER_ACK.N_22\
        );

    \I__757\ : InMux
    port map (
            O => \N__4119\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__756\ : InMux
    port map (
            O => \N__4116\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__755\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__754\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4109\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4106\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__751\ : InMux
    port map (
            O => \N__4101\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__750\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4094\
        );

    \I__749\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4091\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4094\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__746\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4083\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__744\ : InMux
    port map (
            O => \N__4080\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__743\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4073\
        );

    \I__742\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4070\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4073\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4070\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__739\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4062\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__737\ : InMux
    port map (
            O => \N__4059\,
            I => \bfn_9_8_0_\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__735\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4049\
        );

    \I__734\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4046\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4049\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4046\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__731\ : InMux
    port map (
            O => \N__4041\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__730\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4034\
        );

    \I__729\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4034\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__726\ : InMux
    port map (
            O => \N__4026\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__725\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4019\
        );

    \I__724\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4016\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4019\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4016\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__721\ : InMux
    port map (
            O => \N__4011\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__720\ : InMux
    port map (
            O => \N__4008\,
            I => \N__4004\
        );

    \I__719\ : InMux
    port map (
            O => \N__4007\,
            I => \N__4001\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4001\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__716\ : InMux
    port map (
            O => \N__3996\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__715\ : InMux
    port map (
            O => \N__3993\,
            I => \N__3989\
        );

    \I__714\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3986\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3989\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3986\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__711\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3978\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__709\ : InMux
    port map (
            O => \N__3975\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__708\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__3969\,
            I => \U409_TICK.TICK603_11\
        );

    \I__706\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__3960\,
            I => \N__3957\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__702\ : Span12Mux_h
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__701\ : Odrv12
    port map (
            O => \N__3951\,
            I => \A_c_13\
        );

    \I__700\ : IoInMux
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__698\ : IoSpan4Mux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__697\ : Sp12to4
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__696\ : Span12Mux_s7_h
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__695\ : Span12Mux_h
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__3930\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS1_i\
        );

    \I__693\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__689\ : Odrv12
    port map (
            O => \N__3915\,
            I => \A_c_12\
        );

    \I__688\ : IoInMux
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__686\ : Span4Mux_s0_h
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__685\ : Sp12to4
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__684\ : Span12Mux_s11_v
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__683\ : Span12Mux_h
    port map (
            O => \N__3897\,
            I => \N__3894\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__3894\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS0_i\
        );

    \I__681\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3886\
        );

    \I__680\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3883\
        );

    \I__679\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3880\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3886\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3883\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3880\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__3873\,
            I => \N__3867\
        );

    \I__674\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3862\
        );

    \I__673\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3862\
        );

    \I__672\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3859\
        );

    \I__671\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3856\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3862\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3859\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3856\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3849\,
            I => \N__3846\
        );

    \I__666\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3842\
        );

    \I__665\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3839\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3842\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3839\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__662\ : InMux
    port map (
            O => \N__3834\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__661\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3827\
        );

    \I__660\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3824\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3827\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3824\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__657\ : InMux
    port map (
            O => \N__3819\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__656\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3812\
        );

    \I__655\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3809\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3812\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3809\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__652\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3801\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__650\ : InMux
    port map (
            O => \N__3798\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__649\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3791\
        );

    \I__648\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3788\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3791\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3788\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__645\ : InMux
    port map (
            O => \N__3783\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__643\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3773\
        );

    \I__642\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3770\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3773\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3770\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__638\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3759\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__636\ : InMux
    port map (
            O => \N__3756\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__3753\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__3750\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3747\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3727\
        );

    \I__631\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3727\
        );

    \I__630\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3727\
        );

    \I__629\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3727\
        );

    \I__628\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3727\
        );

    \I__627\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3722\
        );

    \I__626\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3722\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3727\,
            I => \U409_TICK.TICK603_14\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3722\,
            I => \U409_TICK.TICK603_14\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__622\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3709\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3713\,
            I => \N__3706\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__3712\,
            I => \N__3700\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3696\
        );

    \I__618\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3691\
        );

    \I__617\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3691\
        );

    \I__616\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3688\
        );

    \I__615\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3681\
        );

    \I__614\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3681\
        );

    \I__613\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3681\
        );

    \I__612\ : Odrv4
    port map (
            O => \N__3696\,
            I => \U409_TICK.TICK603_9\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3691\,
            I => \U409_TICK.TICK603_9\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3688\,
            I => \U409_TICK.TICK603_9\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3681\,
            I => \U409_TICK.TICK603_9\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3672\,
            I => \N__3667\
        );

    \I__607\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3658\
        );

    \I__606\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3658\
        );

    \I__605\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3647\
        );

    \I__604\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3647\
        );

    \I__603\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3647\
        );

    \I__602\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3647\
        );

    \I__601\ : InMux
    port map (
            O => \N__3663\,
            I => \N__3647\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3658\,
            I => \U409_TICK.TICK603_10\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3647\,
            I => \U409_TICK.TICK603_10\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3642\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__3639\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__596\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3621\
        );

    \I__595\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3621\
        );

    \I__594\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3621\
        );

    \I__593\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3621\
        );

    \I__592\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3614\
        );

    \I__591\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3614\
        );

    \I__590\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3614\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3621\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3614\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3609\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__586\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3600\
        );

    \I__585\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3600\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3600\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__583\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3594\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__3591\,
            I => \N__3581\
        );

    \I__580\ : InMux
    port map (
            O => \N__3590\,
            I => \N__3578\
        );

    \I__579\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3569\
        );

    \I__578\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3569\
        );

    \I__577\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3569\
        );

    \I__576\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3569\
        );

    \I__575\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3562\
        );

    \I__574\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3562\
        );

    \I__573\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3562\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3578\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3569\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3562\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__3555\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__568\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3544\
        );

    \I__567\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3537\
        );

    \I__566\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3537\
        );

    \I__565\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3537\
        );

    \I__564\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3532\
        );

    \I__563\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3532\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3544\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3537\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3532\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__559\ : ClkMux
    port map (
            O => \N__3525\,
            I => \N__3513\
        );

    \I__558\ : ClkMux
    port map (
            O => \N__3524\,
            I => \N__3513\
        );

    \I__557\ : ClkMux
    port map (
            O => \N__3523\,
            I => \N__3513\
        );

    \I__556\ : ClkMux
    port map (
            O => \N__3522\,
            I => \N__3513\
        );

    \I__555\ : GlobalMux
    port map (
            O => \N__3513\,
            I => \N__3510\
        );

    \I__554\ : gio2CtrlBuf
    port map (
            O => \N__3510\,
            I => \CLK28_IN_c_g\
        );

    \I__553\ : IoInMux
    port map (
            O => \N__3507\,
            I => \N__3504\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3504\,
            I => \N__3501\
        );

    \I__551\ : Span4Mux_s1_v
    port map (
            O => \N__3501\,
            I => \N__3498\
        );

    \I__550\ : Sp12to4
    port map (
            O => \N__3498\,
            I => \N__3495\
        );

    \I__549\ : Span12Mux_h
    port map (
            O => \N__3495\,
            I => \N__3491\
        );

    \I__548\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3488\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__3491\,
            I => \TICK60_c\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3488\,
            I => \TICK60_c\
        );

    \I__545\ : InMux
    port map (
            O => \N__3483\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3480\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__543\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3474\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__540\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3462\
        );

    \I__539\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3462\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3462\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__537\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3453\
        );

    \I__536\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3448\
        );

    \I__535\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3448\
        );

    \I__534\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3445\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3453\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3448\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3445\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__530\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3430\
        );

    \I__529\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3430\
        );

    \I__528\ : InMux
    port map (
            O => \N__3436\,
            I => \N__3425\
        );

    \I__527\ : InMux
    port map (
            O => \N__3435\,
            I => \N__3425\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3430\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3425\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3420\,
            I => \N__3416\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3419\,
            I => \N__3412\
        );

    \I__522\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3406\
        );

    \I__521\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3406\
        );

    \I__520\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3401\
        );

    \I__519\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3401\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3406\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3401\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__516\ : IoInMux
    port map (
            O => \N__3396\,
            I => \N__3393\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__514\ : Span4Mux_s3_v
    port map (
            O => \N__3390\,
            I => \N__3387\
        );

    \I__513\ : Span4Mux_h
    port map (
            O => \N__3387\,
            I => \N__3384\
        );

    \I__512\ : Sp12to4
    port map (
            O => \N__3384\,
            I => \N__3381\
        );

    \I__511\ : Span12Mux_v
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__510\ : Odrv12
    port map (
            O => \N__3378\,
            I => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3375\,
            I => \N__3370\
        );

    \I__508\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3361\
        );

    \I__507\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3361\
        );

    \I__506\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3361\
        );

    \I__505\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3358\
        );

    \I__504\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3355\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3361\,
            I => \N__3352\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3358\,
            I => \N__3347\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3344\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__3352\,
            I => \N__3341\
        );

    \I__499\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3338\
        );

    \I__498\ : InMux
    port map (
            O => \N__3350\,
            I => \N__3335\
        );

    \I__497\ : Span12Mux_v
    port map (
            O => \N__3347\,
            I => \N__3330\
        );

    \I__496\ : Span12Mux_v
    port map (
            O => \N__3344\,
            I => \N__3330\
        );

    \I__495\ : Sp12to4
    port map (
            O => \N__3341\,
            I => \N__3323\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3323\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3335\,
            I => \N__3323\
        );

    \I__492\ : Odrv12
    port map (
            O => \N__3330\,
            I => \A_c_21\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__3323\,
            I => \A_c_21\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__489\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3312\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3312\,
            I => \N__3308\
        );

    \I__487\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3305\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__3308\,
            I => \U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3305\,
            I => \U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2\
        );

    \I__484\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3297\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3297\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__480\ : IoSpan4Mux
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__479\ : Span4Mux_s0_v
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__477\ : Span12Mux_s11_v
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__476\ : Span12Mux_h
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__3273\,
            I => \nBUFEN_c\
        );

    \I__474\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3264\
        );

    \I__473\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3258\
        );

    \I__472\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3255\
        );

    \I__471\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3252\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3264\,
            I => \N__3249\
        );

    \I__469\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3244\
        );

    \I__468\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3244\
        );

    \I__467\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3241\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3258\,
            I => \N__3238\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3255\,
            I => \N__3233\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3252\,
            I => \N__3233\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__3249\,
            I => \N__3228\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3244\,
            I => \N__3228\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3241\,
            I => \N__3225\
        );

    \I__460\ : Span4Mux_v
    port map (
            O => \N__3238\,
            I => \N__3219\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__3233\,
            I => \N__3219\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__3228\,
            I => \N__3214\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__3225\,
            I => \N__3214\
        );

    \I__456\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3211\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__3219\,
            I => \N__3204\
        );

    \I__454\ : Sp12to4
    port map (
            O => \N__3214\,
            I => \N__3204\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3211\,
            I => \N__3204\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__3204\,
            I => \A_c_23\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__450\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3195\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3195\,
            I => \N__3192\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__3192\,
            I => \N__3188\
        );

    \I__447\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3185\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__3188\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3185\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__444\ : IoInMux
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__442\ : Span4Mux_s3_v
    port map (
            O => \N__3174\,
            I => \N__3171\
        );

    \I__441\ : Span4Mux_h
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__440\ : Span4Mux_h
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__439\ : Sp12to4
    port map (
            O => \N__3165\,
            I => \N__3162\
        );

    \I__438\ : Span12Mux_s11_v
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__3159\,
            I => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\
        );

    \I__436\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3151\
        );

    \I__435\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3148\
        );

    \I__434\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3145\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3151\,
            I => \N__3141\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3148\,
            I => \N__3138\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3145\,
            I => \N__3135\
        );

    \I__430\ : InMux
    port map (
            O => \N__3144\,
            I => \N__3132\
        );

    \I__429\ : Span4Mux_h
    port map (
            O => \N__3141\,
            I => \N__3127\
        );

    \I__428\ : Span4Mux_h
    port map (
            O => \N__3138\,
            I => \N__3122\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__3135\,
            I => \N__3122\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3119\
        );

    \I__425\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3114\
        );

    \I__424\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3114\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__3127\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__422\ : Odrv4
    port map (
            O => \N__3122\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__421\ : Odrv12
    port map (
            O => \N__3119\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3114\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3102\,
            I => \N__3096\
        );

    \I__417\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3093\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3100\,
            I => \N__3090\
        );

    \I__415\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3086\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__3096\,
            I => \N__3081\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3093\,
            I => \N__3081\
        );

    \I__412\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3078\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3089\,
            I => \N__3075\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3086\,
            I => \N__3071\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__3081\,
            I => \N__3068\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3078\,
            I => \N__3065\
        );

    \I__407\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3060\
        );

    \I__406\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3060\
        );

    \I__405\ : Odrv12
    port map (
            O => \N__3071\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__3068\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__403\ : Odrv4
    port map (
            O => \N__3065\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3060\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__3051\,
            I => \N__3047\
        );

    \I__400\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3044\
        );

    \I__399\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3041\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3044\,
            I => \N__3036\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3041\,
            I => \N__3036\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__3033\,
            I => \U409_ADDRESS_DECODE.N_23\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__392\ : Span4Mux_s2_v
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__3021\,
            I => \N__3018\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__389\ : Sp12to4
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__3012\,
            I => \ROMENm_i\
        );

    \I__387\ : InMux
    port map (
            O => \N__3009\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__386\ : InMux
    port map (
            O => \N__3006\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__385\ : InMux
    port map (
            O => \N__3003\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__384\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2997\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2997\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2994\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2985\
        );

    \I__379\ : Span4Mux_s3_v
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__2976\,
            I => \PORTSIZE_0_i\
        );

    \I__375\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2963\
        );

    \I__374\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2963\
        );

    \I__373\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2963\
        );

    \I__372\ : InMux
    port map (
            O => \N__2970\,
            I => \N__2960\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N__2954\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2960\,
            I => \N__2954\
        );

    \I__369\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2951\
        );

    \I__368\ : Span4Mux_v
    port map (
            O => \N__2954\,
            I => \N__2945\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2951\,
            I => \N__2945\
        );

    \I__366\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2942\
        );

    \I__365\ : Span4Mux_h
    port map (
            O => \N__2945\,
            I => \N__2937\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2942\,
            I => \N__2937\
        );

    \I__363\ : Sp12to4
    port map (
            O => \N__2937\,
            I => \N__2934\
        );

    \I__362\ : Span12Mux_v
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__361\ : Odrv12
    port map (
            O => \N__2931\,
            I => \A_c_22\
        );

    \I__360\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2925\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__2922\,
            I => \U409_CIA.g0Z0Z_2_cascade_\
        );

    \I__357\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2916\,
            I => \U409_CIA.g0Z0Z_10\
        );

    \I__355\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2907\
        );

    \I__354\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2907\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2907\,
            I => \N__2904\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__2904\,
            I => \A_c_27\
        );

    \I__351\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2895\
        );

    \I__350\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2895\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2895\,
            I => \N__2892\
        );

    \I__348\ : Odrv12
    port map (
            O => \N__2892\,
            I => \A_c_25\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2889\,
            I => \N__2885\
        );

    \I__346\ : InMux
    port map (
            O => \N__2888\,
            I => \N__2880\
        );

    \I__345\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2880\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__343\ : Span4Mux_v
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__342\ : Span4Mux_v
    port map (
            O => \N__2874\,
            I => \N__2871\
        );

    \I__341\ : Span4Mux_h
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__2868\,
            I => \A_c_26\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__338\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2856\
        );

    \I__337\ : InMux
    port map (
            O => \N__2861\,
            I => \N__2856\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__335\ : Span4Mux_v
    port map (
            O => \N__2853\,
            I => \N__2850\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__333\ : Span4Mux_h
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__332\ : Odrv4
    port map (
            O => \N__2844\,
            I => \A_c_24\
        );

    \I__331\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2835\
        );

    \I__330\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2835\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2835\,
            I => \N__2832\
        );

    \I__328\ : Span4Mux_v
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__327\ : Sp12to4
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__326\ : Odrv12
    port map (
            O => \N__2826\,
            I => \A_c_31\
        );

    \I__325\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2817\
        );

    \I__324\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2817\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__322\ : Sp12to4
    port map (
            O => \N__2814\,
            I => \N__2811\
        );

    \I__321\ : Span12Mux_v
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__320\ : Odrv12
    port map (
            O => \N__2808\,
            I => \A_c_29\
        );

    \I__319\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2802\,
            I => \N__2798\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__2801\,
            I => \N__2795\
        );

    \I__316\ : Span4Mux_v
    port map (
            O => \N__2798\,
            I => \N__2792\
        );

    \I__315\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2789\
        );

    \I__314\ : Span4Mux_h
    port map (
            O => \N__2792\,
            I => \N__2784\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2789\,
            I => \N__2784\
        );

    \I__312\ : Span4Mux_v
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__311\ : Span4Mux_h
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__2778\,
            I => \A_c_30\
        );

    \I__309\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2771\
        );

    \I__308\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2768\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2771\,
            I => \N__2763\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2768\,
            I => \N__2763\
        );

    \I__305\ : Span4Mux_h
    port map (
            O => \N__2763\,
            I => \N__2760\
        );

    \I__304\ : Span4Mux_v
    port map (
            O => \N__2760\,
            I => \N__2757\
        );

    \I__303\ : Span4Mux_v
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__2754\,
            I => \A_c_28\
        );

    \I__301\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2745\
        );

    \I__300\ : InMux
    port map (
            O => \N__2750\,
            I => \N__2745\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__298\ : Span4Mux_v
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__297\ : Span4Mux_h
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__296\ : Span4Mux_v
    port map (
            O => \N__2736\,
            I => \N__2733\
        );

    \I__295\ : Span4Mux_v
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2730\,
            I => \A_c_18\
        );

    \I__293\ : CascadeMux
    port map (
            O => \N__2727\,
            I => \N__2723\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__2726\,
            I => \N__2720\
        );

    \I__291\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2717\
        );

    \I__290\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2714\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2717\,
            I => \N__2709\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2714\,
            I => \N__2709\
        );

    \I__287\ : Span4Mux_h
    port map (
            O => \N__2709\,
            I => \N__2706\
        );

    \I__286\ : Sp12to4
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__285\ : Span12Mux_v
    port map (
            O => \N__2703\,
            I => \N__2700\
        );

    \I__284\ : Odrv12
    port map (
            O => \N__2700\,
            I => \A_c_16\
        );

    \I__283\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2691\
        );

    \I__282\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2691\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2691\,
            I => \N__2688\
        );

    \I__280\ : Sp12to4
    port map (
            O => \N__2688\,
            I => \N__2685\
        );

    \I__279\ : Span12Mux_v
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__278\ : Odrv12
    port map (
            O => \N__2682\,
            I => \A_c_17\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__2679\,
            I => \U409_CIA.g0Z0Z_11_cascade_\
        );

    \I__276\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2673\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2673\,
            I => \N__2670\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2670\,
            I => \U409_CIA.g0Z0Z_8\
        );

    \I__273\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2664\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2664\,
            I => \N__2659\
        );

    \I__271\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2654\
        );

    \I__270\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2654\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2659\,
            I => \N__2651\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2654\,
            I => \N__2648\
        );

    \I__267\ : Sp12to4
    port map (
            O => \N__2651\,
            I => \N__2645\
        );

    \I__266\ : Span4Mux_h
    port map (
            O => \N__2648\,
            I => \N__2642\
        );

    \I__265\ : Span12Mux_s3_h
    port map (
            O => \N__2645\,
            I => \N__2637\
        );

    \I__264\ : Sp12to4
    port map (
            O => \N__2642\,
            I => \N__2637\
        );

    \I__263\ : Span12Mux_v
    port map (
            O => \N__2637\,
            I => \N__2634\
        );

    \I__262\ : Odrv12
    port map (
            O => \N__2634\,
            I => \A_c_19\
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__2631\,
            I => \U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_\
        );

    \I__260\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2625\,
            I => \U409_ADDRESS_DECODE.N_58\
        );

    \I__258\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2618\
        );

    \I__257\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2615\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2618\,
            I => \N__2610\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2615\,
            I => \N__2610\
        );

    \I__254\ : Span4Mux_v
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__253\ : Sp12to4
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__252\ : Span12Mux_h
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__251\ : Span12Mux_v
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__250\ : Span12Mux_h
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__249\ : Odrv12
    port map (
            O => \N__2595\,
            I => \OVL_c\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2592\,
            I => \N__2589\
        );

    \I__247\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2583\
        );

    \I__246\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2583\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2583\,
            I => \N__2580\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2580\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2577\,
            I => \N__2572\
        );

    \I__242\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2569\
        );

    \I__241\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2564\
        );

    \I__240\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2564\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2569\,
            I => \N__2561\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2564\,
            I => \N__2558\
        );

    \I__237\ : Span4Mux_v
    port map (
            O => \N__2561\,
            I => \N__2552\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__2558\,
            I => \N__2552\
        );

    \I__235\ : InMux
    port map (
            O => \N__2557\,
            I => \N__2549\
        );

    \I__234\ : Sp12to4
    port map (
            O => \N__2552\,
            I => \N__2544\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2549\,
            I => \N__2544\
        );

    \I__232\ : Odrv12
    port map (
            O => \N__2544\,
            I => \A_c_20\
        );

    \I__231\ : ClkMux
    port map (
            O => \N__2541\,
            I => \N__2505\
        );

    \I__230\ : ClkMux
    port map (
            O => \N__2540\,
            I => \N__2505\
        );

    \I__229\ : ClkMux
    port map (
            O => \N__2539\,
            I => \N__2505\
        );

    \I__228\ : ClkMux
    port map (
            O => \N__2538\,
            I => \N__2505\
        );

    \I__227\ : ClkMux
    port map (
            O => \N__2537\,
            I => \N__2505\
        );

    \I__226\ : ClkMux
    port map (
            O => \N__2536\,
            I => \N__2505\
        );

    \I__225\ : ClkMux
    port map (
            O => \N__2535\,
            I => \N__2505\
        );

    \I__224\ : ClkMux
    port map (
            O => \N__2534\,
            I => \N__2505\
        );

    \I__223\ : ClkMux
    port map (
            O => \N__2533\,
            I => \N__2505\
        );

    \I__222\ : ClkMux
    port map (
            O => \N__2532\,
            I => \N__2505\
        );

    \I__221\ : ClkMux
    port map (
            O => \N__2531\,
            I => \N__2505\
        );

    \I__220\ : ClkMux
    port map (
            O => \N__2530\,
            I => \N__2505\
        );

    \I__219\ : GlobalMux
    port map (
            O => \N__2505\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__2541\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2540\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2539\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__2534\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2537\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__2535\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2533\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2532\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2530\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            I => \N__2538\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net\,
            I => \N__2536\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2531\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_10_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_5_0_\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2662\,
            in1 => \N__2750\,
            in2 => \N__2726\,
            in3 => \N__2696\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2751\,
            in1 => \N__3270\,
            in2 => \N__2727\,
            in3 => \N__2663\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2576\,
            in1 => \N__2697\,
            in2 => \N__2679\,
            in3 => \N__2676\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__2973\,
            in1 => \N__3374\,
            in2 => \_gnd_net_\,
            in3 => \N__2805\,
            lcout => \U409_CIA.g0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a2_0_2_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2557\,
            in1 => \N__2971\,
            in2 => \_gnd_net_\,
            in3 => \N__3262\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_o2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__2667\,
            in1 => \N__3373\,
            in2 => \N__2631\,
            in3 => \N__2628\,
            lcout => \U409_ADDRESS_DECODE.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a2_1_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__2621\,
            in1 => \N__2972\,
            in2 => \N__3375\,
            in3 => \N__3263\,
            lcout => \U409_ADDRESS_DECODE.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_2_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2970\,
            in1 => \N__3144\,
            in2 => \N__3100\,
            in3 => \N__2622\,
            lcout => \U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3224\,
            in1 => \N__3350\,
            in2 => \N__2577\,
            in3 => \N__2588\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2959\,
            in1 => \N__3351\,
            in2 => \N__2592\,
            in3 => \N__2575\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3131\,
            in1 => \N__3261\,
            in2 => \N__3089\,
            in3 => \N__3191\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__3000\,
            in1 => \_gnd_net_\,
            in2 => \N__2994\,
            in3 => \N__2928\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2950\,
            in1 => \N__3130\,
            in2 => \N__5865\,
            in3 => \N__3074\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2823\,
            in2 => \_gnd_net_\,
            in3 => \N__5874\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2919\,
            in1 => \N__2841\,
            in2 => \N__2922\,
            in3 => \N__2775\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2901\,
            in1 => \N__2913\,
            in2 => \N__2865\,
            in3 => \N__2888\,
            lcout => \U409_CIA.g0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2912\,
            in1 => \N__2900\,
            in2 => \N__2889\,
            in3 => \N__2861\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2840\,
            in1 => \N__2822\,
            in2 => \N__2801\,
            in3 => \N__2774\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__3369\,
            in1 => \N__3269\,
            in2 => \_gnd_net_\,
            in3 => \N__3311\,
            lcout => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__3267\,
            in1 => \N__3368\,
            in2 => \N__3318\,
            in3 => \N__3300\,
            lcout => \nBUFEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3154\,
            in1 => \N__3268\,
            in2 => \N__3201\,
            in3 => \N__3101\,
            lcout => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3105\,
            in1 => \N__3156\,
            in2 => \N__3051\,
            in3 => \N__5866\,
            lcout => \ROMENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3155\,
            in1 => \N__3099\,
            in2 => \N__5873\,
            in3 => \N__3050\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3547\,
            in2 => \N__3591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3435\,
            in2 => \_gnd_net_\,
            in3 => \N__3009\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__3525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3630\,
            in2 => \_gnd_net_\,
            in3 => \N__3006\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3457\,
            in2 => \_gnd_net_\,
            in3 => \N__3003\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__3525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3415\,
            in2 => \_gnd_net_\,
            in3 => \N__3483\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__3632\,
            in1 => \N__3467\,
            in2 => \N__3480\,
            in3 => \N__3584\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101001100"
        )
    port map (
            in0 => \N__3585\,
            in1 => \N__3477\,
            in2 => \N__3471\,
            in3 => \N__3631\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3548\,
            in1 => \N__3458\,
            in2 => \N__3420\,
            in3 => \N__3436\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3590\,
            in2 => \_gnd_net_\,
            in3 => \N__3552\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3523\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4372\,
            in1 => \N__4291\,
            in2 => \N__4333\,
            in3 => \N__4255\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3411\,
            in1 => \N__3437\,
            in2 => \_gnd_net_\,
            in3 => \N__3456\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3588\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3459\,
            in1 => \N__3438\,
            in2 => \N__3419\,
            in3 => \N__3635\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__3634\,
            in1 => \N__3587\,
            in2 => \_gnd_net_\,
            in3 => \N__3550\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__4285\,
            in1 => \N__3636\,
            in2 => \N__3639\,
            in3 => \N__3606\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3633\,
            in1 => \N__3586\,
            in2 => \_gnd_net_\,
            in3 => \N__3549\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4219\,
            in2 => \N__3609\,
            in3 => \N__3605\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__3597\,
            in1 => \N__3589\,
            in2 => \N__3555\,
            in3 => \N__3551\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3871\,
            in2 => \_gnd_net_\,
            in3 => \N__3891\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__3741\,
            in1 => \N__3666\,
            in2 => \N__3717\,
            in3 => \N__3494\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3664\,
            in1 => \N__3744\,
            in2 => \N__3712\,
            in3 => \N__4086\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3740\,
            in1 => \N__3665\,
            in2 => \N__3765\,
            in3 => \N__3703\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__3699\,
            in1 => \N__3742\,
            in2 => \N__3672\,
            in3 => \N__3872\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4077\,
            in1 => \N__4098\,
            in2 => \N__3780\,
            in3 => \N__3993\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3663\,
            in1 => \N__3743\,
            in2 => \N__3753\,
            in3 => \N__3804\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3738\,
            in1 => \N__3671\,
            in2 => \N__3713\,
            in3 => \N__4065\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4113\,
            in1 => \N__4008\,
            in2 => \N__4056\,
            in3 => \N__4176\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3704\,
            in1 => \N__3739\,
            in2 => \N__3750\,
            in3 => \N__4164\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__3795\,
            in1 => \N__3816\,
            in2 => \_gnd_net_\,
            in3 => \N__3870\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3972\,
            in1 => \N__4038\,
            in2 => \N__3747\,
            in3 => \N__3831\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3705\,
            in1 => \N__3670\,
            in2 => \N__3642\,
            in3 => \N__3981\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__3890\,
            in2 => \N__3849\,
            in3 => \N__4151\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3966\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4394\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3889\,
            in2 => \N__3873\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3845\,
            in2 => \_gnd_net_\,
            in3 => \N__3834\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__4836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3830\,
            in2 => \_gnd_net_\,
            in3 => \N__3819\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__4836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3815\,
            in2 => \_gnd_net_\,
            in3 => \N__3798\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3794\,
            in2 => \_gnd_net_\,
            in3 => \N__3783\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__4836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3776\,
            in2 => \_gnd_net_\,
            in3 => \N__3756\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4112\,
            in2 => \_gnd_net_\,
            in3 => \N__4101\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__4836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4097\,
            in2 => \_gnd_net_\,
            in3 => \N__4080\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4076\,
            in2 => \_gnd_net_\,
            in3 => \N__4059\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4052\,
            in2 => \_gnd_net_\,
            in3 => \N__4041\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__4838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4037\,
            in2 => \_gnd_net_\,
            in3 => \N__4026\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__4838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4022\,
            in2 => \_gnd_net_\,
            in3 => \N__4011\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__4838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4007\,
            in2 => \_gnd_net_\,
            in3 => \N__3996\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__4838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3992\,
            in2 => \_gnd_net_\,
            in3 => \N__3975\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4175\,
            in2 => \_gnd_net_\,
            in3 => \N__4158\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4152\,
            in2 => \_gnd_net_\,
            in3 => \N__4155\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5855\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5023\,
            in2 => \_gnd_net_\,
            in3 => \N__4125\,
            lcout => \U409_TRANSFER_ACK.N_22_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI8GRM5_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__5471\,
            in1 => \N__5432\,
            in2 => \N__4140\,
            in3 => \N__4526\,
            lcout => \U409_TRANSFER_ACK.N_24\,
            ltout => \U409_TRANSFER_ACK.N_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111100"
        )
    port map (
            in0 => \N__4527\,
            in1 => \N__4503\,
            in2 => \N__4128\,
            in3 => \N__4479\,
            lcout => \U409_TRANSFER_ACK.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4659\,
            in2 => \N__4730\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4754\,
            in2 => \_gnd_net_\,
            in3 => \N__4119\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__4833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4676\,
            in2 => \_gnd_net_\,
            in3 => \N__4116\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__4833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4430\,
            in2 => \_gnd_net_\,
            in3 => \N__4203\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__4833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4688\,
            in2 => \_gnd_net_\,
            in3 => \N__4200\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4454\,
            in2 => \_gnd_net_\,
            in3 => \N__4197\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4442\,
            in2 => \_gnd_net_\,
            in3 => \N__4194\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__4833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4766\,
            in2 => \_gnd_net_\,
            in3 => \N__4191\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__4833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4850\,
            in2 => \_gnd_net_\,
            in3 => \N__4188\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4619\,
            in2 => \_gnd_net_\,
            in3 => \N__4185\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__4835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4595\,
            in2 => \_gnd_net_\,
            in3 => \N__4182\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4634\,
            in2 => \_gnd_net_\,
            in3 => \N__4179\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__4835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4550\,
            in2 => \_gnd_net_\,
            in3 => \N__4410\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4574\,
            in2 => \_gnd_net_\,
            in3 => \N__4407\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4979\,
            in2 => \_gnd_net_\,
            in3 => \N__4404\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4743\,
            in2 => \_gnd_net_\,
            in3 => \N__4401\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4298\,
            in1 => \N__4380\,
            in2 => \N__4347\,
            in3 => \N__4262\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__4373\,
            in1 => \N__4340\,
            in2 => \N__4302\,
            in3 => \N__4266\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5051\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5051\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4806\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5051\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5214\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5051\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4530\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net\,
            ce => \N__4539\,
            sr => \N__5044\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__4505\,
            in1 => \N__4481\,
            in2 => \_gnd_net_\,
            in3 => \N__4529\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5055\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__4504\,
            in1 => \N__4480\,
            in2 => \_gnd_net_\,
            in3 => \N__4528\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5055\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4506\,
            in1 => \N__4488\,
            in2 => \_gnd_net_\,
            in3 => \N__4482\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5055\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4551\,
            in1 => \N__4851\,
            in2 => \N__4599\,
            in3 => \N__4455\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4875\,
            in1 => \N__4934\,
            in2 => \N__4464\,
            in3 => \N__4461\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4961\,
            in1 => \N__4930\,
            in2 => \N__4665\,
            in3 => \N__4874\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__4443\,
            in2 => \N__4578\,
            in3 => \N__4431\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__4931\,
            in2 => \N__4419\,
            in3 => \N__4416\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4767\,
            in1 => \N__4755\,
            in2 => \N__4731\,
            in3 => \N__4742\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4664\,
            in1 => \N__4729\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4876\,
            in1 => \N__4963\,
            in2 => \N__4706\,
            in3 => \N__4935\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4689\,
            in1 => \N__4677\,
            in2 => \_gnd_net_\,
            in3 => \N__4660\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4641\,
            in1 => \N__4635\,
            in2 => \N__4623\,
            in3 => \N__4620\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__4608\,
            in1 => \N__4877\,
            in2 => \N__4602\,
            in3 => \N__4964\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4879\,
            in1 => \N__4966\,
            in2 => \N__4932\,
            in3 => \N__4584\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4965\,
            in1 => \N__4923\,
            in2 => \N__4563\,
            in3 => \N__4878\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4880\,
            in1 => \N__4967\,
            in2 => \N__4933\,
            in3 => \N__4986\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4968\,
            in1 => \N__4924\,
            in2 => \N__4893\,
            in3 => \N__4881\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5179\,
            in2 => \_gnd_net_\,
            in3 => \N__5099\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__5211\,
            in2 => \N__4809\,
            in3 => \N__5441\,
            lcout => \U409_TRANSFER_ACK.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__5210\,
            in1 => \N__5183\,
            in2 => \N__5159\,
            in3 => \N__5101\,
            lcout => \U409_TRANSFER_ACK.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5100\,
            in1 => \N__4788\,
            in2 => \N__5187\,
            in3 => \N__4805\,
            lcout => \U409_TRANSFER_ACK.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4804\,
            in2 => \_gnd_net_\,
            in3 => \N__4787\,
            lcout => \U409_TRANSFER_ACK.N_29\,
            ltout => \U409_TRANSFER_ACK.N_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__5833\,
            in1 => \N__4776\,
            in2 => \N__4770\,
            in3 => \N__5082\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5185\,
            in2 => \_gnd_net_\,
            in3 => \N__5102\,
            lcout => \U409_TRANSFER_ACK.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5433\,
            in1 => \N__5212\,
            in2 => \N__5157\,
            in3 => \N__5186\,
            lcout => \U409_TRANSFER_ACK.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__5213\,
            in1 => \N__5184\,
            in2 => \N__5158\,
            in3 => \N__5103\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__5077\,
            in1 => \N__5127\,
            in2 => \N__5121\,
            in3 => \N__5118\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__5834\,
            in1 => \_gnd_net_\,
            in2 => \N__5112\,
            in3 => \N__5109\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__5078\,
            in1 => \N__5061\,
            in2 => \_gnd_net_\,
            in3 => \N__5001\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5043\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__5330\,
            in1 => \N__5840\,
            in2 => \_gnd_net_\,
            in3 => \N__5314\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNIUBID_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5000\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNILJA71_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__5315\,
            in1 => \N__5329\,
            in2 => \N__4989\,
            in3 => \N__5234\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5334\,
            in3 => \N__5838\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5331\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101010"
        )
    port map (
            in0 => \N__5285\,
            in1 => \N__5841\,
            in2 => \N__5319\,
            in3 => \N__5274\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5273\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__5262\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__5235\,
            in1 => \N__5223\,
            in2 => \_gnd_net_\,
            in3 => \N__5993\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5754\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNO_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5514\,
            in1 => \N__5346\,
            in2 => \N__5364\,
            in3 => \N__5618\,
            lcout => \U409_TRANSFER_ACK.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIT7KM1_4_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__5513\,
            in1 => \N__6034\,
            in2 => \N__5619\,
            in3 => \N__5552\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CJV2_7_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__5923\,
            in1 => \N__5583\,
            in2 => \N__5217\,
            in3 => \N__5652\,
            lcout => \U409_TRANSFER_ACK.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011101100"
        )
    port map (
            in0 => \N__5681\,
            in1 => \N__5951\,
            in2 => \N__6003\,
            in3 => \N__5666\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5745\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_0_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5680\,
            in2 => \_gnd_net_\,
            in3 => \N__5580\,
            lcout => \U409_TRANSFER_ACK.N_41_4\,
            ltout => \U409_TRANSFER_ACK.N_41_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIGDB12_2_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5478\,
            in1 => \N__5617\,
            in2 => \N__5451\,
            in3 => \N__5515\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI772Q3_2_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5363\,
            in1 => \_gnd_net_\,
            in2 => \N__5448\,
            in3 => \N__5437\,
            lcout => \U409_TRANSFER_ACK.N_44\,
            ltout => \U409_TRANSFER_ACK.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__5581\,
            in1 => \N__6001\,
            in2 => \N__5367\,
            in3 => \N__5562\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5745\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__5516\,
            in1 => \N__5997\,
            in2 => \N__5960\,
            in3 => \N__5487\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5745\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__5998\,
            in1 => \N__5955\,
            in2 => \N__6039\,
            in3 => \N__6012\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5745\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIU8KM1_7_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5550\,
            in1 => \N__5649\,
            in2 => \N__5924\,
            in3 => \N__6033\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__5612\,
            in1 => \N__5512\,
            in2 => \N__5349\,
            in3 => \N__5345\,
            lcout => \U409_TRANSFER_ACK.N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__5999\,
            in1 => \N__5956\,
            in2 => \N__5631\,
            in3 => \N__5650\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__5553\,
            in1 => \N__6000\,
            in2 => \N__5961\,
            in3 => \N__5529\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5682\,
            in2 => \N__5667\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_LUT4_0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5651\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5613\,
            in2 => \_gnd_net_\,
            in3 => \N__5586\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2\,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_LUT4_0_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5582\,
            in2 => \_gnd_net_\,
            in3 => \N__5556\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_LUT4_0_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5551\,
            in2 => \_gnd_net_\,
            in3 => \N__5523\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_LUT4_0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5520\,
            in3 => \N__5481\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_LUT4_0_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6035\,
            in2 => \_gnd_net_\,
            in3 => \N__6006\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5\,
            carryout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__6002\,
            in1 => \N__5950\,
            in2 => \N__5925\,
            in3 => \N__5928\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5832\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5718\,
            lcout => \N_391_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

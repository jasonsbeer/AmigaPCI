// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 6 2025 20:26:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12772;
    wire N__12771;
    wire N__12770;
    wire N__12763;
    wire N__12762;
    wire N__12761;
    wire N__12754;
    wire N__12753;
    wire N__12752;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12736;
    wire N__12735;
    wire N__12734;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12718;
    wire N__12717;
    wire N__12716;
    wire N__12709;
    wire N__12708;
    wire N__12707;
    wire N__12700;
    wire N__12699;
    wire N__12698;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12682;
    wire N__12681;
    wire N__12680;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12664;
    wire N__12663;
    wire N__12662;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12646;
    wire N__12645;
    wire N__12644;
    wire N__12637;
    wire N__12636;
    wire N__12635;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12610;
    wire N__12609;
    wire N__12608;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12574;
    wire N__12573;
    wire N__12572;
    wire N__12565;
    wire N__12564;
    wire N__12563;
    wire N__12556;
    wire N__12555;
    wire N__12554;
    wire N__12547;
    wire N__12546;
    wire N__12545;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12529;
    wire N__12528;
    wire N__12527;
    wire N__12520;
    wire N__12519;
    wire N__12518;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12448;
    wire N__12447;
    wire N__12446;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12430;
    wire N__12429;
    wire N__12428;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12403;
    wire N__12402;
    wire N__12401;
    wire N__12394;
    wire N__12393;
    wire N__12392;
    wire N__12385;
    wire N__12384;
    wire N__12383;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12304;
    wire N__12303;
    wire N__12302;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12277;
    wire N__12276;
    wire N__12275;
    wire N__12268;
    wire N__12267;
    wire N__12266;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12232;
    wire N__12231;
    wire N__12230;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12214;
    wire N__12213;
    wire N__12212;
    wire N__12205;
    wire N__12204;
    wire N__12203;
    wire N__12196;
    wire N__12195;
    wire N__12194;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12142;
    wire N__12141;
    wire N__12140;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12088;
    wire N__12087;
    wire N__12086;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12070;
    wire N__12069;
    wire N__12068;
    wire N__12061;
    wire N__12060;
    wire N__12059;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12034;
    wire N__12033;
    wire N__12032;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12016;
    wire N__12015;
    wire N__12014;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11971;
    wire N__11970;
    wire N__11969;
    wire N__11962;
    wire N__11961;
    wire N__11960;
    wire N__11953;
    wire N__11952;
    wire N__11951;
    wire N__11944;
    wire N__11943;
    wire N__11942;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11917;
    wire N__11916;
    wire N__11915;
    wire N__11898;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11705;
    wire N__11702;
    wire N__11701;
    wire N__11698;
    wire N__11693;
    wire N__11692;
    wire N__11691;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11630;
    wire N__11627;
    wire N__11622;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11613;
    wire N__11612;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11567;
    wire N__11564;
    wire N__11557;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11538;
    wire N__11535;
    wire N__11528;
    wire N__11525;
    wire N__11520;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11468;
    wire N__11467;
    wire N__11466;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11374;
    wire N__11369;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11344;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11279;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11196;
    wire N__11191;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11175;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11155;
    wire N__11150;
    wire N__11147;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11110;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11055;
    wire N__11052;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11024;
    wire N__11021;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10977;
    wire N__10974;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10966;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10952;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10945;
    wire N__10944;
    wire N__10941;
    wire N__10936;
    wire N__10933;
    wire N__10932;
    wire N__10929;
    wire N__10922;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10896;
    wire N__10893;
    wire N__10892;
    wire N__10891;
    wire N__10890;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10883;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10844;
    wire N__10841;
    wire N__10832;
    wire N__10825;
    wire N__10818;
    wire N__10797;
    wire N__10796;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10785;
    wire N__10782;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10743;
    wire N__10742;
    wire N__10741;
    wire N__10738;
    wire N__10737;
    wire N__10736;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10730;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10722;
    wire N__10721;
    wire N__10720;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10714;
    wire N__10713;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10698;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10682;
    wire N__10679;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10643;
    wire N__10642;
    wire N__10631;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10565;
    wire N__10560;
    wire N__10559;
    wire N__10558;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10495;
    wire N__10494;
    wire N__10493;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10410;
    wire N__10409;
    wire N__10408;
    wire N__10407;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10401;
    wire N__10400;
    wire N__10397;
    wire N__10396;
    wire N__10395;
    wire N__10394;
    wire N__10393;
    wire N__10386;
    wire N__10385;
    wire N__10384;
    wire N__10383;
    wire N__10382;
    wire N__10381;
    wire N__10380;
    wire N__10375;
    wire N__10372;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10351;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10312;
    wire N__10309;
    wire N__10304;
    wire N__10301;
    wire N__10300;
    wire N__10297;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10257;
    wire N__10254;
    wire N__10253;
    wire N__10252;
    wire N__10247;
    wire N__10240;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10226;
    wire N__10221;
    wire N__10214;
    wire N__10209;
    wire N__10206;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10128;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10116;
    wire N__10115;
    wire N__10114;
    wire N__10113;
    wire N__10110;
    wire N__10105;
    wire N__10104;
    wire N__10103;
    wire N__10102;
    wire N__10101;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10093;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10071;
    wire N__10066;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10044;
    wire N__10041;
    wire N__10036;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9993;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9986;
    wire N__9985;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9977;
    wire N__9976;
    wire N__9975;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9941;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9831;
    wire N__9828;
    wire N__9827;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9799;
    wire N__9796;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9788;
    wire N__9787;
    wire N__9786;
    wire N__9785;
    wire N__9784;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9774;
    wire N__9773;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9756;
    wire N__9755;
    wire N__9754;
    wire N__9753;
    wire N__9752;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9746;
    wire N__9745;
    wire N__9744;
    wire N__9743;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9602;
    wire N__9601;
    wire N__9598;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9544;
    wire N__9543;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9483;
    wire N__9480;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9339;
    wire N__9336;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9287;
    wire N__9286;
    wire N__9283;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9251;
    wire N__9248;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9158;
    wire N__9155;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9049;
    wire N__9044;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8968;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8950;
    wire N__8949;
    wire N__8942;
    wire N__8939;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8914;
    wire N__8913;
    wire N__8912;
    wire N__8911;
    wire N__8906;
    wire N__8903;
    wire N__8898;
    wire N__8895;
    wire N__8886;
    wire N__8883;
    wire N__8882;
    wire N__8881;
    wire N__8878;
    wire N__8877;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8862;
    wire N__8853;
    wire N__8852;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8841;
    wire N__8838;
    wire N__8837;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8810;
    wire N__8805;
    wire N__8796;
    wire N__8787;
    wire N__8786;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8762;
    wire N__8759;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8688;
    wire N__8687;
    wire N__8686;
    wire N__8685;
    wire N__8682;
    wire N__8675;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8662;
    wire N__8657;
    wire N__8652;
    wire N__8649;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8641;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8598;
    wire N__8595;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8574;
    wire N__8573;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8502;
    wire N__8499;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8393;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8367;
    wire N__8366;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8358;
    wire N__8355;
    wire N__8354;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8342;
    wire N__8339;
    wire N__8338;
    wire N__8335;
    wire N__8334;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8330;
    wire N__8321;
    wire N__8316;
    wire N__8315;
    wire N__8314;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8306;
    wire N__8305;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8291;
    wire N__8290;
    wire N__8287;
    wire N__8286;
    wire N__8285;
    wire N__8284;
    wire N__8279;
    wire N__8272;
    wire N__8269;
    wire N__8260;
    wire N__8257;
    wire N__8252;
    wire N__8241;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8108;
    wire N__8107;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8095;
    wire N__8088;
    wire N__8087;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8067;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8049;
    wire N__8046;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8004;
    wire N__7997;
    wire N__7994;
    wire N__7989;
    wire N__7986;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7954;
    wire N__7951;
    wire N__7946;
    wire N__7941;
    wire N__7940;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7904;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7883;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7799;
    wire N__7798;
    wire N__7793;
    wire N__7790;
    wire N__7789;
    wire N__7788;
    wire N__7787;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7772;
    wire N__7769;
    wire N__7758;
    wire N__7757;
    wire N__7756;
    wire N__7755;
    wire N__7754;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7740;
    wire N__7737;
    wire N__7736;
    wire N__7733;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7721;
    wire N__7720;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7708;
    wire N__7705;
    wire N__7700;
    wire N__7695;
    wire N__7692;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7655;
    wire N__7654;
    wire N__7651;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7609;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7559;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7551;
    wire N__7548;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7524;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7494;
    wire N__7493;
    wire N__7492;
    wire N__7491;
    wire N__7490;
    wire N__7489;
    wire N__7488;
    wire N__7487;
    wire N__7486;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7440;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7404;
    wire N__7401;
    wire N__7396;
    wire N__7393;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7365;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7289;
    wire N__7286;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7238;
    wire N__7235;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7155;
    wire N__7152;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7140;
    wire N__7137;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7125;
    wire N__7122;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7107;
    wire N__7104;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7020;
    wire N__7019;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6988;
    wire N__6987;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6957;
    wire N__6954;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6885;
    wire N__6884;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6632;
    wire N__6631;
    wire N__6628;
    wire N__6627;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6609;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6589;
    wire N__6588;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6574;
    wire N__6567;
    wire N__6564;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6377;
    wire N__6376;
    wire N__6373;
    wire N__6368;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6338;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6311;
    wire N__6308;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6296;
    wire N__6291;
    wire N__6288;
    wire N__6287;
    wire N__6286;
    wire N__6283;
    wire N__6278;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6240;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6221;
    wire N__6220;
    wire N__6217;
    wire N__6216;
    wire N__6215;
    wire N__6214;
    wire N__6213;
    wire N__6212;
    wire N__6211;
    wire N__6210;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6199;
    wire N__6198;
    wire N__6197;
    wire N__6196;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6173;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6160;
    wire N__6155;
    wire N__6150;
    wire N__6139;
    wire N__6136;
    wire N__6125;
    wire N__6114;
    wire N__6099;
    wire N__6098;
    wire N__6097;
    wire N__6096;
    wire N__6095;
    wire N__6094;
    wire N__6093;
    wire N__6090;
    wire N__6089;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6070;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6062;
    wire N__6061;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6050;
    wire N__6049;
    wire N__6040;
    wire N__6031;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6022;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6008;
    wire N__6005;
    wire N__6000;
    wire N__5995;
    wire N__5990;
    wire N__5983;
    wire N__5976;
    wire N__5967;
    wire N__5946;
    wire N__5945;
    wire N__5942;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5877;
    wire N__5876;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5864;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5843;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5817;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5633;
    wire N__5630;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5576;
    wire N__5573;
    wire N__5572;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5550;
    wire N__5549;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5543;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5503;
    wire N__5502;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5484;
    wire N__5479;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5451;
    wire N__5450;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5441;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5433;
    wire N__5432;
    wire N__5429;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5419;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5387;
    wire N__5382;
    wire N__5379;
    wire N__5374;
    wire N__5355;
    wire N__5354;
    wire N__5353;
    wire N__5352;
    wire N__5349;
    wire N__5348;
    wire N__5343;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5328;
    wire N__5325;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5306;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5271;
    wire N__5270;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5250;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5242;
    wire N__5237;
    wire N__5236;
    wire N__5231;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5214;
    wire N__5213;
    wire N__5212;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5159;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5120;
    wire N__5117;
    wire N__5116;
    wire N__5115;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5111;
    wire N__5110;
    wire N__5105;
    wire N__5104;
    wire N__5099;
    wire N__5094;
    wire N__5091;
    wire N__5090;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5086;
    wire N__5085;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5066;
    wire N__5061;
    wire N__5054;
    wire N__5051;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4907;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4884;
    wire N__4881;
    wire N__4880;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4839;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4827;
    wire N__4824;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4812;
    wire N__4809;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4797;
    wire N__4794;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4761;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4691;
    wire N__4690;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4686;
    wire N__4679;
    wire N__4676;
    wire N__4669;
    wire N__4662;
    wire N__4659;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire REGSPACEn_c;
    wire \U712_CHIP_RAM.N_555_cascade_ ;
    wire \U712_CHIP_RAM.N_390_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_2 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ;
    wire bfn_7_7_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire A_c_8;
    wire A_c_2;
    wire A_c_3;
    wire A_c_4;
    wire A_c_7;
    wire A_c_5;
    wire A_c_18;
    wire \U712_CHIP_RAM.N_436_cascade_ ;
    wire \U712_CHIP_RAM.N_194_cascade_ ;
    wire \U712_CHIP_RAM.N_20_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.m101_i_1 ;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire \U712_CHIP_RAM.N_376 ;
    wire \U712_CHIP_RAM.m101_i_0_cascade_ ;
    wire \U712_CHIP_RAM.m101_i_2 ;
    wire \U712_CHIP_RAM.N_304_cascade_ ;
    wire \U712_CHIP_RAM.N_312_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.N_39 ;
    wire \U712_CHIP_RAM.N_326 ;
    wire \U712_CHIP_RAM.N_39_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_307_cascade_ ;
    wire \U712_CHIP_RAM.N_467_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_440 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_1 ;
    wire bfn_8_10_0_;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_3 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_4 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_5 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_7 ;
    wire DBRn_c;
    wire A_c_12;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_6 ;
    wire \U712_CHIP_RAM.N_194 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_378 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_CMDs_0_4 ;
    wire \U712_CHIP_RAM.N_396_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_0_2 ;
    wire \U712_CHIP_RAM.N_397 ;
    wire \U712_CHIP_RAM.N_555 ;
    wire \U712_CHIP_RAM.N_449 ;
    wire \U712_CHIP_RAM.SDRAM_CMDs_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_3 ;
    wire \U712_CHIP_RAM.N_194_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire CMA_c_6;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.m123_i_2 ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.N_190 ;
    wire \U712_CHIP_RAM.N_476 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_344 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.N_551_cascade_ ;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.N_435_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ;
    wire \U712_CHIP_RAM.N_325 ;
    wire \U712_CHIP_RAM.N_321 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_551 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ;
    wire \U712_CHIP_RAM.LATCH_CLK_6 ;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ;
    wire A_c_11;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.m93_i_a2_5 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_0 ;
    wire \U712_CHIP_RAM.m93_i_a2_4 ;
    wire \U712_CHIP_RAM.N_428_cascade_ ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.N_430 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CHIP_RAM.N_335_cascade_ ;
    wire N_202_i;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire N_165_i;
    wire WEn_c;
    wire RASn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire A_c_14;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ;
    wire A_c_9;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.N_361 ;
    wire CMA_c_5;
    wire A_c_10;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire A_c_13;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_435 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ;
    wire \U712_CHIP_RAM.N_467 ;
    wire \U712_CHIP_RAM.DBENn_7_0_0 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire DBDIR_c;
    wire TACK_OUTn;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.N_367 ;
    wire \U712_CHIP_RAM.N_419 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_10_10_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire DMA_CYCLEm;
    wire DBENn_c;
    wire \U712_REG_SM.N_402 ;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire CONSTANT_ONE_NET;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ;
    wire \U712_CHIP_RAM.N_314 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ;
    wire TACK_EN;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_REG_SM.N_373_cascade_ ;
    wire \U712_REG_SM.N_130 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_REG_SM.N_406 ;
    wire C3_c;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_328_cascade_ ;
    wire \U712_REG_SM.N_331_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_328 ;
    wire \U712_REG_SM.N_412 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.REGENn_e_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire REGENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.N_332 ;
    wire CPU_TACKm;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_455_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire \U712_REG_SM.N_373 ;
    wire \U712_REG_SM.N_330_cascade_ ;
    wire \U712_REG_SM.N_413 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_410 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.STATE_COUNTc_0_0 ;
    wire \U712_REG_SM.N_308 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_308_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire DRA_c_3;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire ASn_c;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ;
    wire N_336_i;
    wire DRA_c_0;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DRA_c_5;
    wire AGNUS_REV_c;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DBRn_c_i_0_g;
    wire RAS1n_c;
    wire RAS0n_c;
    wire RESETn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire LDSn_c;
    wire \U712_REG_SM.N_459 ;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire UDSn_c;
    wire CLK80_PLL;
    wire RESETn_c_i_g;
    wire \U712_REG_SM.N_404 ;
    wire N_335_i;
    wire N_337_i;
    wire N_177_i;
    wire N_334;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ;
    wire N_175_i;
    wire N_336;
    wire \U712_CHIP_RAM.m50_i_a2_0_0 ;
    wire \U712_CHIP_RAM.N_337_cascade_ ;
    wire N_200_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire N_334_i;
    wire RnW_c;
    wire DMA_WRITE_CYCLE;
    wire N_379;
    wire CASUn_c;
    wire CASLn_c;
    wire CPU_CYCLEm;
    wire REG_CYCLEm;
    wire N_167_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4344),
            .RESETB(N__7365),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12772),
            .DIN(N__12771),
            .DOUT(N__12770),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12772),
            .PADOUT(N__12771),
            .PADIN(N__12770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7422),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12763),
            .DIN(N__12762),
            .DOUT(N__12761),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12763),
            .PADOUT(N__12762),
            .PADIN(N__12761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12754),
            .DIN(N__12753),
            .DOUT(N__12752),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12754),
            .PADOUT(N__12753),
            .PADIN(N__12752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8226),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12745),
            .DIN(N__12744),
            .DOUT(N__12743),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12745),
            .PADOUT(N__12744),
            .PADIN(N__12743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11142),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12736),
            .DIN(N__12735),
            .DOUT(N__12734),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12736),
            .PADOUT(N__12735),
            .PADIN(N__12734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12727),
            .DIN(N__12726),
            .DOUT(N__12725),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12727),
            .PADOUT(N__12726),
            .PADIN(N__12725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12718),
            .DIN(N__12717),
            .DOUT(N__12716),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12718),
            .PADOUT(N__12717),
            .PADIN(N__12716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12709),
            .DIN(N__12708),
            .DOUT(N__12707),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12709),
            .PADOUT(N__12708),
            .PADIN(N__12707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12700),
            .DIN(N__12699),
            .DOUT(N__12698),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12700),
            .PADOUT(N__12699),
            .PADIN(N__12698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12691),
            .DIN(N__12690),
            .DOUT(N__12689),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12691),
            .PADOUT(N__12690),
            .PADIN(N__12689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12682),
            .DIN(N__12681),
            .DOUT(N__12680),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12682),
            .PADOUT(N__12681),
            .PADIN(N__12680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12673),
            .DIN(N__12672),
            .DOUT(N__12671),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12673),
            .PADOUT(N__12672),
            .PADIN(N__12671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7671),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12664),
            .DIN(N__12663),
            .DOUT(N__12662),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12664),
            .PADOUT(N__12663),
            .PADIN(N__12662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9408),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12655),
            .DIN(N__12654),
            .DOUT(N__12653),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12655),
            .PADOUT(N__12654),
            .PADIN(N__12653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12646),
            .DIN(N__12645),
            .DOUT(N__12644),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12646),
            .PADOUT(N__12645),
            .PADIN(N__12644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5910),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12637),
            .DIN(N__12636),
            .DOUT(N__12635),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12637),
            .PADOUT(N__12636),
            .PADIN(N__12635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12628),
            .DIN(N__12627),
            .DOUT(N__12626),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12628),
            .PADOUT(N__12627),
            .PADIN(N__12626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12619),
            .DIN(N__12618),
            .DOUT(N__12617),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12619),
            .PADOUT(N__12618),
            .PADIN(N__12617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4956),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12610),
            .DIN(N__12609),
            .DOUT(N__12608),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12610),
            .PADOUT(N__12609),
            .PADIN(N__12608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12601),
            .DIN(N__12600),
            .DOUT(N__12599),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12601),
            .PADOUT(N__12600),
            .PADIN(N__12599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12592),
            .DIN(N__12591),
            .DOUT(N__12590),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12592),
            .PADOUT(N__12591),
            .PADIN(N__12590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12583),
            .DIN(N__12582),
            .DOUT(N__12581),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12583),
            .PADOUT(N__12582),
            .PADIN(N__12581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12574),
            .DIN(N__12573),
            .DOUT(N__12572),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12574),
            .PADOUT(N__12573),
            .PADIN(N__12572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7335),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12565),
            .DIN(N__12564),
            .DOUT(N__12563),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12565),
            .PADOUT(N__12564),
            .PADIN(N__12563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12556),
            .DIN(N__12555),
            .DOUT(N__12554),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12556),
            .PADOUT(N__12555),
            .PADIN(N__12554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9630),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12547),
            .DIN(N__12546),
            .DOUT(N__12545),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12547),
            .PADOUT(N__12546),
            .PADIN(N__12545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8045),
            .DIN0(),
            .DOUT0(N__7289),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12538),
            .DIN(N__12537),
            .DOUT(N__12536),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12538),
            .PADOUT(N__12537),
            .PADIN(N__12536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12529),
            .DIN(N__12528),
            .DOUT(N__12527),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12529),
            .PADOUT(N__12528),
            .PADIN(N__12527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12520),
            .DIN(N__12519),
            .DOUT(N__12518),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12520),
            .PADOUT(N__12519),
            .PADIN(N__12518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12511),
            .DIN(N__12510),
            .DOUT(N__12509),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12511),
            .PADOUT(N__12510),
            .PADIN(N__12509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12502),
            .DIN(N__12501),
            .DOUT(N__12500),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12502),
            .PADOUT(N__12501),
            .PADIN(N__12500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12493),
            .DIN(N__12492),
            .DOUT(N__12491),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12493),
            .PADOUT(N__12492),
            .PADIN(N__12491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6441),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12484),
            .DIN(N__12483),
            .DOUT(N__12482),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12484),
            .PADOUT(N__12483),
            .PADIN(N__12482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12475),
            .DIN(N__12474),
            .DOUT(N__12473),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12475),
            .PADOUT(N__12474),
            .PADIN(N__12473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12466),
            .DIN(N__12465),
            .DOUT(N__12464),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12466),
            .PADOUT(N__12465),
            .PADIN(N__12464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12457),
            .DIN(N__12456),
            .DOUT(N__12455),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12457),
            .PADOUT(N__12456),
            .PADIN(N__12455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12448),
            .DIN(N__12447),
            .DOUT(N__12446),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12448),
            .PADOUT(N__12447),
            .PADIN(N__12446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12439),
            .DIN(N__12438),
            .DOUT(N__12437),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12439),
            .PADOUT(N__12438),
            .PADIN(N__12437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12430),
            .DIN(N__12429),
            .DOUT(N__12428),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12430),
            .PADOUT(N__12429),
            .PADIN(N__12428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12421),
            .DIN(N__12420),
            .DOUT(N__12419),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12421),
            .PADOUT(N__12420),
            .PADIN(N__12419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12412),
            .DIN(N__12411),
            .DOUT(N__12410),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12412),
            .PADOUT(N__12411),
            .PADIN(N__12410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9435),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12403),
            .DIN(N__12402),
            .DOUT(N__12401),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12403),
            .PADOUT(N__12402),
            .PADIN(N__12401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6563),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12394),
            .DIN(N__12393),
            .DOUT(N__12392),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12394),
            .PADOUT(N__12393),
            .PADIN(N__12392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12385),
            .DIN(N__12384),
            .DOUT(N__12383),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12385),
            .PADOUT(N__12384),
            .PADIN(N__12383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7878),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12376),
            .DIN(N__12375),
            .DOUT(N__12374),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12376),
            .PADOUT(N__12375),
            .PADIN(N__12374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12367),
            .DIN(N__12366),
            .DOUT(N__12365),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12367),
            .PADOUT(N__12366),
            .PADIN(N__12365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8403),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12358),
            .DIN(N__12357),
            .DOUT(N__12356),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12358),
            .PADOUT(N__12357),
            .PADIN(N__12356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12349),
            .DIN(N__12348),
            .DOUT(N__12347),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12349),
            .PADOUT(N__12348),
            .PADIN(N__12347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12340),
            .DIN(N__12339),
            .DOUT(N__12338),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12340),
            .PADOUT(N__12339),
            .PADIN(N__12338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12331),
            .DIN(N__12330),
            .DOUT(N__12329),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12331),
            .PADOUT(N__12330),
            .PADIN(N__12329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8049),
            .DIN0(),
            .DOUT0(N__7290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12322),
            .DIN(N__12321),
            .DOUT(N__12320),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12322),
            .PADOUT(N__12321),
            .PADIN(N__12320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6423),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12313),
            .DIN(N__12312),
            .DOUT(N__12311),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12313),
            .PADOUT(N__12312),
            .PADIN(N__12311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6867),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12304),
            .DIN(N__12303),
            .DOUT(N__12302),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12304),
            .PADOUT(N__12303),
            .PADIN(N__12302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11844),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12295),
            .DIN(N__12294),
            .DOUT(N__12293),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12295),
            .PADOUT(N__12294),
            .PADIN(N__12293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12286),
            .DIN(N__12285),
            .DOUT(N__12284),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12286),
            .PADOUT(N__12285),
            .PADIN(N__12284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12277),
            .DIN(N__12276),
            .DOUT(N__12275),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12277),
            .PADOUT(N__12276),
            .PADIN(N__12275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5805),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12268),
            .DIN(N__12267),
            .DOUT(N__12266),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12268),
            .PADOUT(N__12267),
            .PADIN(N__12266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12259),
            .DIN(N__12258),
            .DOUT(N__12257),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12259),
            .PADOUT(N__12258),
            .PADIN(N__12257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12250),
            .DIN(N__12249),
            .DOUT(N__12248),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12250),
            .PADOUT(N__12249),
            .PADIN(N__12248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6747),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12241),
            .DIN(N__12240),
            .DOUT(N__12239),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12241),
            .PADOUT(N__12240),
            .PADIN(N__12239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12232),
            .DIN(N__12231),
            .DOUT(N__12230),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12232),
            .PADOUT(N__12231),
            .PADIN(N__12230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12223),
            .DIN(N__12222),
            .DOUT(N__12221),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12223),
            .PADOUT(N__12222),
            .PADIN(N__12221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11787),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12214),
            .DIN(N__12213),
            .DOUT(N__12212),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12214),
            .PADOUT(N__12213),
            .PADIN(N__12212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8035),
            .DIN0(),
            .DOUT0(N__7285),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12205),
            .DIN(N__12204),
            .DOUT(N__12203),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12205),
            .PADOUT(N__12204),
            .PADIN(N__12203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7842),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12196),
            .DIN(N__12195),
            .DOUT(N__12194),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12196),
            .PADOUT(N__12195),
            .PADIN(N__12194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12187),
            .DIN(N__12186),
            .DOUT(N__12185),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12187),
            .PADOUT(N__12186),
            .PADIN(N__12185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12178),
            .DIN(N__12177),
            .DOUT(N__12176),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12178),
            .PADOUT(N__12177),
            .PADIN(N__12176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5700),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12169),
            .DIN(N__12168),
            .DOUT(N__12167),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12169),
            .PADOUT(N__12168),
            .PADIN(N__12167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12160),
            .DIN(N__12159),
            .DOUT(N__12158),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12160),
            .PADOUT(N__12159),
            .PADIN(N__12158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12151),
            .DIN(N__12150),
            .DOUT(N__12149),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12151),
            .PADOUT(N__12150),
            .PADIN(N__12149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6813),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12142),
            .DIN(N__12141),
            .DOUT(N__12140),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12142),
            .PADOUT(N__12141),
            .PADIN(N__12140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12133),
            .DIN(N__12132),
            .DOUT(N__12131),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12133),
            .PADOUT(N__12132),
            .PADIN(N__12131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12124),
            .DIN(N__12123),
            .DOUT(N__12122),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12124),
            .PADOUT(N__12123),
            .PADIN(N__12122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6837),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12115),
            .DIN(N__12114),
            .DOUT(N__12113),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12115),
            .PADOUT(N__12114),
            .PADIN(N__12113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10023),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12106),
            .DIN(N__12105),
            .DOUT(N__12104),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12106),
            .PADOUT(N__12105),
            .PADIN(N__12104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11274),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12097),
            .DIN(N__12096),
            .DOUT(N__12095),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12097),
            .PADOUT(N__12096),
            .PADIN(N__12095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4446),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12088),
            .DIN(N__12087),
            .DOUT(N__12086),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12088),
            .PADOUT(N__12087),
            .PADIN(N__12086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12079),
            .DIN(N__12078),
            .DOUT(N__12077),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12079),
            .PADOUT(N__12078),
            .PADIN(N__12077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12070),
            .DIN(N__12069),
            .DOUT(N__12068),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12070),
            .PADOUT(N__12069),
            .PADIN(N__12068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5028),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12061),
            .DIN(N__12060),
            .DOUT(N__12059),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12061),
            .PADOUT(N__12060),
            .PADIN(N__12059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12052),
            .DIN(N__12051),
            .DOUT(N__12050),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12052),
            .PADOUT(N__12051),
            .PADIN(N__12050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12043),
            .DIN(N__12042),
            .DOUT(N__12041),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12043),
            .PADOUT(N__12042),
            .PADIN(N__12041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12034),
            .DIN(N__12033),
            .DOUT(N__12032),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12034),
            .PADOUT(N__12033),
            .PADIN(N__12032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10170),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12025),
            .DIN(N__12024),
            .DOUT(N__12023),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12025),
            .PADOUT(N__12024),
            .PADIN(N__12023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12016),
            .DIN(N__12015),
            .DOUT(N__12014),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12016),
            .PADOUT(N__12015),
            .PADIN(N__12014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12007),
            .DIN(N__12006),
            .DOUT(N__12005),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12007),
            .PADOUT(N__12006),
            .PADIN(N__12005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8513),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11998),
            .DIN(N__11997),
            .DOUT(N__11996),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11998),
            .PADOUT(N__11997),
            .PADIN(N__11996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11989),
            .DIN(N__11988),
            .DOUT(N__11987),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11989),
            .PADOUT(N__11988),
            .PADIN(N__11987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6669),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11980),
            .DIN(N__11979),
            .DOUT(N__11978),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11980),
            .PADOUT(N__11979),
            .PADIN(N__11978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11971),
            .DIN(N__11970),
            .DOUT(N__11969),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11971),
            .PADOUT(N__11970),
            .PADIN(N__11969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11962),
            .DIN(N__11961),
            .DOUT(N__11960),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11962),
            .PADOUT(N__11961),
            .PADIN(N__11960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11953),
            .DIN(N__11952),
            .DOUT(N__11951),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11953),
            .PADOUT(N__11952),
            .PADIN(N__11951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11944),
            .DIN(N__11943),
            .DOUT(N__11942),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11944),
            .PADOUT(N__11943),
            .PADIN(N__11942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8498),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11935),
            .DIN(N__11934),
            .DOUT(N__11933),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11935),
            .PADOUT(N__11934),
            .PADIN(N__11933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11859),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11926),
            .DIN(N__11925),
            .DOUT(N__11924),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11926),
            .PADOUT(N__11925),
            .PADIN(N__11924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6501),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11917),
            .DIN(N__11916),
            .DOUT(N__11915),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11917),
            .PADOUT(N__11916),
            .PADIN(N__11915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5655),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2899 (
            .O(N__11898),
            .I(N__11894));
    InMux I__2898 (
            .O(N__11897),
            .I(N__11891));
    LocalMux I__2897 (
            .O(N__11894),
            .I(N__11888));
    LocalMux I__2896 (
            .O(N__11891),
            .I(N__11885));
    Span12Mux_v I__2895 (
            .O(N__11888),
            .I(N__11881));
    Span4Mux_v I__2894 (
            .O(N__11885),
            .I(N__11878));
    CascadeMux I__2893 (
            .O(N__11884),
            .I(N__11875));
    Span12Mux_h I__2892 (
            .O(N__11881),
            .I(N__11872));
    Span4Mux_v I__2891 (
            .O(N__11878),
            .I(N__11869));
    InMux I__2890 (
            .O(N__11875),
            .I(N__11866));
    Odrv12 I__2889 (
            .O(N__11872),
            .I(REG_CYCLEm));
    Odrv4 I__2888 (
            .O(N__11869),
            .I(REG_CYCLEm));
    LocalMux I__2887 (
            .O(N__11866),
            .I(REG_CYCLEm));
    IoInMux I__2886 (
            .O(N__11859),
            .I(N__11856));
    LocalMux I__2885 (
            .O(N__11856),
            .I(N__11853));
    Span4Mux_s3_v I__2884 (
            .O(N__11853),
            .I(N__11850));
    Span4Mux_v I__2883 (
            .O(N__11850),
            .I(N__11847));
    Odrv4 I__2882 (
            .O(N__11847),
            .I(N_167_i));
    IoInMux I__2881 (
            .O(N__11844),
            .I(N__11841));
    LocalMux I__2880 (
            .O(N__11841),
            .I(N__11838));
    Span4Mux_s3_h I__2879 (
            .O(N__11838),
            .I(N__11835));
    Span4Mux_h I__2878 (
            .O(N__11835),
            .I(N__11832));
    Span4Mux_h I__2877 (
            .O(N__11832),
            .I(N__11829));
    Sp12to4 I__2876 (
            .O(N__11829),
            .I(N__11826));
    Span12Mux_v I__2875 (
            .O(N__11826),
            .I(N__11823));
    Odrv12 I__2874 (
            .O(N__11823),
            .I(N_177_i));
    CascadeMux I__2873 (
            .O(N__11820),
            .I(N__11817));
    InMux I__2872 (
            .O(N__11817),
            .I(N__11814));
    LocalMux I__2871 (
            .O(N__11814),
            .I(N__11811));
    Odrv4 I__2870 (
            .O(N__11811),
            .I(N_334));
    InMux I__2869 (
            .O(N__11808),
            .I(N__11805));
    LocalMux I__2868 (
            .O(N__11805),
            .I(N__11801));
    InMux I__2867 (
            .O(N__11804),
            .I(N__11798));
    Span4Mux_h I__2866 (
            .O(N__11801),
            .I(N__11793));
    LocalMux I__2865 (
            .O(N__11798),
            .I(N__11793));
    Span4Mux_h I__2864 (
            .O(N__11793),
            .I(N__11790));
    Odrv4 I__2863 (
            .O(N__11790),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ));
    IoInMux I__2862 (
            .O(N__11787),
            .I(N__11784));
    LocalMux I__2861 (
            .O(N__11784),
            .I(N__11781));
    IoSpan4Mux I__2860 (
            .O(N__11781),
            .I(N__11778));
    Span4Mux_s3_h I__2859 (
            .O(N__11778),
            .I(N__11775));
    Span4Mux_v I__2858 (
            .O(N__11775),
            .I(N__11772));
    Span4Mux_h I__2857 (
            .O(N__11772),
            .I(N__11769));
    Odrv4 I__2856 (
            .O(N__11769),
            .I(N_175_i));
    CascadeMux I__2855 (
            .O(N__11766),
            .I(N__11763));
    InMux I__2854 (
            .O(N__11763),
            .I(N__11760));
    LocalMux I__2853 (
            .O(N__11760),
            .I(N__11757));
    Odrv4 I__2852 (
            .O(N__11757),
            .I(N_336));
    InMux I__2851 (
            .O(N__11754),
            .I(N__11751));
    LocalMux I__2850 (
            .O(N__11751),
            .I(N__11748));
    Span4Mux_v I__2849 (
            .O(N__11748),
            .I(N__11744));
    InMux I__2848 (
            .O(N__11747),
            .I(N__11741));
    Sp12to4 I__2847 (
            .O(N__11744),
            .I(N__11738));
    LocalMux I__2846 (
            .O(N__11741),
            .I(N__11735));
    Odrv12 I__2845 (
            .O(N__11738),
            .I(\U712_CHIP_RAM.m50_i_a2_0_0 ));
    Odrv4 I__2844 (
            .O(N__11735),
            .I(\U712_CHIP_RAM.m50_i_a2_0_0 ));
    CascadeMux I__2843 (
            .O(N__11730),
            .I(\U712_CHIP_RAM.N_337_cascade_ ));
    IoInMux I__2842 (
            .O(N__11727),
            .I(N__11724));
    LocalMux I__2841 (
            .O(N__11724),
            .I(N__11721));
    IoSpan4Mux I__2840 (
            .O(N__11721),
            .I(N__11718));
    Sp12to4 I__2839 (
            .O(N__11718),
            .I(N__11715));
    Span12Mux_s7_v I__2838 (
            .O(N__11715),
            .I(N__11712));
    Span12Mux_v I__2837 (
            .O(N__11712),
            .I(N__11709));
    Odrv12 I__2836 (
            .O(N__11709),
            .I(N_200_i));
    CascadeMux I__2835 (
            .O(N__11706),
            .I(N__11702));
    InMux I__2834 (
            .O(N__11705),
            .I(N__11698));
    InMux I__2833 (
            .O(N__11702),
            .I(N__11693));
    InMux I__2832 (
            .O(N__11701),
            .I(N__11693));
    LocalMux I__2831 (
            .O(N__11698),
            .I(N__11685));
    LocalMux I__2830 (
            .O(N__11693),
            .I(N__11682));
    InMux I__2829 (
            .O(N__11692),
            .I(N__11679));
    InMux I__2828 (
            .O(N__11691),
            .I(N__11674));
    InMux I__2827 (
            .O(N__11690),
            .I(N__11674));
    InMux I__2826 (
            .O(N__11689),
            .I(N__11671));
    InMux I__2825 (
            .O(N__11688),
            .I(N__11668));
    Span4Mux_v I__2824 (
            .O(N__11685),
            .I(N__11665));
    Span4Mux_v I__2823 (
            .O(N__11682),
            .I(N__11662));
    LocalMux I__2822 (
            .O(N__11679),
            .I(N__11659));
    LocalMux I__2821 (
            .O(N__11674),
            .I(N__11654));
    LocalMux I__2820 (
            .O(N__11671),
            .I(N__11654));
    LocalMux I__2819 (
            .O(N__11668),
            .I(N__11651));
    Span4Mux_v I__2818 (
            .O(N__11665),
            .I(N__11648));
    Span4Mux_v I__2817 (
            .O(N__11662),
            .I(N__11643));
    Span4Mux_v I__2816 (
            .O(N__11659),
            .I(N__11643));
    Span4Mux_v I__2815 (
            .O(N__11654),
            .I(N__11640));
    Span4Mux_v I__2814 (
            .O(N__11651),
            .I(N__11637));
    Sp12to4 I__2813 (
            .O(N__11648),
            .I(N__11630));
    Sp12to4 I__2812 (
            .O(N__11643),
            .I(N__11630));
    Sp12to4 I__2811 (
            .O(N__11640),
            .I(N__11630));
    Span4Mux_v I__2810 (
            .O(N__11637),
            .I(N__11627));
    Span12Mux_h I__2809 (
            .O(N__11630),
            .I(N__11622));
    Sp12to4 I__2808 (
            .O(N__11627),
            .I(N__11622));
    Odrv12 I__2807 (
            .O(N__11622),
            .I(A_c_1));
    CascadeMux I__2806 (
            .O(N__11619),
            .I(N__11613));
    InMux I__2805 (
            .O(N__11618),
            .I(N__11609));
    CascadeMux I__2804 (
            .O(N__11617),
            .I(N__11604));
    InMux I__2803 (
            .O(N__11616),
            .I(N__11598));
    InMux I__2802 (
            .O(N__11613),
            .I(N__11595));
    InMux I__2801 (
            .O(N__11612),
            .I(N__11592));
    LocalMux I__2800 (
            .O(N__11609),
            .I(N__11589));
    InMux I__2799 (
            .O(N__11608),
            .I(N__11584));
    InMux I__2798 (
            .O(N__11607),
            .I(N__11584));
    InMux I__2797 (
            .O(N__11604),
            .I(N__11581));
    InMux I__2796 (
            .O(N__11603),
            .I(N__11578));
    InMux I__2795 (
            .O(N__11602),
            .I(N__11575));
    CascadeMux I__2794 (
            .O(N__11601),
            .I(N__11572));
    LocalMux I__2793 (
            .O(N__11598),
            .I(N__11567));
    LocalMux I__2792 (
            .O(N__11595),
            .I(N__11567));
    LocalMux I__2791 (
            .O(N__11592),
            .I(N__11564));
    Span4Mux_h I__2790 (
            .O(N__11589),
            .I(N__11557));
    LocalMux I__2789 (
            .O(N__11584),
            .I(N__11557));
    LocalMux I__2788 (
            .O(N__11581),
            .I(N__11557));
    LocalMux I__2787 (
            .O(N__11578),
            .I(N__11552));
    LocalMux I__2786 (
            .O(N__11575),
            .I(N__11552));
    InMux I__2785 (
            .O(N__11572),
            .I(N__11549));
    Span4Mux_v I__2784 (
            .O(N__11567),
            .I(N__11546));
    Span4Mux_v I__2783 (
            .O(N__11564),
            .I(N__11543));
    Span4Mux_v I__2782 (
            .O(N__11557),
            .I(N__11538));
    Span4Mux_v I__2781 (
            .O(N__11552),
            .I(N__11538));
    LocalMux I__2780 (
            .O(N__11549),
            .I(N__11535));
    Sp12to4 I__2779 (
            .O(N__11546),
            .I(N__11528));
    Sp12to4 I__2778 (
            .O(N__11543),
            .I(N__11528));
    Sp12to4 I__2777 (
            .O(N__11538),
            .I(N__11528));
    Span4Mux_v I__2776 (
            .O(N__11535),
            .I(N__11525));
    Span12Mux_h I__2775 (
            .O(N__11528),
            .I(N__11520));
    Sp12to4 I__2774 (
            .O(N__11525),
            .I(N__11520));
    Odrv12 I__2773 (
            .O(N__11520),
            .I(A_c_0));
    InMux I__2772 (
            .O(N__11517),
            .I(N__11512));
    CascadeMux I__2771 (
            .O(N__11516),
            .I(N__11509));
    InMux I__2770 (
            .O(N__11515),
            .I(N__11506));
    LocalMux I__2769 (
            .O(N__11512),
            .I(N__11503));
    InMux I__2768 (
            .O(N__11509),
            .I(N__11500));
    LocalMux I__2767 (
            .O(N__11506),
            .I(N__11494));
    Span4Mux_v I__2766 (
            .O(N__11503),
            .I(N__11491));
    LocalMux I__2765 (
            .O(N__11500),
            .I(N__11488));
    InMux I__2764 (
            .O(N__11499),
            .I(N__11483));
    InMux I__2763 (
            .O(N__11498),
            .I(N__11483));
    InMux I__2762 (
            .O(N__11497),
            .I(N__11478));
    Span4Mux_v I__2761 (
            .O(N__11494),
            .I(N__11475));
    Span4Mux_v I__2760 (
            .O(N__11491),
            .I(N__11468));
    Span4Mux_h I__2759 (
            .O(N__11488),
            .I(N__11468));
    LocalMux I__2758 (
            .O(N__11483),
            .I(N__11468));
    InMux I__2757 (
            .O(N__11482),
            .I(N__11461));
    InMux I__2756 (
            .O(N__11481),
            .I(N__11461));
    LocalMux I__2755 (
            .O(N__11478),
            .I(N__11458));
    Span4Mux_v I__2754 (
            .O(N__11475),
            .I(N__11455));
    Span4Mux_h I__2753 (
            .O(N__11468),
            .I(N__11452));
    InMux I__2752 (
            .O(N__11467),
            .I(N__11449));
    InMux I__2751 (
            .O(N__11466),
            .I(N__11446));
    LocalMux I__2750 (
            .O(N__11461),
            .I(N__11443));
    Sp12to4 I__2749 (
            .O(N__11458),
            .I(N__11440));
    Span4Mux_v I__2748 (
            .O(N__11455),
            .I(N__11437));
    Span4Mux_v I__2747 (
            .O(N__11452),
            .I(N__11434));
    LocalMux I__2746 (
            .O(N__11449),
            .I(N__11429));
    LocalMux I__2745 (
            .O(N__11446),
            .I(N__11429));
    Span12Mux_v I__2744 (
            .O(N__11443),
            .I(N__11426));
    Span12Mux_v I__2743 (
            .O(N__11440),
            .I(N__11423));
    Sp12to4 I__2742 (
            .O(N__11437),
            .I(N__11416));
    Sp12to4 I__2741 (
            .O(N__11434),
            .I(N__11416));
    Span12Mux_v I__2740 (
            .O(N__11429),
            .I(N__11416));
    Span12Mux_h I__2739 (
            .O(N__11426),
            .I(N__11413));
    Span12Mux_h I__2738 (
            .O(N__11423),
            .I(N__11410));
    Span12Mux_h I__2737 (
            .O(N__11416),
            .I(N__11407));
    Odrv12 I__2736 (
            .O(N__11413),
            .I(SIZ_c_1));
    Odrv12 I__2735 (
            .O(N__11410),
            .I(SIZ_c_1));
    Odrv12 I__2734 (
            .O(N__11407),
            .I(SIZ_c_1));
    CascadeMux I__2733 (
            .O(N__11400),
            .I(N__11394));
    InMux I__2732 (
            .O(N__11399),
            .I(N__11391));
    InMux I__2731 (
            .O(N__11398),
            .I(N__11388));
    InMux I__2730 (
            .O(N__11397),
            .I(N__11385));
    InMux I__2729 (
            .O(N__11394),
            .I(N__11382));
    LocalMux I__2728 (
            .O(N__11391),
            .I(N__11374));
    LocalMux I__2727 (
            .O(N__11388),
            .I(N__11374));
    LocalMux I__2726 (
            .O(N__11385),
            .I(N__11369));
    LocalMux I__2725 (
            .O(N__11382),
            .I(N__11369));
    CascadeMux I__2724 (
            .O(N__11381),
            .I(N__11365));
    CascadeMux I__2723 (
            .O(N__11380),
            .I(N__11362));
    CascadeMux I__2722 (
            .O(N__11379),
            .I(N__11359));
    Span4Mux_v I__2721 (
            .O(N__11374),
            .I(N__11355));
    Span4Mux_v I__2720 (
            .O(N__11369),
            .I(N__11352));
    InMux I__2719 (
            .O(N__11368),
            .I(N__11349));
    InMux I__2718 (
            .O(N__11365),
            .I(N__11344));
    InMux I__2717 (
            .O(N__11362),
            .I(N__11344));
    InMux I__2716 (
            .O(N__11359),
            .I(N__11340));
    InMux I__2715 (
            .O(N__11358),
            .I(N__11337));
    Span4Mux_v I__2714 (
            .O(N__11355),
            .I(N__11328));
    Span4Mux_v I__2713 (
            .O(N__11352),
            .I(N__11328));
    LocalMux I__2712 (
            .O(N__11349),
            .I(N__11328));
    LocalMux I__2711 (
            .O(N__11344),
            .I(N__11328));
    InMux I__2710 (
            .O(N__11343),
            .I(N__11325));
    LocalMux I__2709 (
            .O(N__11340),
            .I(N__11322));
    LocalMux I__2708 (
            .O(N__11337),
            .I(N__11319));
    Span4Mux_h I__2707 (
            .O(N__11328),
            .I(N__11314));
    LocalMux I__2706 (
            .O(N__11325),
            .I(N__11314));
    Span4Mux_v I__2705 (
            .O(N__11322),
            .I(N__11311));
    Span4Mux_v I__2704 (
            .O(N__11319),
            .I(N__11308));
    Span4Mux_h I__2703 (
            .O(N__11314),
            .I(N__11305));
    Sp12to4 I__2702 (
            .O(N__11311),
            .I(N__11302));
    Span4Mux_v I__2701 (
            .O(N__11308),
            .I(N__11299));
    Span4Mux_v I__2700 (
            .O(N__11305),
            .I(N__11296));
    Span12Mux_h I__2699 (
            .O(N__11302),
            .I(N__11293));
    Span4Mux_v I__2698 (
            .O(N__11299),
            .I(N__11290));
    Span4Mux_h I__2697 (
            .O(N__11296),
            .I(N__11287));
    Span12Mux_v I__2696 (
            .O(N__11293),
            .I(N__11284));
    Sp12to4 I__2695 (
            .O(N__11290),
            .I(N__11279));
    Sp12to4 I__2694 (
            .O(N__11287),
            .I(N__11279));
    Odrv12 I__2693 (
            .O(N__11284),
            .I(SIZ_c_0));
    Odrv12 I__2692 (
            .O(N__11279),
            .I(SIZ_c_0));
    IoInMux I__2691 (
            .O(N__11274),
            .I(N__11271));
    LocalMux I__2690 (
            .O(N__11271),
            .I(N__11268));
    Span4Mux_s2_v I__2689 (
            .O(N__11268),
            .I(N__11265));
    Span4Mux_v I__2688 (
            .O(N__11265),
            .I(N__11262));
    Odrv4 I__2687 (
            .O(N__11262),
            .I(N_334_i));
    CascadeMux I__2686 (
            .O(N__11259),
            .I(N__11254));
    InMux I__2685 (
            .O(N__11258),
            .I(N__11251));
    InMux I__2684 (
            .O(N__11257),
            .I(N__11247));
    InMux I__2683 (
            .O(N__11254),
            .I(N__11244));
    LocalMux I__2682 (
            .O(N__11251),
            .I(N__11241));
    InMux I__2681 (
            .O(N__11250),
            .I(N__11238));
    LocalMux I__2680 (
            .O(N__11247),
            .I(N__11235));
    LocalMux I__2679 (
            .O(N__11244),
            .I(N__11231));
    Span4Mux_v I__2678 (
            .O(N__11241),
            .I(N__11228));
    LocalMux I__2677 (
            .O(N__11238),
            .I(N__11225));
    Span4Mux_v I__2676 (
            .O(N__11235),
            .I(N__11222));
    InMux I__2675 (
            .O(N__11234),
            .I(N__11219));
    Span4Mux_v I__2674 (
            .O(N__11231),
            .I(N__11216));
    Span4Mux_v I__2673 (
            .O(N__11228),
            .I(N__11213));
    Span4Mux_v I__2672 (
            .O(N__11225),
            .I(N__11210));
    Sp12to4 I__2671 (
            .O(N__11222),
            .I(N__11207));
    LocalMux I__2670 (
            .O(N__11219),
            .I(N__11204));
    Span4Mux_h I__2669 (
            .O(N__11216),
            .I(N__11201));
    Span4Mux_v I__2668 (
            .O(N__11213),
            .I(N__11196));
    Span4Mux_h I__2667 (
            .O(N__11210),
            .I(N__11196));
    Span12Mux_h I__2666 (
            .O(N__11207),
            .I(N__11191));
    Span12Mux_v I__2665 (
            .O(N__11204),
            .I(N__11191));
    Sp12to4 I__2664 (
            .O(N__11201),
            .I(N__11186));
    Sp12to4 I__2663 (
            .O(N__11196),
            .I(N__11186));
    Span12Mux_h I__2662 (
            .O(N__11191),
            .I(N__11183));
    Span12Mux_h I__2661 (
            .O(N__11186),
            .I(N__11180));
    Odrv12 I__2660 (
            .O(N__11183),
            .I(RnW_c));
    Odrv12 I__2659 (
            .O(N__11180),
            .I(RnW_c));
    InMux I__2658 (
            .O(N__11175),
            .I(N__11171));
    InMux I__2657 (
            .O(N__11174),
            .I(N__11168));
    LocalMux I__2656 (
            .O(N__11171),
            .I(N__11165));
    LocalMux I__2655 (
            .O(N__11168),
            .I(N__11162));
    Span12Mux_s6_h I__2654 (
            .O(N__11165),
            .I(N__11159));
    Sp12to4 I__2653 (
            .O(N__11162),
            .I(N__11156));
    Span12Mux_v I__2652 (
            .O(N__11159),
            .I(N__11150));
    Span12Mux_v I__2651 (
            .O(N__11156),
            .I(N__11150));
    InMux I__2650 (
            .O(N__11155),
            .I(N__11147));
    Odrv12 I__2649 (
            .O(N__11150),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2648 (
            .O(N__11147),
            .I(DMA_WRITE_CYCLE));
    IoInMux I__2647 (
            .O(N__11142),
            .I(N__11139));
    LocalMux I__2646 (
            .O(N__11139),
            .I(N__11136));
    IoSpan4Mux I__2645 (
            .O(N__11136),
            .I(N__11133));
    Span4Mux_s3_h I__2644 (
            .O(N__11133),
            .I(N__11130));
    Odrv4 I__2643 (
            .O(N__11130),
            .I(N_379));
    InMux I__2642 (
            .O(N__11127),
            .I(N__11124));
    LocalMux I__2641 (
            .O(N__11124),
            .I(N__11117));
    InMux I__2640 (
            .O(N__11123),
            .I(N__11114));
    InMux I__2639 (
            .O(N__11122),
            .I(N__11111));
    InMux I__2638 (
            .O(N__11121),
            .I(N__11105));
    InMux I__2637 (
            .O(N__11120),
            .I(N__11105));
    Sp12to4 I__2636 (
            .O(N__11117),
            .I(N__11102));
    LocalMux I__2635 (
            .O(N__11114),
            .I(N__11099));
    LocalMux I__2634 (
            .O(N__11111),
            .I(N__11096));
    InMux I__2633 (
            .O(N__11110),
            .I(N__11093));
    LocalMux I__2632 (
            .O(N__11105),
            .I(N__11090));
    Span12Mux_v I__2631 (
            .O(N__11102),
            .I(N__11087));
    Span12Mux_h I__2630 (
            .O(N__11099),
            .I(N__11084));
    Span12Mux_h I__2629 (
            .O(N__11096),
            .I(N__11079));
    LocalMux I__2628 (
            .O(N__11093),
            .I(N__11079));
    Span4Mux_h I__2627 (
            .O(N__11090),
            .I(N__11076));
    Span12Mux_h I__2626 (
            .O(N__11087),
            .I(N__11073));
    Span12Mux_v I__2625 (
            .O(N__11084),
            .I(N__11070));
    Span12Mux_v I__2624 (
            .O(N__11079),
            .I(N__11067));
    Span4Mux_v I__2623 (
            .O(N__11076),
            .I(N__11064));
    Odrv12 I__2622 (
            .O(N__11073),
            .I(CASUn_c));
    Odrv12 I__2621 (
            .O(N__11070),
            .I(CASUn_c));
    Odrv12 I__2620 (
            .O(N__11067),
            .I(CASUn_c));
    Odrv4 I__2619 (
            .O(N__11064),
            .I(CASUn_c));
    InMux I__2618 (
            .O(N__11055),
            .I(N__11052));
    LocalMux I__2617 (
            .O(N__11052),
            .I(N__11048));
    InMux I__2616 (
            .O(N__11051),
            .I(N__11045));
    Span4Mux_v I__2615 (
            .O(N__11048),
            .I(N__11040));
    LocalMux I__2614 (
            .O(N__11045),
            .I(N__11037));
    InMux I__2613 (
            .O(N__11044),
            .I(N__11034));
    InMux I__2612 (
            .O(N__11043),
            .I(N__11031));
    Span4Mux_v I__2611 (
            .O(N__11040),
            .I(N__11024));
    Span4Mux_v I__2610 (
            .O(N__11037),
            .I(N__11024));
    LocalMux I__2609 (
            .O(N__11034),
            .I(N__11024));
    LocalMux I__2608 (
            .O(N__11031),
            .I(N__11021));
    Span4Mux_v I__2607 (
            .O(N__11024),
            .I(N__11017));
    Span4Mux_v I__2606 (
            .O(N__11021),
            .I(N__11014));
    CascadeMux I__2605 (
            .O(N__11020),
            .I(N__11010));
    Span4Mux_v I__2604 (
            .O(N__11017),
            .I(N__11007));
    Sp12to4 I__2603 (
            .O(N__11014),
            .I(N__11004));
    InMux I__2602 (
            .O(N__11013),
            .I(N__11001));
    InMux I__2601 (
            .O(N__11010),
            .I(N__10998));
    Sp12to4 I__2600 (
            .O(N__11007),
            .I(N__10995));
    Span12Mux_h I__2599 (
            .O(N__11004),
            .I(N__10988));
    LocalMux I__2598 (
            .O(N__11001),
            .I(N__10988));
    LocalMux I__2597 (
            .O(N__10998),
            .I(N__10988));
    Span12Mux_h I__2596 (
            .O(N__10995),
            .I(N__10985));
    Span12Mux_v I__2595 (
            .O(N__10988),
            .I(N__10982));
    Odrv12 I__2594 (
            .O(N__10985),
            .I(CASLn_c));
    Odrv12 I__2593 (
            .O(N__10982),
            .I(CASLn_c));
    CascadeMux I__2592 (
            .O(N__10977),
            .I(N__10974));
    InMux I__2591 (
            .O(N__10974),
            .I(N__10970));
    InMux I__2590 (
            .O(N__10973),
            .I(N__10967));
    LocalMux I__2589 (
            .O(N__10970),
            .I(N__10962));
    LocalMux I__2588 (
            .O(N__10967),
            .I(N__10959));
    InMux I__2587 (
            .O(N__10966),
            .I(N__10956));
    InMux I__2586 (
            .O(N__10965),
            .I(N__10953));
    Span4Mux_v I__2585 (
            .O(N__10962),
            .I(N__10941));
    Span4Mux_v I__2584 (
            .O(N__10959),
            .I(N__10936));
    LocalMux I__2583 (
            .O(N__10956),
            .I(N__10936));
    LocalMux I__2582 (
            .O(N__10953),
            .I(N__10933));
    InMux I__2581 (
            .O(N__10952),
            .I(N__10929));
    InMux I__2580 (
            .O(N__10951),
            .I(N__10922));
    InMux I__2579 (
            .O(N__10950),
            .I(N__10922));
    InMux I__2578 (
            .O(N__10949),
            .I(N__10922));
    InMux I__2577 (
            .O(N__10948),
            .I(N__10917));
    InMux I__2576 (
            .O(N__10947),
            .I(N__10917));
    InMux I__2575 (
            .O(N__10946),
            .I(N__10914));
    CascadeMux I__2574 (
            .O(N__10945),
            .I(N__10911));
    InMux I__2573 (
            .O(N__10944),
            .I(N__10906));
    Sp12to4 I__2572 (
            .O(N__10941),
            .I(N__10903));
    Span4Mux_v I__2571 (
            .O(N__10936),
            .I(N__10900));
    Span4Mux_v I__2570 (
            .O(N__10933),
            .I(N__10897));
    InMux I__2569 (
            .O(N__10932),
            .I(N__10893));
    LocalMux I__2568 (
            .O(N__10929),
            .I(N__10883));
    LocalMux I__2567 (
            .O(N__10922),
            .I(N__10878));
    LocalMux I__2566 (
            .O(N__10917),
            .I(N__10878));
    LocalMux I__2565 (
            .O(N__10914),
            .I(N__10875));
    InMux I__2564 (
            .O(N__10911),
            .I(N__10872));
    InMux I__2563 (
            .O(N__10910),
            .I(N__10867));
    InMux I__2562 (
            .O(N__10909),
            .I(N__10867));
    LocalMux I__2561 (
            .O(N__10906),
            .I(N__10864));
    Span12Mux_h I__2560 (
            .O(N__10903),
            .I(N__10861));
    Span4Mux_h I__2559 (
            .O(N__10900),
            .I(N__10858));
    Span4Mux_h I__2558 (
            .O(N__10897),
            .I(N__10855));
    InMux I__2557 (
            .O(N__10896),
            .I(N__10852));
    LocalMux I__2556 (
            .O(N__10893),
            .I(N__10849));
    InMux I__2555 (
            .O(N__10892),
            .I(N__10844));
    InMux I__2554 (
            .O(N__10891),
            .I(N__10844));
    InMux I__2553 (
            .O(N__10890),
            .I(N__10841));
    InMux I__2552 (
            .O(N__10889),
            .I(N__10832));
    InMux I__2551 (
            .O(N__10888),
            .I(N__10832));
    InMux I__2550 (
            .O(N__10887),
            .I(N__10832));
    InMux I__2549 (
            .O(N__10886),
            .I(N__10832));
    Span4Mux_v I__2548 (
            .O(N__10883),
            .I(N__10825));
    Span4Mux_v I__2547 (
            .O(N__10878),
            .I(N__10825));
    Span4Mux_h I__2546 (
            .O(N__10875),
            .I(N__10825));
    LocalMux I__2545 (
            .O(N__10872),
            .I(N__10818));
    LocalMux I__2544 (
            .O(N__10867),
            .I(N__10818));
    Span4Mux_h I__2543 (
            .O(N__10864),
            .I(N__10818));
    Odrv12 I__2542 (
            .O(N__10861),
            .I(CPU_CYCLEm));
    Odrv4 I__2541 (
            .O(N__10858),
            .I(CPU_CYCLEm));
    Odrv4 I__2540 (
            .O(N__10855),
            .I(CPU_CYCLEm));
    LocalMux I__2539 (
            .O(N__10852),
            .I(CPU_CYCLEm));
    Odrv4 I__2538 (
            .O(N__10849),
            .I(CPU_CYCLEm));
    LocalMux I__2537 (
            .O(N__10844),
            .I(CPU_CYCLEm));
    LocalMux I__2536 (
            .O(N__10841),
            .I(CPU_CYCLEm));
    LocalMux I__2535 (
            .O(N__10832),
            .I(CPU_CYCLEm));
    Odrv4 I__2534 (
            .O(N__10825),
            .I(CPU_CYCLEm));
    Odrv4 I__2533 (
            .O(N__10818),
            .I(CPU_CYCLEm));
    InMux I__2532 (
            .O(N__10797),
            .I(N__10792));
    InMux I__2531 (
            .O(N__10796),
            .I(N__10789));
    InMux I__2530 (
            .O(N__10795),
            .I(N__10786));
    LocalMux I__2529 (
            .O(N__10792),
            .I(N__10782));
    LocalMux I__2528 (
            .O(N__10789),
            .I(N__10777));
    LocalMux I__2527 (
            .O(N__10786),
            .I(N__10777));
    InMux I__2526 (
            .O(N__10785),
            .I(N__10774));
    Span4Mux_h I__2525 (
            .O(N__10782),
            .I(N__10771));
    Span4Mux_v I__2524 (
            .O(N__10777),
            .I(N__10766));
    LocalMux I__2523 (
            .O(N__10774),
            .I(N__10766));
    Sp12to4 I__2522 (
            .O(N__10771),
            .I(N__10763));
    Span4Mux_h I__2521 (
            .O(N__10766),
            .I(N__10760));
    Span12Mux_v I__2520 (
            .O(N__10763),
            .I(N__10757));
    Sp12to4 I__2519 (
            .O(N__10760),
            .I(N__10754));
    Span12Mux_h I__2518 (
            .O(N__10757),
            .I(N__10751));
    Span12Mux_v I__2517 (
            .O(N__10754),
            .I(N__10748));
    Odrv12 I__2516 (
            .O(N__10751),
            .I(DRA_c_5));
    Odrv12 I__2515 (
            .O(N__10748),
            .I(DRA_c_5));
    CascadeMux I__2514 (
            .O(N__10743),
            .I(N__10738));
    CascadeMux I__2513 (
            .O(N__10742),
            .I(N__10730));
    InMux I__2512 (
            .O(N__10741),
            .I(N__10726));
    InMux I__2511 (
            .O(N__10738),
            .I(N__10723));
    CascadeMux I__2510 (
            .O(N__10737),
            .I(N__10717));
    InMux I__2509 (
            .O(N__10736),
            .I(N__10709));
    InMux I__2508 (
            .O(N__10735),
            .I(N__10706));
    InMux I__2507 (
            .O(N__10734),
            .I(N__10703));
    InMux I__2506 (
            .O(N__10733),
            .I(N__10698));
    InMux I__2505 (
            .O(N__10730),
            .I(N__10693));
    InMux I__2504 (
            .O(N__10729),
            .I(N__10693));
    LocalMux I__2503 (
            .O(N__10726),
            .I(N__10690));
    LocalMux I__2502 (
            .O(N__10723),
            .I(N__10687));
    InMux I__2501 (
            .O(N__10722),
            .I(N__10682));
    InMux I__2500 (
            .O(N__10721),
            .I(N__10682));
    InMux I__2499 (
            .O(N__10720),
            .I(N__10679));
    InMux I__2498 (
            .O(N__10717),
            .I(N__10672));
    InMux I__2497 (
            .O(N__10716),
            .I(N__10672));
    InMux I__2496 (
            .O(N__10715),
            .I(N__10672));
    InMux I__2495 (
            .O(N__10714),
            .I(N__10669));
    InMux I__2494 (
            .O(N__10713),
            .I(N__10666));
    InMux I__2493 (
            .O(N__10712),
            .I(N__10662));
    LocalMux I__2492 (
            .O(N__10709),
            .I(N__10659));
    LocalMux I__2491 (
            .O(N__10706),
            .I(N__10654));
    LocalMux I__2490 (
            .O(N__10703),
            .I(N__10654));
    InMux I__2489 (
            .O(N__10702),
            .I(N__10651));
    InMux I__2488 (
            .O(N__10701),
            .I(N__10648));
    LocalMux I__2487 (
            .O(N__10698),
            .I(N__10643));
    LocalMux I__2486 (
            .O(N__10693),
            .I(N__10643));
    Span4Mux_v I__2485 (
            .O(N__10690),
            .I(N__10631));
    Span4Mux_v I__2484 (
            .O(N__10687),
            .I(N__10631));
    LocalMux I__2483 (
            .O(N__10682),
            .I(N__10631));
    LocalMux I__2482 (
            .O(N__10679),
            .I(N__10631));
    LocalMux I__2481 (
            .O(N__10672),
            .I(N__10631));
    LocalMux I__2480 (
            .O(N__10669),
            .I(N__10626));
    LocalMux I__2479 (
            .O(N__10666),
            .I(N__10626));
    InMux I__2478 (
            .O(N__10665),
            .I(N__10623));
    LocalMux I__2477 (
            .O(N__10662),
            .I(N__10620));
    Span4Mux_h I__2476 (
            .O(N__10659),
            .I(N__10617));
    Span4Mux_v I__2475 (
            .O(N__10654),
            .I(N__10610));
    LocalMux I__2474 (
            .O(N__10651),
            .I(N__10610));
    LocalMux I__2473 (
            .O(N__10648),
            .I(N__10610));
    Span4Mux_v I__2472 (
            .O(N__10643),
            .I(N__10607));
    InMux I__2471 (
            .O(N__10642),
            .I(N__10604));
    Span4Mux_h I__2470 (
            .O(N__10631),
            .I(N__10595));
    Span4Mux_v I__2469 (
            .O(N__10626),
            .I(N__10595));
    LocalMux I__2468 (
            .O(N__10623),
            .I(N__10595));
    Span4Mux_v I__2467 (
            .O(N__10620),
            .I(N__10595));
    Sp12to4 I__2466 (
            .O(N__10617),
            .I(N__10592));
    Sp12to4 I__2465 (
            .O(N__10610),
            .I(N__10589));
    Sp12to4 I__2464 (
            .O(N__10607),
            .I(N__10582));
    LocalMux I__2463 (
            .O(N__10604),
            .I(N__10582));
    Sp12to4 I__2462 (
            .O(N__10595),
            .I(N__10582));
    Span12Mux_v I__2461 (
            .O(N__10592),
            .I(N__10579));
    Span12Mux_v I__2460 (
            .O(N__10589),
            .I(N__10576));
    Span12Mux_h I__2459 (
            .O(N__10582),
            .I(N__10573));
    Span12Mux_h I__2458 (
            .O(N__10579),
            .I(N__10570));
    Span12Mux_h I__2457 (
            .O(N__10576),
            .I(N__10565));
    Span12Mux_v I__2456 (
            .O(N__10573),
            .I(N__10565));
    Odrv12 I__2455 (
            .O(N__10570),
            .I(AGNUS_REV_c));
    Odrv12 I__2454 (
            .O(N__10565),
            .I(AGNUS_REV_c));
    InMux I__2453 (
            .O(N__10560),
            .I(N__10554));
    InMux I__2452 (
            .O(N__10559),
            .I(N__10551));
    InMux I__2451 (
            .O(N__10558),
            .I(N__10546));
    InMux I__2450 (
            .O(N__10557),
            .I(N__10546));
    LocalMux I__2449 (
            .O(N__10554),
            .I(N__10543));
    LocalMux I__2448 (
            .O(N__10551),
            .I(N__10540));
    LocalMux I__2447 (
            .O(N__10546),
            .I(N__10537));
    Span4Mux_h I__2446 (
            .O(N__10543),
            .I(N__10532));
    Span4Mux_v I__2445 (
            .O(N__10540),
            .I(N__10532));
    Sp12to4 I__2444 (
            .O(N__10537),
            .I(N__10529));
    Span4Mux_v I__2443 (
            .O(N__10532),
            .I(N__10526));
    Span12Mux_v I__2442 (
            .O(N__10529),
            .I(N__10521));
    Sp12to4 I__2441 (
            .O(N__10526),
            .I(N__10521));
    Span12Mux_h I__2440 (
            .O(N__10521),
            .I(N__10518));
    Odrv12 I__2439 (
            .O(N__10518),
            .I(DRA_c_6));
    InMux I__2438 (
            .O(N__10515),
            .I(N__10512));
    LocalMux I__2437 (
            .O(N__10512),
            .I(N__10509));
    Odrv12 I__2436 (
            .O(N__10509),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    CEMux I__2435 (
            .O(N__10506),
            .I(N__10464));
    CEMux I__2434 (
            .O(N__10505),
            .I(N__10464));
    CEMux I__2433 (
            .O(N__10504),
            .I(N__10464));
    CEMux I__2432 (
            .O(N__10503),
            .I(N__10464));
    CEMux I__2431 (
            .O(N__10502),
            .I(N__10464));
    CEMux I__2430 (
            .O(N__10501),
            .I(N__10464));
    CEMux I__2429 (
            .O(N__10500),
            .I(N__10464));
    CEMux I__2428 (
            .O(N__10499),
            .I(N__10464));
    CEMux I__2427 (
            .O(N__10498),
            .I(N__10464));
    CEMux I__2426 (
            .O(N__10497),
            .I(N__10464));
    CEMux I__2425 (
            .O(N__10496),
            .I(N__10464));
    CEMux I__2424 (
            .O(N__10495),
            .I(N__10464));
    CEMux I__2423 (
            .O(N__10494),
            .I(N__10464));
    CEMux I__2422 (
            .O(N__10493),
            .I(N__10464));
    GlobalMux I__2421 (
            .O(N__10464),
            .I(N__10461));
    gio2CtrlBuf I__2420 (
            .O(N__10461),
            .I(DBRn_c_i_0_g));
    InMux I__2419 (
            .O(N__10458),
            .I(N__10455));
    LocalMux I__2418 (
            .O(N__10455),
            .I(N__10452));
    Span12Mux_h I__2417 (
            .O(N__10452),
            .I(N__10449));
    Odrv12 I__2416 (
            .O(N__10449),
            .I(RAS1n_c));
    InMux I__2415 (
            .O(N__10446),
            .I(N__10442));
    InMux I__2414 (
            .O(N__10445),
            .I(N__10439));
    LocalMux I__2413 (
            .O(N__10442),
            .I(N__10436));
    LocalMux I__2412 (
            .O(N__10439),
            .I(N__10433));
    Span4Mux_v I__2411 (
            .O(N__10436),
            .I(N__10428));
    Span4Mux_v I__2410 (
            .O(N__10433),
            .I(N__10428));
    Sp12to4 I__2409 (
            .O(N__10428),
            .I(N__10425));
    Span12Mux_h I__2408 (
            .O(N__10425),
            .I(N__10422));
    Odrv12 I__2407 (
            .O(N__10422),
            .I(RAS0n_c));
    CascadeMux I__2406 (
            .O(N__10419),
            .I(N__10414));
    CascadeMux I__2405 (
            .O(N__10418),
            .I(N__10411));
    CascadeMux I__2404 (
            .O(N__10417),
            .I(N__10401));
    InMux I__2403 (
            .O(N__10414),
            .I(N__10397));
    InMux I__2402 (
            .O(N__10411),
            .I(N__10386));
    InMux I__2401 (
            .O(N__10410),
            .I(N__10386));
    InMux I__2400 (
            .O(N__10409),
            .I(N__10386));
    InMux I__2399 (
            .O(N__10408),
            .I(N__10375));
    InMux I__2398 (
            .O(N__10407),
            .I(N__10375));
    CascadeMux I__2397 (
            .O(N__10406),
            .I(N__10372));
    InMux I__2396 (
            .O(N__10405),
            .I(N__10367));
    InMux I__2395 (
            .O(N__10404),
            .I(N__10367));
    InMux I__2394 (
            .O(N__10401),
            .I(N__10364));
    InMux I__2393 (
            .O(N__10400),
            .I(N__10361));
    LocalMux I__2392 (
            .O(N__10397),
            .I(N__10358));
    InMux I__2391 (
            .O(N__10396),
            .I(N__10351));
    InMux I__2390 (
            .O(N__10395),
            .I(N__10351));
    InMux I__2389 (
            .O(N__10394),
            .I(N__10351));
    InMux I__2388 (
            .O(N__10393),
            .I(N__10347));
    LocalMux I__2387 (
            .O(N__10386),
            .I(N__10344));
    InMux I__2386 (
            .O(N__10385),
            .I(N__10341));
    InMux I__2385 (
            .O(N__10384),
            .I(N__10338));
    InMux I__2384 (
            .O(N__10383),
            .I(N__10335));
    InMux I__2383 (
            .O(N__10382),
            .I(N__10328));
    InMux I__2382 (
            .O(N__10381),
            .I(N__10328));
    InMux I__2381 (
            .O(N__10380),
            .I(N__10328));
    LocalMux I__2380 (
            .O(N__10375),
            .I(N__10322));
    InMux I__2379 (
            .O(N__10372),
            .I(N__10319));
    LocalMux I__2378 (
            .O(N__10367),
            .I(N__10312));
    LocalMux I__2377 (
            .O(N__10364),
            .I(N__10312));
    LocalMux I__2376 (
            .O(N__10361),
            .I(N__10309));
    Span4Mux_h I__2375 (
            .O(N__10358),
            .I(N__10304));
    LocalMux I__2374 (
            .O(N__10351),
            .I(N__10304));
    InMux I__2373 (
            .O(N__10350),
            .I(N__10301));
    LocalMux I__2372 (
            .O(N__10347),
            .I(N__10297));
    Span4Mux_v I__2371 (
            .O(N__10344),
            .I(N__10286));
    LocalMux I__2370 (
            .O(N__10341),
            .I(N__10286));
    LocalMux I__2369 (
            .O(N__10338),
            .I(N__10286));
    LocalMux I__2368 (
            .O(N__10335),
            .I(N__10286));
    LocalMux I__2367 (
            .O(N__10328),
            .I(N__10286));
    InMux I__2366 (
            .O(N__10327),
            .I(N__10283));
    InMux I__2365 (
            .O(N__10326),
            .I(N__10280));
    InMux I__2364 (
            .O(N__10325),
            .I(N__10277));
    Span4Mux_h I__2363 (
            .O(N__10322),
            .I(N__10272));
    LocalMux I__2362 (
            .O(N__10319),
            .I(N__10272));
    InMux I__2361 (
            .O(N__10318),
            .I(N__10269));
    InMux I__2360 (
            .O(N__10317),
            .I(N__10266));
    Span4Mux_h I__2359 (
            .O(N__10312),
            .I(N__10257));
    Span4Mux_v I__2358 (
            .O(N__10309),
            .I(N__10257));
    Span4Mux_v I__2357 (
            .O(N__10304),
            .I(N__10257));
    LocalMux I__2356 (
            .O(N__10301),
            .I(N__10257));
    InMux I__2355 (
            .O(N__10300),
            .I(N__10254));
    Span4Mux_v I__2354 (
            .O(N__10297),
            .I(N__10247));
    Span4Mux_v I__2353 (
            .O(N__10286),
            .I(N__10247));
    LocalMux I__2352 (
            .O(N__10283),
            .I(N__10240));
    LocalMux I__2351 (
            .O(N__10280),
            .I(N__10240));
    LocalMux I__2350 (
            .O(N__10277),
            .I(N__10240));
    Span4Mux_h I__2349 (
            .O(N__10272),
            .I(N__10233));
    LocalMux I__2348 (
            .O(N__10269),
            .I(N__10233));
    LocalMux I__2347 (
            .O(N__10266),
            .I(N__10233));
    Span4Mux_h I__2346 (
            .O(N__10257),
            .I(N__10226));
    LocalMux I__2345 (
            .O(N__10254),
            .I(N__10226));
    InMux I__2344 (
            .O(N__10253),
            .I(N__10221));
    InMux I__2343 (
            .O(N__10252),
            .I(N__10221));
    Span4Mux_h I__2342 (
            .O(N__10247),
            .I(N__10214));
    Span4Mux_v I__2341 (
            .O(N__10240),
            .I(N__10214));
    Span4Mux_v I__2340 (
            .O(N__10233),
            .I(N__10214));
    InMux I__2339 (
            .O(N__10232),
            .I(N__10209));
    InMux I__2338 (
            .O(N__10231),
            .I(N__10209));
    Sp12to4 I__2337 (
            .O(N__10226),
            .I(N__10206));
    LocalMux I__2336 (
            .O(N__10221),
            .I(N__10199));
    Sp12to4 I__2335 (
            .O(N__10214),
            .I(N__10199));
    LocalMux I__2334 (
            .O(N__10209),
            .I(N__10199));
    Span12Mux_v I__2333 (
            .O(N__10206),
            .I(N__10196));
    Span12Mux_h I__2332 (
            .O(N__10199),
            .I(N__10193));
    Span12Mux_h I__2331 (
            .O(N__10196),
            .I(N__10190));
    Odrv12 I__2330 (
            .O(N__10193),
            .I(RESETn_c));
    Odrv12 I__2329 (
            .O(N__10190),
            .I(RESETn_c));
    InMux I__2328 (
            .O(N__10185),
            .I(N__10182));
    LocalMux I__2327 (
            .O(N__10182),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2326 (
            .O(N__10179),
            .I(N__10176));
    LocalMux I__2325 (
            .O(N__10176),
            .I(N__10173));
    Odrv4 I__2324 (
            .O(N__10173),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    IoInMux I__2323 (
            .O(N__10170),
            .I(N__10167));
    LocalMux I__2322 (
            .O(N__10167),
            .I(N__10164));
    Span4Mux_s1_v I__2321 (
            .O(N__10164),
            .I(N__10161));
    Sp12to4 I__2320 (
            .O(N__10161),
            .I(N__10158));
    Span12Mux_h I__2319 (
            .O(N__10158),
            .I(N__10155));
    Span12Mux_v I__2318 (
            .O(N__10155),
            .I(N__10151));
    InMux I__2317 (
            .O(N__10154),
            .I(N__10148));
    Odrv12 I__2316 (
            .O(N__10151),
            .I(LDSn_c));
    LocalMux I__2315 (
            .O(N__10148),
            .I(LDSn_c));
    InMux I__2314 (
            .O(N__10143),
            .I(N__10140));
    LocalMux I__2313 (
            .O(N__10140),
            .I(\U712_REG_SM.N_459 ));
    CascadeMux I__2312 (
            .O(N__10137),
            .I(N__10133));
    InMux I__2311 (
            .O(N__10136),
            .I(N__10128));
    InMux I__2310 (
            .O(N__10133),
            .I(N__10128));
    LocalMux I__2309 (
            .O(N__10128),
            .I(N__10124));
    InMux I__2308 (
            .O(N__10127),
            .I(N__10121));
    Odrv12 I__2307 (
            .O(N__10124),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    LocalMux I__2306 (
            .O(N__10121),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    InMux I__2305 (
            .O(N__10116),
            .I(N__10110));
    InMux I__2304 (
            .O(N__10115),
            .I(N__10105));
    InMux I__2303 (
            .O(N__10114),
            .I(N__10105));
    CascadeMux I__2302 (
            .O(N__10113),
            .I(N__10093));
    LocalMux I__2301 (
            .O(N__10110),
            .I(N__10088));
    LocalMux I__2300 (
            .O(N__10105),
            .I(N__10088));
    CascadeMux I__2299 (
            .O(N__10104),
            .I(N__10085));
    InMux I__2298 (
            .O(N__10103),
            .I(N__10082));
    InMux I__2297 (
            .O(N__10102),
            .I(N__10079));
    InMux I__2296 (
            .O(N__10101),
            .I(N__10076));
    InMux I__2295 (
            .O(N__10100),
            .I(N__10071));
    InMux I__2294 (
            .O(N__10099),
            .I(N__10071));
    InMux I__2293 (
            .O(N__10098),
            .I(N__10066));
    InMux I__2292 (
            .O(N__10097),
            .I(N__10066));
    CascadeMux I__2291 (
            .O(N__10096),
            .I(N__10062));
    InMux I__2290 (
            .O(N__10093),
            .I(N__10059));
    Span4Mux_h I__2289 (
            .O(N__10088),
            .I(N__10056));
    InMux I__2288 (
            .O(N__10085),
            .I(N__10053));
    LocalMux I__2287 (
            .O(N__10082),
            .I(N__10044));
    LocalMux I__2286 (
            .O(N__10079),
            .I(N__10044));
    LocalMux I__2285 (
            .O(N__10076),
            .I(N__10044));
    LocalMux I__2284 (
            .O(N__10071),
            .I(N__10044));
    LocalMux I__2283 (
            .O(N__10066),
            .I(N__10041));
    InMux I__2282 (
            .O(N__10065),
            .I(N__10036));
    InMux I__2281 (
            .O(N__10062),
            .I(N__10036));
    LocalMux I__2280 (
            .O(N__10059),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2279 (
            .O(N__10056),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2278 (
            .O(N__10053),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2277 (
            .O(N__10044),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv12 I__2276 (
            .O(N__10041),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2275 (
            .O(N__10036),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__2274 (
            .O(N__10023),
            .I(N__10020));
    LocalMux I__2273 (
            .O(N__10020),
            .I(N__10017));
    IoSpan4Mux I__2272 (
            .O(N__10017),
            .I(N__10014));
    Span4Mux_s2_v I__2271 (
            .O(N__10014),
            .I(N__10011));
    Sp12to4 I__2270 (
            .O(N__10011),
            .I(N__10007));
    CascadeMux I__2269 (
            .O(N__10010),
            .I(N__10004));
    Span12Mux_v I__2268 (
            .O(N__10007),
            .I(N__10001));
    InMux I__2267 (
            .O(N__10004),
            .I(N__9998));
    Odrv12 I__2266 (
            .O(N__10001),
            .I(UDSn_c));
    LocalMux I__2265 (
            .O(N__9998),
            .I(UDSn_c));
    InMux I__2264 (
            .O(N__9993),
            .I(N__9990));
    LocalMux I__2263 (
            .O(N__9990),
            .I(N__9950));
    ClkMux I__2262 (
            .O(N__9989),
            .I(N__9831));
    ClkMux I__2261 (
            .O(N__9988),
            .I(N__9831));
    ClkMux I__2260 (
            .O(N__9987),
            .I(N__9831));
    ClkMux I__2259 (
            .O(N__9986),
            .I(N__9831));
    ClkMux I__2258 (
            .O(N__9985),
            .I(N__9831));
    ClkMux I__2257 (
            .O(N__9984),
            .I(N__9831));
    ClkMux I__2256 (
            .O(N__9983),
            .I(N__9831));
    ClkMux I__2255 (
            .O(N__9982),
            .I(N__9831));
    ClkMux I__2254 (
            .O(N__9981),
            .I(N__9831));
    ClkMux I__2253 (
            .O(N__9980),
            .I(N__9831));
    ClkMux I__2252 (
            .O(N__9979),
            .I(N__9831));
    ClkMux I__2251 (
            .O(N__9978),
            .I(N__9831));
    ClkMux I__2250 (
            .O(N__9977),
            .I(N__9831));
    ClkMux I__2249 (
            .O(N__9976),
            .I(N__9831));
    ClkMux I__2248 (
            .O(N__9975),
            .I(N__9831));
    ClkMux I__2247 (
            .O(N__9974),
            .I(N__9831));
    ClkMux I__2246 (
            .O(N__9973),
            .I(N__9831));
    ClkMux I__2245 (
            .O(N__9972),
            .I(N__9831));
    ClkMux I__2244 (
            .O(N__9971),
            .I(N__9831));
    ClkMux I__2243 (
            .O(N__9970),
            .I(N__9831));
    ClkMux I__2242 (
            .O(N__9969),
            .I(N__9831));
    ClkMux I__2241 (
            .O(N__9968),
            .I(N__9831));
    ClkMux I__2240 (
            .O(N__9967),
            .I(N__9831));
    ClkMux I__2239 (
            .O(N__9966),
            .I(N__9831));
    ClkMux I__2238 (
            .O(N__9965),
            .I(N__9831));
    ClkMux I__2237 (
            .O(N__9964),
            .I(N__9831));
    ClkMux I__2236 (
            .O(N__9963),
            .I(N__9831));
    ClkMux I__2235 (
            .O(N__9962),
            .I(N__9831));
    ClkMux I__2234 (
            .O(N__9961),
            .I(N__9831));
    ClkMux I__2233 (
            .O(N__9960),
            .I(N__9831));
    ClkMux I__2232 (
            .O(N__9959),
            .I(N__9831));
    ClkMux I__2231 (
            .O(N__9958),
            .I(N__9831));
    ClkMux I__2230 (
            .O(N__9957),
            .I(N__9831));
    ClkMux I__2229 (
            .O(N__9956),
            .I(N__9831));
    ClkMux I__2228 (
            .O(N__9955),
            .I(N__9831));
    ClkMux I__2227 (
            .O(N__9954),
            .I(N__9831));
    ClkMux I__2226 (
            .O(N__9953),
            .I(N__9831));
    Glb2LocalMux I__2225 (
            .O(N__9950),
            .I(N__9831));
    ClkMux I__2224 (
            .O(N__9949),
            .I(N__9831));
    ClkMux I__2223 (
            .O(N__9948),
            .I(N__9831));
    ClkMux I__2222 (
            .O(N__9947),
            .I(N__9831));
    ClkMux I__2221 (
            .O(N__9946),
            .I(N__9831));
    ClkMux I__2220 (
            .O(N__9945),
            .I(N__9831));
    ClkMux I__2219 (
            .O(N__9944),
            .I(N__9831));
    ClkMux I__2218 (
            .O(N__9943),
            .I(N__9831));
    ClkMux I__2217 (
            .O(N__9942),
            .I(N__9831));
    ClkMux I__2216 (
            .O(N__9941),
            .I(N__9831));
    ClkMux I__2215 (
            .O(N__9940),
            .I(N__9831));
    ClkMux I__2214 (
            .O(N__9939),
            .I(N__9831));
    ClkMux I__2213 (
            .O(N__9938),
            .I(N__9831));
    ClkMux I__2212 (
            .O(N__9937),
            .I(N__9831));
    ClkMux I__2211 (
            .O(N__9936),
            .I(N__9831));
    GlobalMux I__2210 (
            .O(N__9831),
            .I(CLK80_PLL));
    InMux I__2209 (
            .O(N__9828),
            .I(N__9820));
    InMux I__2208 (
            .O(N__9827),
            .I(N__9817));
    InMux I__2207 (
            .O(N__9826),
            .I(N__9814));
    InMux I__2206 (
            .O(N__9825),
            .I(N__9811));
    InMux I__2205 (
            .O(N__9824),
            .I(N__9808));
    InMux I__2204 (
            .O(N__9823),
            .I(N__9805));
    LocalMux I__2203 (
            .O(N__9820),
            .I(N__9802));
    LocalMux I__2202 (
            .O(N__9817),
            .I(N__9796));
    LocalMux I__2201 (
            .O(N__9814),
            .I(N__9788));
    LocalMux I__2200 (
            .O(N__9811),
            .I(N__9781));
    LocalMux I__2199 (
            .O(N__9808),
            .I(N__9770));
    LocalMux I__2198 (
            .O(N__9805),
            .I(N__9746));
    Glb2LocalMux I__2197 (
            .O(N__9802),
            .I(N__9642));
    SRMux I__2196 (
            .O(N__9801),
            .I(N__9642));
    SRMux I__2195 (
            .O(N__9800),
            .I(N__9642));
    SRMux I__2194 (
            .O(N__9799),
            .I(N__9642));
    Glb2LocalMux I__2193 (
            .O(N__9796),
            .I(N__9642));
    SRMux I__2192 (
            .O(N__9795),
            .I(N__9642));
    SRMux I__2191 (
            .O(N__9794),
            .I(N__9642));
    SRMux I__2190 (
            .O(N__9793),
            .I(N__9642));
    SRMux I__2189 (
            .O(N__9792),
            .I(N__9642));
    SRMux I__2188 (
            .O(N__9791),
            .I(N__9642));
    Glb2LocalMux I__2187 (
            .O(N__9788),
            .I(N__9642));
    SRMux I__2186 (
            .O(N__9787),
            .I(N__9642));
    SRMux I__2185 (
            .O(N__9786),
            .I(N__9642));
    SRMux I__2184 (
            .O(N__9785),
            .I(N__9642));
    SRMux I__2183 (
            .O(N__9784),
            .I(N__9642));
    Glb2LocalMux I__2182 (
            .O(N__9781),
            .I(N__9642));
    SRMux I__2181 (
            .O(N__9780),
            .I(N__9642));
    SRMux I__2180 (
            .O(N__9779),
            .I(N__9642));
    SRMux I__2179 (
            .O(N__9778),
            .I(N__9642));
    SRMux I__2178 (
            .O(N__9777),
            .I(N__9642));
    SRMux I__2177 (
            .O(N__9776),
            .I(N__9642));
    SRMux I__2176 (
            .O(N__9775),
            .I(N__9642));
    SRMux I__2175 (
            .O(N__9774),
            .I(N__9642));
    SRMux I__2174 (
            .O(N__9773),
            .I(N__9642));
    Glb2LocalMux I__2173 (
            .O(N__9770),
            .I(N__9642));
    SRMux I__2172 (
            .O(N__9769),
            .I(N__9642));
    SRMux I__2171 (
            .O(N__9768),
            .I(N__9642));
    SRMux I__2170 (
            .O(N__9767),
            .I(N__9642));
    SRMux I__2169 (
            .O(N__9766),
            .I(N__9642));
    SRMux I__2168 (
            .O(N__9765),
            .I(N__9642));
    SRMux I__2167 (
            .O(N__9764),
            .I(N__9642));
    SRMux I__2166 (
            .O(N__9763),
            .I(N__9642));
    SRMux I__2165 (
            .O(N__9762),
            .I(N__9642));
    SRMux I__2164 (
            .O(N__9761),
            .I(N__9642));
    SRMux I__2163 (
            .O(N__9760),
            .I(N__9642));
    SRMux I__2162 (
            .O(N__9759),
            .I(N__9642));
    SRMux I__2161 (
            .O(N__9758),
            .I(N__9642));
    SRMux I__2160 (
            .O(N__9757),
            .I(N__9642));
    SRMux I__2159 (
            .O(N__9756),
            .I(N__9642));
    SRMux I__2158 (
            .O(N__9755),
            .I(N__9642));
    SRMux I__2157 (
            .O(N__9754),
            .I(N__9642));
    SRMux I__2156 (
            .O(N__9753),
            .I(N__9642));
    SRMux I__2155 (
            .O(N__9752),
            .I(N__9642));
    SRMux I__2154 (
            .O(N__9751),
            .I(N__9642));
    SRMux I__2153 (
            .O(N__9750),
            .I(N__9642));
    SRMux I__2152 (
            .O(N__9749),
            .I(N__9642));
    Glb2LocalMux I__2151 (
            .O(N__9746),
            .I(N__9642));
    SRMux I__2150 (
            .O(N__9745),
            .I(N__9642));
    SRMux I__2149 (
            .O(N__9744),
            .I(N__9642));
    SRMux I__2148 (
            .O(N__9743),
            .I(N__9642));
    GlobalMux I__2147 (
            .O(N__9642),
            .I(N__9639));
    gio2CtrlBuf I__2146 (
            .O(N__9639),
            .I(RESETn_c_i_g));
    InMux I__2145 (
            .O(N__9636),
            .I(N__9633));
    LocalMux I__2144 (
            .O(N__9633),
            .I(\U712_REG_SM.N_404 ));
    IoInMux I__2143 (
            .O(N__9630),
            .I(N__9627));
    LocalMux I__2142 (
            .O(N__9627),
            .I(N__9624));
    Span4Mux_s0_v I__2141 (
            .O(N__9624),
            .I(N__9621));
    Span4Mux_v I__2140 (
            .O(N__9621),
            .I(N__9618));
    Odrv4 I__2139 (
            .O(N__9618),
            .I(N_335_i));
    IoInMux I__2138 (
            .O(N__9615),
            .I(N__9612));
    LocalMux I__2137 (
            .O(N__9612),
            .I(N__9609));
    Span4Mux_s3_v I__2136 (
            .O(N__9609),
            .I(N__9606));
    Odrv4 I__2135 (
            .O(N__9606),
            .I(N_337_i));
    InMux I__2134 (
            .O(N__9603),
            .I(N__9598));
    InMux I__2133 (
            .O(N__9602),
            .I(N__9593));
    InMux I__2132 (
            .O(N__9601),
            .I(N__9593));
    LocalMux I__2131 (
            .O(N__9598),
            .I(N__9590));
    LocalMux I__2130 (
            .O(N__9593),
            .I(N__9586));
    Span4Mux_v I__2129 (
            .O(N__9590),
            .I(N__9583));
    InMux I__2128 (
            .O(N__9589),
            .I(N__9580));
    Span4Mux_h I__2127 (
            .O(N__9586),
            .I(N__9577));
    Sp12to4 I__2126 (
            .O(N__9583),
            .I(N__9574));
    LocalMux I__2125 (
            .O(N__9580),
            .I(N__9569));
    Sp12to4 I__2124 (
            .O(N__9577),
            .I(N__9569));
    Span12Mux_h I__2123 (
            .O(N__9574),
            .I(N__9566));
    Span12Mux_v I__2122 (
            .O(N__9569),
            .I(N__9563));
    Span12Mux_v I__2121 (
            .O(N__9566),
            .I(N__9560));
    Span12Mux_h I__2120 (
            .O(N__9563),
            .I(N__9557));
    Odrv12 I__2119 (
            .O(N__9560),
            .I(DRA_c_3));
    Odrv12 I__2118 (
            .O(N__9557),
            .I(DRA_c_3));
    InMux I__2117 (
            .O(N__9552),
            .I(N__9548));
    InMux I__2116 (
            .O(N__9551),
            .I(N__9545));
    LocalMux I__2115 (
            .O(N__9548),
            .I(N__9538));
    LocalMux I__2114 (
            .O(N__9545),
            .I(N__9538));
    InMux I__2113 (
            .O(N__9544),
            .I(N__9535));
    InMux I__2112 (
            .O(N__9543),
            .I(N__9532));
    Span4Mux_v I__2111 (
            .O(N__9538),
            .I(N__9529));
    LocalMux I__2110 (
            .O(N__9535),
            .I(N__9526));
    LocalMux I__2109 (
            .O(N__9532),
            .I(N__9521));
    Sp12to4 I__2108 (
            .O(N__9529),
            .I(N__9521));
    Span12Mux_h I__2107 (
            .O(N__9526),
            .I(N__9518));
    Span12Mux_h I__2106 (
            .O(N__9521),
            .I(N__9515));
    Span12Mux_v I__2105 (
            .O(N__9518),
            .I(N__9512));
    Span12Mux_v I__2104 (
            .O(N__9515),
            .I(N__9509));
    Odrv12 I__2103 (
            .O(N__9512),
            .I(DRA_c_2));
    Odrv12 I__2102 (
            .O(N__9509),
            .I(DRA_c_2));
    InMux I__2101 (
            .O(N__9504),
            .I(N__9501));
    LocalMux I__2100 (
            .O(N__9501),
            .I(N__9498));
    Odrv4 I__2099 (
            .O(N__9498),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2098 (
            .O(N__9495),
            .I(N__9490));
    InMux I__2097 (
            .O(N__9494),
            .I(N__9487));
    InMux I__2096 (
            .O(N__9493),
            .I(N__9484));
    LocalMux I__2095 (
            .O(N__9490),
            .I(N__9480));
    LocalMux I__2094 (
            .O(N__9487),
            .I(N__9475));
    LocalMux I__2093 (
            .O(N__9484),
            .I(N__9475));
    InMux I__2092 (
            .O(N__9483),
            .I(N__9472));
    Span4Mux_v I__2091 (
            .O(N__9480),
            .I(N__9469));
    Sp12to4 I__2090 (
            .O(N__9475),
            .I(N__9464));
    LocalMux I__2089 (
            .O(N__9472),
            .I(N__9464));
    Sp12to4 I__2088 (
            .O(N__9469),
            .I(N__9461));
    Span12Mux_v I__2087 (
            .O(N__9464),
            .I(N__9458));
    Span12Mux_h I__2086 (
            .O(N__9461),
            .I(N__9455));
    Span12Mux_h I__2085 (
            .O(N__9458),
            .I(N__9452));
    Odrv12 I__2084 (
            .O(N__9455),
            .I(DRA_c_8));
    Odrv12 I__2083 (
            .O(N__9452),
            .I(DRA_c_8));
    InMux I__2082 (
            .O(N__9447),
            .I(N__9444));
    LocalMux I__2081 (
            .O(N__9444),
            .I(N__9441));
    Span4Mux_h I__2080 (
            .O(N__9441),
            .I(N__9438));
    Odrv4 I__2079 (
            .O(N__9438),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    IoInMux I__2078 (
            .O(N__9435),
            .I(N__9432));
    LocalMux I__2077 (
            .O(N__9432),
            .I(N__9429));
    IoSpan4Mux I__2076 (
            .O(N__9429),
            .I(N__9426));
    Sp12to4 I__2075 (
            .O(N__9426),
            .I(N__9423));
    Span12Mux_v I__2074 (
            .O(N__9423),
            .I(N__9420));
    Span12Mux_h I__2073 (
            .O(N__9420),
            .I(N__9417));
    Odrv12 I__2072 (
            .O(N__9417),
            .I(ASn_c));
    CEMux I__2071 (
            .O(N__9414),
            .I(N__9411));
    LocalMux I__2070 (
            .O(N__9411),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ));
    IoInMux I__2069 (
            .O(N__9408),
            .I(N__9405));
    LocalMux I__2068 (
            .O(N__9405),
            .I(N__9402));
    Span4Mux_s3_v I__2067 (
            .O(N__9402),
            .I(N__9399));
    Odrv4 I__2066 (
            .O(N__9399),
            .I(N_336_i));
    InMux I__2065 (
            .O(N__9396),
            .I(N__9393));
    LocalMux I__2064 (
            .O(N__9393),
            .I(N__9389));
    InMux I__2063 (
            .O(N__9392),
            .I(N__9386));
    Span4Mux_v I__2062 (
            .O(N__9389),
            .I(N__9383));
    LocalMux I__2061 (
            .O(N__9386),
            .I(N__9380));
    Span4Mux_v I__2060 (
            .O(N__9383),
            .I(N__9377));
    Span4Mux_v I__2059 (
            .O(N__9380),
            .I(N__9374));
    Sp12to4 I__2058 (
            .O(N__9377),
            .I(N__9371));
    Sp12to4 I__2057 (
            .O(N__9374),
            .I(N__9368));
    Span12Mux_h I__2056 (
            .O(N__9371),
            .I(N__9365));
    Span12Mux_v I__2055 (
            .O(N__9368),
            .I(N__9362));
    Span12Mux_v I__2054 (
            .O(N__9365),
            .I(N__9359));
    Span12Mux_h I__2053 (
            .O(N__9362),
            .I(N__9356));
    Odrv12 I__2052 (
            .O(N__9359),
            .I(DRA_c_0));
    Odrv12 I__2051 (
            .O(N__9356),
            .I(DRA_c_0));
    InMux I__2050 (
            .O(N__9351),
            .I(N__9346));
    InMux I__2049 (
            .O(N__9350),
            .I(N__9343));
    InMux I__2048 (
            .O(N__9349),
            .I(N__9340));
    LocalMux I__2047 (
            .O(N__9346),
            .I(N__9336));
    LocalMux I__2046 (
            .O(N__9343),
            .I(N__9331));
    LocalMux I__2045 (
            .O(N__9340),
            .I(N__9331));
    InMux I__2044 (
            .O(N__9339),
            .I(N__9328));
    Span4Mux_v I__2043 (
            .O(N__9336),
            .I(N__9325));
    Span4Mux_h I__2042 (
            .O(N__9331),
            .I(N__9320));
    LocalMux I__2041 (
            .O(N__9328),
            .I(N__9320));
    Span4Mux_h I__2040 (
            .O(N__9325),
            .I(N__9317));
    Span4Mux_h I__2039 (
            .O(N__9320),
            .I(N__9314));
    Sp12to4 I__2038 (
            .O(N__9317),
            .I(N__9311));
    Span4Mux_v I__2037 (
            .O(N__9314),
            .I(N__9308));
    Span12Mux_s10_h I__2036 (
            .O(N__9311),
            .I(N__9303));
    Sp12to4 I__2035 (
            .O(N__9308),
            .I(N__9303));
    Span12Mux_v I__2034 (
            .O(N__9303),
            .I(N__9300));
    Odrv12 I__2033 (
            .O(N__9300),
            .I(DRA_c_1));
    InMux I__2032 (
            .O(N__9297),
            .I(N__9294));
    LocalMux I__2031 (
            .O(N__9294),
            .I(N__9291));
    Odrv12 I__2030 (
            .O(N__9291),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2029 (
            .O(N__9288),
            .I(N__9283));
    InMux I__2028 (
            .O(N__9287),
            .I(N__9279));
    InMux I__2027 (
            .O(N__9286),
            .I(N__9276));
    LocalMux I__2026 (
            .O(N__9283),
            .I(N__9273));
    InMux I__2025 (
            .O(N__9282),
            .I(N__9270));
    LocalMux I__2024 (
            .O(N__9279),
            .I(N__9265));
    LocalMux I__2023 (
            .O(N__9276),
            .I(N__9265));
    Span4Mux_v I__2022 (
            .O(N__9273),
            .I(N__9262));
    LocalMux I__2021 (
            .O(N__9270),
            .I(N__9259));
    Span4Mux_v I__2020 (
            .O(N__9265),
            .I(N__9256));
    Span4Mux_v I__2019 (
            .O(N__9262),
            .I(N__9251));
    Span4Mux_v I__2018 (
            .O(N__9259),
            .I(N__9251));
    Span4Mux_v I__2017 (
            .O(N__9256),
            .I(N__9248));
    Sp12to4 I__2016 (
            .O(N__9251),
            .I(N__9243));
    Sp12to4 I__2015 (
            .O(N__9248),
            .I(N__9243));
    Span12Mux_h I__2014 (
            .O(N__9243),
            .I(N__9240));
    Span12Mux_v I__2013 (
            .O(N__9240),
            .I(N__9237));
    Odrv12 I__2012 (
            .O(N__9237),
            .I(DRA_c_9));
    InMux I__2011 (
            .O(N__9234),
            .I(N__9231));
    LocalMux I__2010 (
            .O(N__9231),
            .I(N__9228));
    Span4Mux_h I__2009 (
            .O(N__9228),
            .I(N__9225));
    Odrv4 I__2008 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2007 (
            .O(N__9222),
            .I(N__9201));
    ClkMux I__2006 (
            .O(N__9221),
            .I(N__9201));
    ClkMux I__2005 (
            .O(N__9220),
            .I(N__9201));
    ClkMux I__2004 (
            .O(N__9219),
            .I(N__9201));
    ClkMux I__2003 (
            .O(N__9218),
            .I(N__9201));
    ClkMux I__2002 (
            .O(N__9217),
            .I(N__9201));
    ClkMux I__2001 (
            .O(N__9216),
            .I(N__9201));
    GlobalMux I__2000 (
            .O(N__9201),
            .I(N__9198));
    gio2CtrlBuf I__1999 (
            .O(N__9198),
            .I(C3_c_g));
    IoInMux I__1998 (
            .O(N__9195),
            .I(N__9192));
    LocalMux I__1997 (
            .O(N__9192),
            .I(N__9189));
    Span12Mux_s6_v I__1996 (
            .O(N__9189),
            .I(N__9186));
    Odrv12 I__1995 (
            .O(N__9186),
            .I(RESETn_c_i));
    CascadeMux I__1994 (
            .O(N__9183),
            .I(N__9180));
    InMux I__1993 (
            .O(N__9180),
            .I(N__9177));
    LocalMux I__1992 (
            .O(N__9177),
            .I(N__9174));
    Odrv12 I__1991 (
            .O(N__9174),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1990 (
            .O(N__9171),
            .I(N__9167));
    InMux I__1989 (
            .O(N__9170),
            .I(N__9164));
    LocalMux I__1988 (
            .O(N__9167),
            .I(N__9158));
    LocalMux I__1987 (
            .O(N__9164),
            .I(N__9158));
    InMux I__1986 (
            .O(N__9163),
            .I(N__9155));
    Span4Mux_v I__1985 (
            .O(N__9158),
            .I(N__9151));
    LocalMux I__1984 (
            .O(N__9155),
            .I(N__9148));
    InMux I__1983 (
            .O(N__9154),
            .I(N__9145));
    Sp12to4 I__1982 (
            .O(N__9151),
            .I(N__9142));
    Sp12to4 I__1981 (
            .O(N__9148),
            .I(N__9137));
    LocalMux I__1980 (
            .O(N__9145),
            .I(N__9137));
    Span12Mux_h I__1979 (
            .O(N__9142),
            .I(N__9134));
    Span12Mux_v I__1978 (
            .O(N__9137),
            .I(N__9131));
    Span12Mux_v I__1977 (
            .O(N__9134),
            .I(N__9126));
    Span12Mux_h I__1976 (
            .O(N__9131),
            .I(N__9126));
    Odrv12 I__1975 (
            .O(N__9126),
            .I(DRA_c_4));
    InMux I__1974 (
            .O(N__9123),
            .I(N__9120));
    LocalMux I__1973 (
            .O(N__9120),
            .I(N__9117));
    Span4Mux_h I__1972 (
            .O(N__9117),
            .I(N__9114));
    Odrv4 I__1971 (
            .O(N__9114),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1970 (
            .O(N__9111),
            .I(N__9108));
    LocalMux I__1969 (
            .O(N__9108),
            .I(N__9105));
    Span4Mux_h I__1968 (
            .O(N__9105),
            .I(N__9102));
    Odrv4 I__1967 (
            .O(N__9102),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1966 (
            .O(N__9099),
            .I(N__9096));
    LocalMux I__1965 (
            .O(N__9096),
            .I(N__9093));
    Odrv12 I__1964 (
            .O(N__9093),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1963 (
            .O(N__9090),
            .I(N__9087));
    LocalMux I__1962 (
            .O(N__9087),
            .I(N__9084));
    Odrv12 I__1961 (
            .O(N__9084),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1960 (
            .O(N__9081),
            .I(N__9078));
    LocalMux I__1959 (
            .O(N__9078),
            .I(N__9075));
    Span4Mux_v I__1958 (
            .O(N__9075),
            .I(N__9072));
    Odrv4 I__1957 (
            .O(N__9072),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1956 (
            .O(N__9069),
            .I(N__9063));
    InMux I__1955 (
            .O(N__9068),
            .I(N__9060));
    InMux I__1954 (
            .O(N__9067),
            .I(N__9057));
    InMux I__1953 (
            .O(N__9066),
            .I(N__9054));
    LocalMux I__1952 (
            .O(N__9063),
            .I(N__9049));
    LocalMux I__1951 (
            .O(N__9060),
            .I(N__9049));
    LocalMux I__1950 (
            .O(N__9057),
            .I(N__9044));
    LocalMux I__1949 (
            .O(N__9054),
            .I(N__9044));
    Span4Mux_v I__1948 (
            .O(N__9049),
            .I(N__9039));
    Span4Mux_v I__1947 (
            .O(N__9044),
            .I(N__9039));
    Sp12to4 I__1946 (
            .O(N__9039),
            .I(N__9036));
    Span12Mux_h I__1945 (
            .O(N__9036),
            .I(N__9033));
    Odrv12 I__1944 (
            .O(N__9033),
            .I(DRA_c_7));
    InMux I__1943 (
            .O(N__9030),
            .I(N__9027));
    LocalMux I__1942 (
            .O(N__9027),
            .I(N__9024));
    Odrv4 I__1941 (
            .O(N__9024),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1940 (
            .O(N__9021),
            .I(N__9018));
    LocalMux I__1939 (
            .O(N__9018),
            .I(N__9015));
    Odrv12 I__1938 (
            .O(N__9015),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__1937 (
            .O(N__9012),
            .I(N__9009));
    LocalMux I__1936 (
            .O(N__9009),
            .I(\U712_REG_SM.N_373 ));
    CascadeMux I__1935 (
            .O(N__9006),
            .I(\U712_REG_SM.N_330_cascade_ ));
    InMux I__1934 (
            .O(N__9003),
            .I(N__9000));
    LocalMux I__1933 (
            .O(N__9000),
            .I(\U712_REG_SM.N_413 ));
    InMux I__1932 (
            .O(N__8997),
            .I(N__8990));
    InMux I__1931 (
            .O(N__8996),
            .I(N__8987));
    InMux I__1930 (
            .O(N__8995),
            .I(N__8984));
    InMux I__1929 (
            .O(N__8994),
            .I(N__8979));
    InMux I__1928 (
            .O(N__8993),
            .I(N__8979));
    LocalMux I__1927 (
            .O(N__8990),
            .I(N__8976));
    LocalMux I__1926 (
            .O(N__8987),
            .I(N__8973));
    LocalMux I__1925 (
            .O(N__8984),
            .I(N__8968));
    LocalMux I__1924 (
            .O(N__8979),
            .I(N__8968));
    Odrv4 I__1923 (
            .O(N__8976),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1922 (
            .O(N__8973),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1921 (
            .O(N__8968),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1920 (
            .O(N__8961),
            .I(N__8958));
    LocalMux I__1919 (
            .O(N__8958),
            .I(\U712_REG_SM.N_410 ));
    CascadeMux I__1918 (
            .O(N__8955),
            .I(N__8950));
    InMux I__1917 (
            .O(N__8954),
            .I(N__8942));
    InMux I__1916 (
            .O(N__8953),
            .I(N__8942));
    InMux I__1915 (
            .O(N__8950),
            .I(N__8942));
    InMux I__1914 (
            .O(N__8949),
            .I(N__8939));
    LocalMux I__1913 (
            .O(N__8942),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1912 (
            .O(N__8939),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__1911 (
            .O(N__8934),
            .I(N__8931));
    LocalMux I__1910 (
            .O(N__8931),
            .I(\U712_REG_SM.STATE_COUNTc_0_0 ));
    InMux I__1909 (
            .O(N__8928),
            .I(N__8925));
    LocalMux I__1908 (
            .O(N__8925),
            .I(\U712_REG_SM.N_308 ));
    InMux I__1907 (
            .O(N__8922),
            .I(N__8918));
    InMux I__1906 (
            .O(N__8921),
            .I(N__8915));
    LocalMux I__1905 (
            .O(N__8918),
            .I(N__8906));
    LocalMux I__1904 (
            .O(N__8915),
            .I(N__8906));
    InMux I__1903 (
            .O(N__8914),
            .I(N__8903));
    InMux I__1902 (
            .O(N__8913),
            .I(N__8898));
    InMux I__1901 (
            .O(N__8912),
            .I(N__8898));
    InMux I__1900 (
            .O(N__8911),
            .I(N__8895));
    Odrv4 I__1899 (
            .O(N__8906),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1898 (
            .O(N__8903),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1897 (
            .O(N__8898),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1896 (
            .O(N__8895),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__1895 (
            .O(N__8886),
            .I(\U712_REG_SM.N_308_cascade_ ));
    InMux I__1894 (
            .O(N__8883),
            .I(N__8878));
    InMux I__1893 (
            .O(N__8882),
            .I(N__8873));
    InMux I__1892 (
            .O(N__8881),
            .I(N__8870));
    LocalMux I__1891 (
            .O(N__8878),
            .I(N__8867));
    InMux I__1890 (
            .O(N__8877),
            .I(N__8862));
    InMux I__1889 (
            .O(N__8876),
            .I(N__8862));
    LocalMux I__1888 (
            .O(N__8873),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1887 (
            .O(N__8870),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__1886 (
            .O(N__8867),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1885 (
            .O(N__8862),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1884 (
            .O(N__8853),
            .I(N__8849));
    CascadeMux I__1883 (
            .O(N__8852),
            .I(N__8838));
    InMux I__1882 (
            .O(N__8849),
            .I(N__8833));
    InMux I__1881 (
            .O(N__8848),
            .I(N__8830));
    InMux I__1880 (
            .O(N__8847),
            .I(N__8825));
    InMux I__1879 (
            .O(N__8846),
            .I(N__8825));
    InMux I__1878 (
            .O(N__8845),
            .I(N__8822));
    InMux I__1877 (
            .O(N__8844),
            .I(N__8819));
    InMux I__1876 (
            .O(N__8843),
            .I(N__8810));
    InMux I__1875 (
            .O(N__8842),
            .I(N__8810));
    InMux I__1874 (
            .O(N__8841),
            .I(N__8810));
    InMux I__1873 (
            .O(N__8838),
            .I(N__8810));
    InMux I__1872 (
            .O(N__8837),
            .I(N__8805));
    InMux I__1871 (
            .O(N__8836),
            .I(N__8805));
    LocalMux I__1870 (
            .O(N__8833),
            .I(N__8796));
    LocalMux I__1869 (
            .O(N__8830),
            .I(N__8796));
    LocalMux I__1868 (
            .O(N__8825),
            .I(N__8796));
    LocalMux I__1867 (
            .O(N__8822),
            .I(N__8796));
    LocalMux I__1866 (
            .O(N__8819),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1865 (
            .O(N__8810),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1864 (
            .O(N__8805),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1863 (
            .O(N__8796),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__1862 (
            .O(N__8787),
            .I(N__8782));
    CascadeMux I__1861 (
            .O(N__8786),
            .I(N__8779));
    InMux I__1860 (
            .O(N__8785),
            .I(N__8773));
    InMux I__1859 (
            .O(N__8782),
            .I(N__8770));
    InMux I__1858 (
            .O(N__8779),
            .I(N__8767));
    InMux I__1857 (
            .O(N__8778),
            .I(N__8762));
    InMux I__1856 (
            .O(N__8777),
            .I(N__8762));
    InMux I__1855 (
            .O(N__8776),
            .I(N__8759));
    LocalMux I__1854 (
            .O(N__8773),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1853 (
            .O(N__8770),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1852 (
            .O(N__8767),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1851 (
            .O(N__8762),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1850 (
            .O(N__8759),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    InMux I__1849 (
            .O(N__8748),
            .I(N__8745));
    LocalMux I__1848 (
            .O(N__8745),
            .I(N__8742));
    Span4Mux_h I__1847 (
            .O(N__8742),
            .I(N__8739));
    Odrv4 I__1846 (
            .O(N__8739),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1845 (
            .O(N__8736),
            .I(N__8733));
    LocalMux I__1844 (
            .O(N__8733),
            .I(N__8730));
    Odrv4 I__1843 (
            .O(N__8730),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1842 (
            .O(N__8727),
            .I(N__8724));
    LocalMux I__1841 (
            .O(N__8724),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1840 (
            .O(N__8721),
            .I(N__8718));
    LocalMux I__1839 (
            .O(N__8718),
            .I(\U712_CYCLE_TERM.N_332 ));
    InMux I__1838 (
            .O(N__8715),
            .I(N__8705));
    InMux I__1837 (
            .O(N__8714),
            .I(N__8705));
    InMux I__1836 (
            .O(N__8713),
            .I(N__8705));
    CascadeMux I__1835 (
            .O(N__8712),
            .I(N__8702));
    LocalMux I__1834 (
            .O(N__8705),
            .I(N__8699));
    InMux I__1833 (
            .O(N__8702),
            .I(N__8696));
    Span4Mux_h I__1832 (
            .O(N__8699),
            .I(N__8693));
    LocalMux I__1831 (
            .O(N__8696),
            .I(CPU_TACKm));
    Odrv4 I__1830 (
            .O(N__8693),
            .I(CPU_TACKm));
    InMux I__1829 (
            .O(N__8688),
            .I(N__8682));
    InMux I__1828 (
            .O(N__8687),
            .I(N__8675));
    InMux I__1827 (
            .O(N__8686),
            .I(N__8675));
    InMux I__1826 (
            .O(N__8685),
            .I(N__8675));
    LocalMux I__1825 (
            .O(N__8682),
            .I(REG_TACK));
    LocalMux I__1824 (
            .O(N__8675),
            .I(REG_TACK));
    CascadeMux I__1823 (
            .O(N__8670),
            .I(N__8667));
    InMux I__1822 (
            .O(N__8667),
            .I(N__8662));
    InMux I__1821 (
            .O(N__8666),
            .I(N__8657));
    InMux I__1820 (
            .O(N__8665),
            .I(N__8657));
    LocalMux I__1819 (
            .O(N__8662),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1818 (
            .O(N__8657),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__1817 (
            .O(N__8652),
            .I(\U712_CYCLE_TERM.N_455_cascade_ ));
    InMux I__1816 (
            .O(N__8649),
            .I(N__8645));
    InMux I__1815 (
            .O(N__8648),
            .I(N__8642));
    LocalMux I__1814 (
            .O(N__8645),
            .I(N__8637));
    LocalMux I__1813 (
            .O(N__8642),
            .I(N__8634));
    InMux I__1812 (
            .O(N__8641),
            .I(N__8631));
    InMux I__1811 (
            .O(N__8640),
            .I(N__8628));
    Odrv4 I__1810 (
            .O(N__8637),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__1809 (
            .O(N__8634),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1808 (
            .O(N__8631),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1807 (
            .O(N__8628),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1806 (
            .O(N__8619),
            .I(N__8616));
    LocalMux I__1805 (
            .O(N__8616),
            .I(N__8612));
    InMux I__1804 (
            .O(N__8615),
            .I(N__8609));
    Span4Mux_v I__1803 (
            .O(N__8612),
            .I(N__8606));
    LocalMux I__1802 (
            .O(N__8609),
            .I(N__8603));
    Span4Mux_h I__1801 (
            .O(N__8606),
            .I(N__8598));
    Span4Mux_h I__1800 (
            .O(N__8603),
            .I(N__8598));
    Odrv4 I__1799 (
            .O(N__8598),
            .I(DBRn_c_i));
    InMux I__1798 (
            .O(N__8595),
            .I(N__8591));
    CascadeMux I__1797 (
            .O(N__8594),
            .I(N__8588));
    LocalMux I__1796 (
            .O(N__8591),
            .I(N__8585));
    InMux I__1795 (
            .O(N__8588),
            .I(N__8582));
    Span4Mux_h I__1794 (
            .O(N__8585),
            .I(N__8579));
    LocalMux I__1793 (
            .O(N__8582),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__1792 (
            .O(N__8579),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1791 (
            .O(N__8574),
            .I(N__8570));
    InMux I__1790 (
            .O(N__8573),
            .I(N__8565));
    LocalMux I__1789 (
            .O(N__8570),
            .I(N__8562));
    InMux I__1788 (
            .O(N__8569),
            .I(N__8559));
    InMux I__1787 (
            .O(N__8568),
            .I(N__8556));
    LocalMux I__1786 (
            .O(N__8565),
            .I(N__8553));
    Span4Mux_v I__1785 (
            .O(N__8562),
            .I(N__8550));
    LocalMux I__1784 (
            .O(N__8559),
            .I(N__8543));
    LocalMux I__1783 (
            .O(N__8556),
            .I(N__8543));
    Span4Mux_h I__1782 (
            .O(N__8553),
            .I(N__8543));
    Span4Mux_v I__1781 (
            .O(N__8550),
            .I(N__8540));
    Span4Mux_v I__1780 (
            .O(N__8543),
            .I(N__8537));
    Span4Mux_v I__1779 (
            .O(N__8540),
            .I(N__8534));
    Span4Mux_v I__1778 (
            .O(N__8537),
            .I(N__8531));
    IoSpan4Mux I__1777 (
            .O(N__8534),
            .I(N__8528));
    Span4Mux_v I__1776 (
            .O(N__8531),
            .I(N__8525));
    Odrv4 I__1775 (
            .O(N__8528),
            .I(CLK40_PLL_i));
    Odrv4 I__1774 (
            .O(N__8525),
            .I(CLK40_PLL_i));
    IoInMux I__1773 (
            .O(N__8520),
            .I(N__8517));
    LocalMux I__1772 (
            .O(N__8517),
            .I(N__8514));
    IoSpan4Mux I__1771 (
            .O(N__8514),
            .I(N__8510));
    IoInMux I__1770 (
            .O(N__8513),
            .I(N__8507));
    Span4Mux_s3_h I__1769 (
            .O(N__8510),
            .I(N__8502));
    LocalMux I__1768 (
            .O(N__8507),
            .I(N__8502));
    Span4Mux_s2_v I__1767 (
            .O(N__8502),
            .I(N__8499));
    Span4Mux_v I__1766 (
            .O(N__8499),
            .I(N__8495));
    IoInMux I__1765 (
            .O(N__8498),
            .I(N__8492));
    Sp12to4 I__1764 (
            .O(N__8495),
            .I(N__8489));
    LocalMux I__1763 (
            .O(N__8492),
            .I(N__8486));
    Span12Mux_h I__1762 (
            .O(N__8489),
            .I(N__8483));
    Span12Mux_s9_h I__1761 (
            .O(N__8486),
            .I(N__8480));
    Odrv12 I__1760 (
            .O(N__8483),
            .I(CLK40_PLL_i_i));
    Odrv12 I__1759 (
            .O(N__8480),
            .I(CLK40_PLL_i_i));
    InMux I__1758 (
            .O(N__8475),
            .I(N__8472));
    LocalMux I__1757 (
            .O(N__8472),
            .I(\U712_REG_SM.N_412 ));
    InMux I__1756 (
            .O(N__8469),
            .I(N__8465));
    IoInMux I__1755 (
            .O(N__8468),
            .I(N__8462));
    LocalMux I__1754 (
            .O(N__8465),
            .I(N__8459));
    LocalMux I__1753 (
            .O(N__8462),
            .I(N__8456));
    Sp12to4 I__1752 (
            .O(N__8459),
            .I(N__8453));
    IoSpan4Mux I__1751 (
            .O(N__8456),
            .I(N__8450));
    Span12Mux_v I__1750 (
            .O(N__8453),
            .I(N__8447));
    IoSpan4Mux I__1749 (
            .O(N__8450),
            .I(N__8444));
    Span12Mux_h I__1748 (
            .O(N__8447),
            .I(N__8441));
    IoSpan4Mux I__1747 (
            .O(N__8444),
            .I(N__8438));
    Odrv12 I__1746 (
            .O(N__8441),
            .I(C1_c));
    Odrv4 I__1745 (
            .O(N__8438),
            .I(C1_c));
    InMux I__1744 (
            .O(N__8433),
            .I(N__8430));
    LocalMux I__1743 (
            .O(N__8430),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__1742 (
            .O(N__8427),
            .I(N__8424));
    LocalMux I__1741 (
            .O(N__8424),
            .I(N__8421));
    Odrv4 I__1740 (
            .O(N__8421),
            .I(\U712_REG_SM.REGENn_e_1 ));
    InMux I__1739 (
            .O(N__8418),
            .I(N__8415));
    LocalMux I__1738 (
            .O(N__8415),
            .I(N__8411));
    InMux I__1737 (
            .O(N__8414),
            .I(N__8408));
    Odrv4 I__1736 (
            .O(N__8411),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    LocalMux I__1735 (
            .O(N__8408),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    IoInMux I__1734 (
            .O(N__8403),
            .I(N__8400));
    LocalMux I__1733 (
            .O(N__8400),
            .I(N__8397));
    Span4Mux_s0_v I__1732 (
            .O(N__8397),
            .I(N__8394));
    Sp12to4 I__1731 (
            .O(N__8394),
            .I(N__8390));
    InMux I__1730 (
            .O(N__8393),
            .I(N__8386));
    Span12Mux_h I__1729 (
            .O(N__8390),
            .I(N__8383));
    InMux I__1728 (
            .O(N__8389),
            .I(N__8380));
    LocalMux I__1727 (
            .O(N__8386),
            .I(N__8377));
    Odrv12 I__1726 (
            .O(N__8383),
            .I(REGENn_c));
    LocalMux I__1725 (
            .O(N__8380),
            .I(REGENn_c));
    Odrv4 I__1724 (
            .O(N__8377),
            .I(REGENn_c));
    CascadeMux I__1723 (
            .O(N__8370),
            .I(N__8362));
    CascadeMux I__1722 (
            .O(N__8369),
            .I(N__8359));
    CascadeMux I__1721 (
            .O(N__8368),
            .I(N__8355));
    CascadeMux I__1720 (
            .O(N__8367),
            .I(N__8350));
    InMux I__1719 (
            .O(N__8366),
            .I(N__8347));
    InMux I__1718 (
            .O(N__8365),
            .I(N__8342));
    InMux I__1717 (
            .O(N__8362),
            .I(N__8342));
    InMux I__1716 (
            .O(N__8359),
            .I(N__8339));
    InMux I__1715 (
            .O(N__8358),
            .I(N__8335));
    InMux I__1714 (
            .O(N__8355),
            .I(N__8321));
    InMux I__1713 (
            .O(N__8354),
            .I(N__8321));
    InMux I__1712 (
            .O(N__8353),
            .I(N__8321));
    InMux I__1711 (
            .O(N__8350),
            .I(N__8321));
    LocalMux I__1710 (
            .O(N__8347),
            .I(N__8316));
    LocalMux I__1709 (
            .O(N__8342),
            .I(N__8316));
    LocalMux I__1708 (
            .O(N__8339),
            .I(N__8310));
    CascadeMux I__1707 (
            .O(N__8338),
            .I(N__8307));
    LocalMux I__1706 (
            .O(N__8335),
            .I(N__8301));
    InMux I__1705 (
            .O(N__8334),
            .I(N__8298));
    InMux I__1704 (
            .O(N__8333),
            .I(N__8291));
    InMux I__1703 (
            .O(N__8332),
            .I(N__8291));
    InMux I__1702 (
            .O(N__8331),
            .I(N__8291));
    CascadeMux I__1701 (
            .O(N__8330),
            .I(N__8287));
    LocalMux I__1700 (
            .O(N__8321),
            .I(N__8279));
    Span4Mux_v I__1699 (
            .O(N__8316),
            .I(N__8279));
    InMux I__1698 (
            .O(N__8315),
            .I(N__8272));
    InMux I__1697 (
            .O(N__8314),
            .I(N__8272));
    InMux I__1696 (
            .O(N__8313),
            .I(N__8272));
    Span4Mux_h I__1695 (
            .O(N__8310),
            .I(N__8269));
    InMux I__1694 (
            .O(N__8307),
            .I(N__8260));
    InMux I__1693 (
            .O(N__8306),
            .I(N__8260));
    InMux I__1692 (
            .O(N__8305),
            .I(N__8260));
    InMux I__1691 (
            .O(N__8304),
            .I(N__8260));
    Span4Mux_v I__1690 (
            .O(N__8301),
            .I(N__8257));
    LocalMux I__1689 (
            .O(N__8298),
            .I(N__8252));
    LocalMux I__1688 (
            .O(N__8291),
            .I(N__8252));
    InMux I__1687 (
            .O(N__8290),
            .I(N__8241));
    InMux I__1686 (
            .O(N__8287),
            .I(N__8241));
    InMux I__1685 (
            .O(N__8286),
            .I(N__8241));
    InMux I__1684 (
            .O(N__8285),
            .I(N__8241));
    InMux I__1683 (
            .O(N__8284),
            .I(N__8241));
    Odrv4 I__1682 (
            .O(N__8279),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1681 (
            .O(N__8272),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1680 (
            .O(N__8269),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1679 (
            .O(N__8260),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1678 (
            .O(N__8257),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1677 (
            .O(N__8252),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1676 (
            .O(N__8241),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1675 (
            .O(N__8226),
            .I(N__8223));
    LocalMux I__1674 (
            .O(N__8223),
            .I(N__8220));
    Span12Mux_s8_v I__1673 (
            .O(N__8220),
            .I(N__8217));
    Span12Mux_h I__1672 (
            .O(N__8217),
            .I(N__8214));
    Odrv12 I__1671 (
            .O(N__8214),
            .I(CASn_c));
    InMux I__1670 (
            .O(N__8211),
            .I(N__8208));
    LocalMux I__1669 (
            .O(N__8208),
            .I(N__8205));
    Odrv4 I__1668 (
            .O(N__8205),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1667 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1666 (
            .O(N__8199),
            .I(N__8195));
    InMux I__1665 (
            .O(N__8198),
            .I(N__8192));
    Span4Mux_v I__1664 (
            .O(N__8195),
            .I(N__8187));
    LocalMux I__1663 (
            .O(N__8192),
            .I(N__8187));
    Odrv4 I__1662 (
            .O(N__8187),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1661 (
            .O(N__8184),
            .I(N__8181));
    LocalMux I__1660 (
            .O(N__8181),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1659 (
            .O(N__8178),
            .I(N__8175));
    LocalMux I__1658 (
            .O(N__8175),
            .I(N__8172));
    Odrv4 I__1657 (
            .O(N__8172),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    IoInMux I__1656 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__1655 (
            .O(N__8166),
            .I(N__8163));
    IoSpan4Mux I__1654 (
            .O(N__8163),
            .I(N__8160));
    Span4Mux_s3_h I__1653 (
            .O(N__8160),
            .I(N__8157));
    Span4Mux_h I__1652 (
            .O(N__8157),
            .I(N__8154));
    Sp12to4 I__1651 (
            .O(N__8154),
            .I(N__8150));
    InMux I__1650 (
            .O(N__8153),
            .I(N__8147));
    Span12Mux_h I__1649 (
            .O(N__8150),
            .I(N__8142));
    LocalMux I__1648 (
            .O(N__8147),
            .I(N__8142));
    Span12Mux_h I__1647 (
            .O(N__8142),
            .I(N__8139));
    Span12Mux_v I__1646 (
            .O(N__8139),
            .I(N__8136));
    Odrv12 I__1645 (
            .O(N__8136),
            .I(C3_c));
    InMux I__1644 (
            .O(N__8133),
            .I(N__8129));
    InMux I__1643 (
            .O(N__8132),
            .I(N__8126));
    LocalMux I__1642 (
            .O(N__8129),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__1641 (
            .O(N__8126),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__1640 (
            .O(N__8121),
            .I(N__8118));
    LocalMux I__1639 (
            .O(N__8118),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__1638 (
            .O(N__8115),
            .I(\U712_REG_SM.N_328_cascade_ ));
    CascadeMux I__1637 (
            .O(N__8112),
            .I(\U712_REG_SM.N_331_cascade_ ));
    InMux I__1636 (
            .O(N__8109),
            .I(N__8103));
    InMux I__1635 (
            .O(N__8108),
            .I(N__8100));
    InMux I__1634 (
            .O(N__8107),
            .I(N__8095));
    InMux I__1633 (
            .O(N__8106),
            .I(N__8095));
    LocalMux I__1632 (
            .O(N__8103),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1631 (
            .O(N__8100),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1630 (
            .O(N__8095),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__1629 (
            .O(N__8088),
            .I(N__8083));
    InMux I__1628 (
            .O(N__8087),
            .I(N__8080));
    InMux I__1627 (
            .O(N__8086),
            .I(N__8077));
    LocalMux I__1626 (
            .O(N__8083),
            .I(N__8074));
    LocalMux I__1625 (
            .O(N__8080),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1624 (
            .O(N__8077),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    Odrv4 I__1623 (
            .O(N__8074),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    CascadeMux I__1622 (
            .O(N__8067),
            .I(N__8063));
    InMux I__1621 (
            .O(N__8066),
            .I(N__8060));
    InMux I__1620 (
            .O(N__8063),
            .I(N__8057));
    LocalMux I__1619 (
            .O(N__8060),
            .I(N__8054));
    LocalMux I__1618 (
            .O(N__8057),
            .I(\U712_REG_SM.N_328 ));
    Odrv4 I__1617 (
            .O(N__8054),
            .I(\U712_REG_SM.N_328 ));
    IoInMux I__1616 (
            .O(N__8049),
            .I(N__8046));
    LocalMux I__1615 (
            .O(N__8046),
            .I(N__8042));
    IoInMux I__1614 (
            .O(N__8045),
            .I(N__8039));
    IoSpan4Mux I__1613 (
            .O(N__8042),
            .I(N__8036));
    LocalMux I__1612 (
            .O(N__8039),
            .I(N__8032));
    Span4Mux_s2_v I__1611 (
            .O(N__8036),
            .I(N__8029));
    IoInMux I__1610 (
            .O(N__8035),
            .I(N__8026));
    IoSpan4Mux I__1609 (
            .O(N__8032),
            .I(N__8023));
    Sp12to4 I__1608 (
            .O(N__8029),
            .I(N__8020));
    LocalMux I__1607 (
            .O(N__8026),
            .I(N__8017));
    Span4Mux_s3_v I__1606 (
            .O(N__8023),
            .I(N__8014));
    Span12Mux_h I__1605 (
            .O(N__8020),
            .I(N__8011));
    Span12Mux_s7_h I__1604 (
            .O(N__8017),
            .I(N__8008));
    Sp12to4 I__1603 (
            .O(N__8014),
            .I(N__8005));
    Span12Mux_v I__1602 (
            .O(N__8011),
            .I(N__7997));
    Span12Mux_v I__1601 (
            .O(N__8008),
            .I(N__7997));
    Span12Mux_v I__1600 (
            .O(N__8005),
            .I(N__7997));
    InMux I__1599 (
            .O(N__8004),
            .I(N__7994));
    Odrv12 I__1598 (
            .O(N__7997),
            .I(TACK_EN));
    LocalMux I__1597 (
            .O(N__7994),
            .I(TACK_EN));
    InMux I__1596 (
            .O(N__7989),
            .I(N__7986));
    LocalMux I__1595 (
            .O(N__7986),
            .I(N__7982));
    InMux I__1594 (
            .O(N__7985),
            .I(N__7979));
    Odrv4 I__1593 (
            .O(N__7982),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1592 (
            .O(N__7979),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__1591 (
            .O(N__7974),
            .I(\U712_REG_SM.N_373_cascade_ ));
    InMux I__1590 (
            .O(N__7971),
            .I(N__7968));
    LocalMux I__1589 (
            .O(N__7968),
            .I(\U712_REG_SM.N_130 ));
    CascadeMux I__1588 (
            .O(N__7965),
            .I(N__7962));
    InMux I__1587 (
            .O(N__7962),
            .I(N__7958));
    CascadeMux I__1586 (
            .O(N__7961),
            .I(N__7955));
    LocalMux I__1585 (
            .O(N__7958),
            .I(N__7951));
    InMux I__1584 (
            .O(N__7955),
            .I(N__7946));
    InMux I__1583 (
            .O(N__7954),
            .I(N__7946));
    Odrv4 I__1582 (
            .O(N__7951),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1581 (
            .O(N__7946),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1580 (
            .O(N__7941),
            .I(N__7935));
    InMux I__1579 (
            .O(N__7940),
            .I(N__7935));
    LocalMux I__1578 (
            .O(N__7935),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    CascadeMux I__1577 (
            .O(N__7932),
            .I(N__7929));
    InMux I__1576 (
            .O(N__7929),
            .I(N__7926));
    LocalMux I__1575 (
            .O(N__7926),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__1574 (
            .O(N__7923),
            .I(N__7920));
    InMux I__1573 (
            .O(N__7920),
            .I(N__7917));
    LocalMux I__1572 (
            .O(N__7917),
            .I(\U712_REG_SM.N_406 ));
    InMux I__1571 (
            .O(N__7914),
            .I(N__7910));
    InMux I__1570 (
            .O(N__7913),
            .I(N__7907));
    LocalMux I__1569 (
            .O(N__7910),
            .I(N__7899));
    LocalMux I__1568 (
            .O(N__7907),
            .I(N__7899));
    InMux I__1567 (
            .O(N__7906),
            .I(N__7896));
    InMux I__1566 (
            .O(N__7905),
            .I(N__7893));
    InMux I__1565 (
            .O(N__7904),
            .I(N__7890));
    Span4Mux_v I__1564 (
            .O(N__7899),
            .I(N__7883));
    LocalMux I__1563 (
            .O(N__7896),
            .I(N__7883));
    LocalMux I__1562 (
            .O(N__7893),
            .I(N__7883));
    LocalMux I__1561 (
            .O(N__7890),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1560 (
            .O(N__7883),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1559 (
            .O(N__7878),
            .I(N__7875));
    LocalMux I__1558 (
            .O(N__7875),
            .I(N__7872));
    Span4Mux_s3_v I__1557 (
            .O(N__7872),
            .I(N__7869));
    Span4Mux_v I__1556 (
            .O(N__7869),
            .I(N__7866));
    Span4Mux_h I__1555 (
            .O(N__7866),
            .I(N__7863));
    Span4Mux_h I__1554 (
            .O(N__7863),
            .I(N__7860));
    Odrv4 I__1553 (
            .O(N__7860),
            .I(CMA_c_10));
    InMux I__1552 (
            .O(N__7857),
            .I(N__7854));
    LocalMux I__1551 (
            .O(N__7854),
            .I(N__7851));
    Span4Mux_h I__1550 (
            .O(N__7851),
            .I(N__7848));
    Odrv4 I__1549 (
            .O(N__7848),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    CascadeMux I__1548 (
            .O(N__7845),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ));
    IoInMux I__1547 (
            .O(N__7842),
            .I(N__7839));
    LocalMux I__1546 (
            .O(N__7839),
            .I(N__7836));
    Span12Mux_s5_v I__1545 (
            .O(N__7836),
            .I(N__7833));
    Odrv12 I__1544 (
            .O(N__7833),
            .I(CMA_c_2));
    InMux I__1543 (
            .O(N__7830),
            .I(N__7827));
    LocalMux I__1542 (
            .O(N__7827),
            .I(N__7824));
    Odrv4 I__1541 (
            .O(N__7824),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    IoInMux I__1540 (
            .O(N__7821),
            .I(N__7818));
    LocalMux I__1539 (
            .O(N__7818),
            .I(N__7815));
    IoSpan4Mux I__1538 (
            .O(N__7815),
            .I(N__7812));
    Span4Mux_s3_h I__1537 (
            .O(N__7812),
            .I(N__7809));
    Sp12to4 I__1536 (
            .O(N__7809),
            .I(N__7806));
    Span12Mux_h I__1535 (
            .O(N__7806),
            .I(N__7803));
    Odrv12 I__1534 (
            .O(N__7803),
            .I(CMA_c_4));
    InMux I__1533 (
            .O(N__7800),
            .I(N__7793));
    InMux I__1532 (
            .O(N__7799),
            .I(N__7793));
    InMux I__1531 (
            .O(N__7798),
            .I(N__7790));
    LocalMux I__1530 (
            .O(N__7793),
            .I(N__7783));
    LocalMux I__1529 (
            .O(N__7790),
            .I(N__7780));
    InMux I__1528 (
            .O(N__7789),
            .I(N__7777));
    InMux I__1527 (
            .O(N__7788),
            .I(N__7772));
    InMux I__1526 (
            .O(N__7787),
            .I(N__7772));
    InMux I__1525 (
            .O(N__7786),
            .I(N__7769));
    Odrv4 I__1524 (
            .O(N__7783),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    Odrv12 I__1523 (
            .O(N__7780),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1522 (
            .O(N__7777),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1521 (
            .O(N__7772),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1520 (
            .O(N__7769),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    CascadeMux I__1519 (
            .O(N__7758),
            .I(N__7750));
    CascadeMux I__1518 (
            .O(N__7757),
            .I(N__7747));
    CascadeMux I__1517 (
            .O(N__7756),
            .I(N__7744));
    CascadeMux I__1516 (
            .O(N__7755),
            .I(N__7741));
    CascadeMux I__1515 (
            .O(N__7754),
            .I(N__7737));
    CascadeMux I__1514 (
            .O(N__7753),
            .I(N__7733));
    InMux I__1513 (
            .O(N__7750),
            .I(N__7728));
    InMux I__1512 (
            .O(N__7747),
            .I(N__7728));
    InMux I__1511 (
            .O(N__7744),
            .I(N__7725));
    InMux I__1510 (
            .O(N__7741),
            .I(N__7722));
    InMux I__1509 (
            .O(N__7740),
            .I(N__7716));
    InMux I__1508 (
            .O(N__7737),
            .I(N__7713));
    InMux I__1507 (
            .O(N__7736),
            .I(N__7708));
    InMux I__1506 (
            .O(N__7733),
            .I(N__7708));
    LocalMux I__1505 (
            .O(N__7728),
            .I(N__7705));
    LocalMux I__1504 (
            .O(N__7725),
            .I(N__7700));
    LocalMux I__1503 (
            .O(N__7722),
            .I(N__7700));
    InMux I__1502 (
            .O(N__7721),
            .I(N__7695));
    InMux I__1501 (
            .O(N__7720),
            .I(N__7695));
    InMux I__1500 (
            .O(N__7719),
            .I(N__7692));
    LocalMux I__1499 (
            .O(N__7716),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1498 (
            .O(N__7713),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1497 (
            .O(N__7708),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__1496 (
            .O(N__7705),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__1495 (
            .O(N__7700),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1494 (
            .O(N__7695),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1493 (
            .O(N__7692),
            .I(\U712_CHIP_RAM.N_314 ));
    InMux I__1492 (
            .O(N__7677),
            .I(N__7674));
    LocalMux I__1491 (
            .O(N__7674),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1490 (
            .O(N__7671),
            .I(N__7668));
    LocalMux I__1489 (
            .O(N__7668),
            .I(N__7665));
    Span12Mux_s5_h I__1488 (
            .O(N__7665),
            .I(N__7662));
    Span12Mux_h I__1487 (
            .O(N__7662),
            .I(N__7659));
    Odrv12 I__1486 (
            .O(N__7659),
            .I(CMA_c_7));
    CEMux I__1485 (
            .O(N__7656),
            .I(N__7651));
    CEMux I__1484 (
            .O(N__7655),
            .I(N__7647));
    CEMux I__1483 (
            .O(N__7654),
            .I(N__7644));
    LocalMux I__1482 (
            .O(N__7651),
            .I(N__7640));
    CEMux I__1481 (
            .O(N__7650),
            .I(N__7637));
    LocalMux I__1480 (
            .O(N__7647),
            .I(N__7634));
    LocalMux I__1479 (
            .O(N__7644),
            .I(N__7631));
    CEMux I__1478 (
            .O(N__7643),
            .I(N__7628));
    Span4Mux_v I__1477 (
            .O(N__7640),
            .I(N__7625));
    LocalMux I__1476 (
            .O(N__7637),
            .I(N__7622));
    Span4Mux_v I__1475 (
            .O(N__7634),
            .I(N__7619));
    Span4Mux_v I__1474 (
            .O(N__7631),
            .I(N__7616));
    LocalMux I__1473 (
            .O(N__7628),
            .I(N__7609));
    Span4Mux_v I__1472 (
            .O(N__7625),
            .I(N__7609));
    Span4Mux_h I__1471 (
            .O(N__7622),
            .I(N__7609));
    Odrv4 I__1470 (
            .O(N__7619),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1469 (
            .O(N__7616),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1468 (
            .O(N__7609),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    InMux I__1467 (
            .O(N__7602),
            .I(N__7599));
    LocalMux I__1466 (
            .O(N__7599),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1465 (
            .O(N__7596),
            .I(N__7593));
    LocalMux I__1464 (
            .O(N__7593),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__1463 (
            .O(N__7590),
            .I(N__7587));
    LocalMux I__1462 (
            .O(N__7587),
            .I(N__7584));
    Span4Mux_h I__1461 (
            .O(N__7584),
            .I(N__7581));
    Span4Mux_v I__1460 (
            .O(N__7581),
            .I(N__7578));
    Sp12to4 I__1459 (
            .O(N__7578),
            .I(N__7575));
    Span12Mux_h I__1458 (
            .O(N__7575),
            .I(N__7572));
    Odrv12 I__1457 (
            .O(N__7572),
            .I(A_c_6));
    InMux I__1456 (
            .O(N__7569),
            .I(N__7566));
    LocalMux I__1455 (
            .O(N__7566),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CEMux I__1454 (
            .O(N__7563),
            .I(N__7560));
    LocalMux I__1453 (
            .O(N__7560),
            .I(N__7555));
    CEMux I__1452 (
            .O(N__7559),
            .I(N__7552));
    CEMux I__1451 (
            .O(N__7558),
            .I(N__7548));
    Span4Mux_h I__1450 (
            .O(N__7555),
            .I(N__7543));
    LocalMux I__1449 (
            .O(N__7552),
            .I(N__7543));
    CEMux I__1448 (
            .O(N__7551),
            .I(N__7540));
    LocalMux I__1447 (
            .O(N__7548),
            .I(N__7537));
    Span4Mux_v I__1446 (
            .O(N__7543),
            .I(N__7534));
    LocalMux I__1445 (
            .O(N__7540),
            .I(N__7531));
    Odrv12 I__1444 (
            .O(N__7537),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__1443 (
            .O(N__7534),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__1442 (
            .O(N__7531),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    InMux I__1441 (
            .O(N__7524),
            .I(N__7520));
    InMux I__1440 (
            .O(N__7523),
            .I(N__7517));
    LocalMux I__1439 (
            .O(N__7520),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1438 (
            .O(N__7517),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1437 (
            .O(N__7512),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1436 (
            .O(N__7509),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__1435 (
            .O(N__7506),
            .I(N__7502));
    InMux I__1434 (
            .O(N__7505),
            .I(N__7499));
    LocalMux I__1433 (
            .O(N__7502),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1432 (
            .O(N__7499),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__1431 (
            .O(N__7494),
            .I(N__7467));
    ClkMux I__1430 (
            .O(N__7493),
            .I(N__7467));
    ClkMux I__1429 (
            .O(N__7492),
            .I(N__7467));
    ClkMux I__1428 (
            .O(N__7491),
            .I(N__7467));
    ClkMux I__1427 (
            .O(N__7490),
            .I(N__7467));
    ClkMux I__1426 (
            .O(N__7489),
            .I(N__7467));
    ClkMux I__1425 (
            .O(N__7488),
            .I(N__7467));
    ClkMux I__1424 (
            .O(N__7487),
            .I(N__7467));
    ClkMux I__1423 (
            .O(N__7486),
            .I(N__7467));
    GlobalMux I__1422 (
            .O(N__7467),
            .I(N__7464));
    gio2CtrlBuf I__1421 (
            .O(N__7464),
            .I(C1_c_g));
    SRMux I__1420 (
            .O(N__7461),
            .I(N__7458));
    LocalMux I__1419 (
            .O(N__7458),
            .I(N__7455));
    Odrv12 I__1418 (
            .O(N__7455),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1417 (
            .O(N__7452),
            .I(N__7449));
    LocalMux I__1416 (
            .O(N__7449),
            .I(N__7445));
    InMux I__1415 (
            .O(N__7448),
            .I(N__7442));
    Span4Mux_h I__1414 (
            .O(N__7445),
            .I(N__7435));
    LocalMux I__1413 (
            .O(N__7442),
            .I(N__7435));
    InMux I__1412 (
            .O(N__7441),
            .I(N__7432));
    InMux I__1411 (
            .O(N__7440),
            .I(N__7429));
    Odrv4 I__1410 (
            .O(N__7435),
            .I(DMA_CYCLEm));
    LocalMux I__1409 (
            .O(N__7432),
            .I(DMA_CYCLEm));
    LocalMux I__1408 (
            .O(N__7429),
            .I(DMA_CYCLEm));
    IoInMux I__1407 (
            .O(N__7422),
            .I(N__7419));
    LocalMux I__1406 (
            .O(N__7419),
            .I(N__7416));
    Sp12to4 I__1405 (
            .O(N__7416),
            .I(N__7411));
    InMux I__1404 (
            .O(N__7415),
            .I(N__7408));
    InMux I__1403 (
            .O(N__7414),
            .I(N__7405));
    Span12Mux_v I__1402 (
            .O(N__7411),
            .I(N__7401));
    LocalMux I__1401 (
            .O(N__7408),
            .I(N__7396));
    LocalMux I__1400 (
            .O(N__7405),
            .I(N__7396));
    InMux I__1399 (
            .O(N__7404),
            .I(N__7393));
    Odrv12 I__1398 (
            .O(N__7401),
            .I(DBENn_c));
    Odrv4 I__1397 (
            .O(N__7396),
            .I(DBENn_c));
    LocalMux I__1396 (
            .O(N__7393),
            .I(DBENn_c));
    InMux I__1395 (
            .O(N__7386),
            .I(N__7383));
    LocalMux I__1394 (
            .O(N__7383),
            .I(N__7380));
    Odrv12 I__1393 (
            .O(N__7380),
            .I(\U712_REG_SM.N_402 ));
    InMux I__1392 (
            .O(N__7377),
            .I(N__7373));
    InMux I__1391 (
            .O(N__7376),
            .I(N__7370));
    LocalMux I__1390 (
            .O(N__7373),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__1389 (
            .O(N__7370),
            .I(\U712_REG_SM.START_RSTZ0 ));
    IoInMux I__1388 (
            .O(N__7365),
            .I(N__7361));
    InMux I__1387 (
            .O(N__7364),
            .I(N__7358));
    LocalMux I__1386 (
            .O(N__7361),
            .I(N__7355));
    LocalMux I__1385 (
            .O(N__7358),
            .I(N__7352));
    Span4Mux_s2_v I__1384 (
            .O(N__7355),
            .I(N__7349));
    Span4Mux_v I__1383 (
            .O(N__7352),
            .I(N__7346));
    Span4Mux_h I__1382 (
            .O(N__7349),
            .I(N__7343));
    Span4Mux_v I__1381 (
            .O(N__7346),
            .I(N__7340));
    Odrv4 I__1380 (
            .O(N__7343),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1379 (
            .O(N__7340),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1378 (
            .O(N__7335),
            .I(N__7332));
    LocalMux I__1377 (
            .O(N__7332),
            .I(N__7329));
    Span4Mux_s2_v I__1376 (
            .O(N__7329),
            .I(N__7326));
    Span4Mux_v I__1375 (
            .O(N__7326),
            .I(N__7323));
    Span4Mux_h I__1374 (
            .O(N__7323),
            .I(N__7320));
    Span4Mux_h I__1373 (
            .O(N__7320),
            .I(N__7317));
    Odrv4 I__1372 (
            .O(N__7317),
            .I(CRCSn_c));
    InMux I__1371 (
            .O(N__7314),
            .I(N__7311));
    LocalMux I__1370 (
            .O(N__7311),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1369 (
            .O(N__7308),
            .I(N__7305));
    LocalMux I__1368 (
            .O(N__7305),
            .I(N__7302));
    Span4Mux_s0_v I__1367 (
            .O(N__7302),
            .I(N__7299));
    Sp12to4 I__1366 (
            .O(N__7299),
            .I(N__7296));
    Span12Mux_h I__1365 (
            .O(N__7296),
            .I(N__7293));
    Odrv12 I__1364 (
            .O(N__7293),
            .I(CMA_c_0));
    IoInMux I__1363 (
            .O(N__7290),
            .I(N__7286));
    IoInMux I__1362 (
            .O(N__7289),
            .I(N__7282));
    LocalMux I__1361 (
            .O(N__7286),
            .I(N__7279));
    IoInMux I__1360 (
            .O(N__7285),
            .I(N__7276));
    LocalMux I__1359 (
            .O(N__7282),
            .I(N__7273));
    Span4Mux_s1_v I__1358 (
            .O(N__7279),
            .I(N__7270));
    LocalMux I__1357 (
            .O(N__7276),
            .I(N__7267));
    IoSpan4Mux I__1356 (
            .O(N__7273),
            .I(N__7264));
    Sp12to4 I__1355 (
            .O(N__7270),
            .I(N__7261));
    Span4Mux_s2_h I__1354 (
            .O(N__7267),
            .I(N__7258));
    Span4Mux_s0_v I__1353 (
            .O(N__7264),
            .I(N__7255));
    Span12Mux_h I__1352 (
            .O(N__7261),
            .I(N__7252));
    Sp12to4 I__1351 (
            .O(N__7258),
            .I(N__7249));
    Sp12to4 I__1350 (
            .O(N__7255),
            .I(N__7246));
    Span12Mux_v I__1349 (
            .O(N__7252),
            .I(N__7238));
    Span12Mux_v I__1348 (
            .O(N__7249),
            .I(N__7238));
    Span12Mux_v I__1347 (
            .O(N__7246),
            .I(N__7238));
    InMux I__1346 (
            .O(N__7245),
            .I(N__7235));
    Odrv12 I__1345 (
            .O(N__7238),
            .I(TACK_OUTn));
    LocalMux I__1344 (
            .O(N__7235),
            .I(TACK_OUTn));
    InMux I__1343 (
            .O(N__7230),
            .I(N__7227));
    LocalMux I__1342 (
            .O(N__7227),
            .I(N__7224));
    Odrv12 I__1341 (
            .O(N__7224),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1340 (
            .O(N__7221),
            .I(N__7218));
    LocalMux I__1339 (
            .O(N__7218),
            .I(N__7215));
    Odrv4 I__1338 (
            .O(N__7215),
            .I(\U712_CHIP_RAM.N_367 ));
    InMux I__1337 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1336 (
            .O(N__7209),
            .I(N__7206));
    Span4Mux_v I__1335 (
            .O(N__7206),
            .I(N__7203));
    Odrv4 I__1334 (
            .O(N__7203),
            .I(\U712_CHIP_RAM.N_419 ));
    CascadeMux I__1333 (
            .O(N__7200),
            .I(N__7197));
    InMux I__1332 (
            .O(N__7197),
            .I(N__7193));
    InMux I__1331 (
            .O(N__7196),
            .I(N__7189));
    LocalMux I__1330 (
            .O(N__7193),
            .I(N__7186));
    InMux I__1329 (
            .O(N__7192),
            .I(N__7183));
    LocalMux I__1328 (
            .O(N__7189),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__1327 (
            .O(N__7186),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1326 (
            .O(N__7183),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__1325 (
            .O(N__7176),
            .I(N__7173));
    LocalMux I__1324 (
            .O(N__7173),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1323 (
            .O(N__7170),
            .I(bfn_10_10_0_));
    InMux I__1322 (
            .O(N__7167),
            .I(N__7163));
    InMux I__1321 (
            .O(N__7166),
            .I(N__7160));
    LocalMux I__1320 (
            .O(N__7163),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__1319 (
            .O(N__7160),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1318 (
            .O(N__7155),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1317 (
            .O(N__7152),
            .I(N__7148));
    InMux I__1316 (
            .O(N__7151),
            .I(N__7145));
    LocalMux I__1315 (
            .O(N__7148),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__1314 (
            .O(N__7145),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__1313 (
            .O(N__7140),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1312 (
            .O(N__7137),
            .I(N__7133));
    InMux I__1311 (
            .O(N__7136),
            .I(N__7130));
    LocalMux I__1310 (
            .O(N__7133),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1309 (
            .O(N__7130),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1308 (
            .O(N__7125),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1307 (
            .O(N__7122),
            .I(N__7118));
    InMux I__1306 (
            .O(N__7121),
            .I(N__7115));
    InMux I__1305 (
            .O(N__7118),
            .I(N__7112));
    LocalMux I__1304 (
            .O(N__7115),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1303 (
            .O(N__7112),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1302 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1301 (
            .O(N__7104),
            .I(N__7100));
    InMux I__1300 (
            .O(N__7103),
            .I(N__7097));
    LocalMux I__1299 (
            .O(N__7100),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1298 (
            .O(N__7097),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1297 (
            .O(N__7092),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1296 (
            .O(N__7089),
            .I(N__7086));
    LocalMux I__1295 (
            .O(N__7086),
            .I(N__7083));
    Span4Mux_v I__1294 (
            .O(N__7083),
            .I(N__7080));
    Span4Mux_v I__1293 (
            .O(N__7080),
            .I(N__7077));
    Sp12to4 I__1292 (
            .O(N__7077),
            .I(N__7074));
    Span12Mux_h I__1291 (
            .O(N__7074),
            .I(N__7071));
    Odrv12 I__1290 (
            .O(N__7071),
            .I(A_c_15));
    InMux I__1289 (
            .O(N__7068),
            .I(N__7065));
    LocalMux I__1288 (
            .O(N__7065),
            .I(N__7062));
    Span4Mux_v I__1287 (
            .O(N__7062),
            .I(N__7059));
    Odrv4 I__1286 (
            .O(N__7059),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    CascadeMux I__1285 (
            .O(N__7056),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1284 (
            .O(N__7053),
            .I(N__7050));
    LocalMux I__1283 (
            .O(N__7050),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    InMux I__1282 (
            .O(N__7047),
            .I(N__7044));
    LocalMux I__1281 (
            .O(N__7044),
            .I(N__7041));
    Span12Mux_v I__1280 (
            .O(N__7041),
            .I(N__7038));
    Span12Mux_h I__1279 (
            .O(N__7038),
            .I(N__7035));
    Odrv12 I__1278 (
            .O(N__7035),
            .I(A_c_20));
    InMux I__1277 (
            .O(N__7032),
            .I(N__7028));
    InMux I__1276 (
            .O(N__7031),
            .I(N__7025));
    LocalMux I__1275 (
            .O(N__7028),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    LocalMux I__1274 (
            .O(N__7025),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__1273 (
            .O(N__7020),
            .I(N__7014));
    InMux I__1272 (
            .O(N__7019),
            .I(N__7014));
    LocalMux I__1271 (
            .O(N__7014),
            .I(N__7011));
    Odrv4 I__1270 (
            .O(N__7011),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    InMux I__1269 (
            .O(N__7008),
            .I(N__7005));
    LocalMux I__1268 (
            .O(N__7005),
            .I(\U712_CHIP_RAM.N_435 ));
    InMux I__1267 (
            .O(N__7002),
            .I(N__6999));
    LocalMux I__1266 (
            .O(N__6999),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ));
    CascadeMux I__1265 (
            .O(N__6996),
            .I(N__6992));
    CascadeMux I__1264 (
            .O(N__6995),
            .I(N__6989));
    InMux I__1263 (
            .O(N__6992),
            .I(N__6983));
    InMux I__1262 (
            .O(N__6989),
            .I(N__6980));
    CascadeMux I__1261 (
            .O(N__6988),
            .I(N__6976));
    CascadeMux I__1260 (
            .O(N__6987),
            .I(N__6973));
    CascadeMux I__1259 (
            .O(N__6986),
            .I(N__6970));
    LocalMux I__1258 (
            .O(N__6983),
            .I(N__6967));
    LocalMux I__1257 (
            .O(N__6980),
            .I(N__6964));
    InMux I__1256 (
            .O(N__6979),
            .I(N__6957));
    InMux I__1255 (
            .O(N__6976),
            .I(N__6957));
    InMux I__1254 (
            .O(N__6973),
            .I(N__6957));
    InMux I__1253 (
            .O(N__6970),
            .I(N__6954));
    Odrv4 I__1252 (
            .O(N__6967),
            .I(\U712_CHIP_RAM.N_467 ));
    Odrv4 I__1251 (
            .O(N__6964),
            .I(\U712_CHIP_RAM.N_467 ));
    LocalMux I__1250 (
            .O(N__6957),
            .I(\U712_CHIP_RAM.N_467 ));
    LocalMux I__1249 (
            .O(N__6954),
            .I(\U712_CHIP_RAM.N_467 ));
    InMux I__1248 (
            .O(N__6945),
            .I(N__6942));
    LocalMux I__1247 (
            .O(N__6942),
            .I(N__6939));
    Span4Mux_h I__1246 (
            .O(N__6939),
            .I(N__6936));
    Odrv4 I__1245 (
            .O(N__6936),
            .I(\U712_CHIP_RAM.DBENn_7_0_0 ));
    InMux I__1244 (
            .O(N__6933),
            .I(N__6929));
    InMux I__1243 (
            .O(N__6932),
            .I(N__6926));
    LocalMux I__1242 (
            .O(N__6929),
            .I(N__6922));
    LocalMux I__1241 (
            .O(N__6926),
            .I(N__6919));
    InMux I__1240 (
            .O(N__6925),
            .I(N__6916));
    Span4Mux_v I__1239 (
            .O(N__6922),
            .I(N__6913));
    Span4Mux_v I__1238 (
            .O(N__6919),
            .I(N__6910));
    LocalMux I__1237 (
            .O(N__6916),
            .I(N__6907));
    Sp12to4 I__1236 (
            .O(N__6913),
            .I(N__6902));
    Sp12to4 I__1235 (
            .O(N__6910),
            .I(N__6902));
    Span12Mux_h I__1234 (
            .O(N__6907),
            .I(N__6899));
    Span12Mux_h I__1233 (
            .O(N__6902),
            .I(N__6896));
    Span12Mux_v I__1232 (
            .O(N__6899),
            .I(N__6893));
    Span12Mux_v I__1231 (
            .O(N__6896),
            .I(N__6890));
    Odrv12 I__1230 (
            .O(N__6893),
            .I(AWEn_c));
    Odrv12 I__1229 (
            .O(N__6890),
            .I(AWEn_c));
    InMux I__1228 (
            .O(N__6885),
            .I(N__6880));
    InMux I__1227 (
            .O(N__6884),
            .I(N__6877));
    InMux I__1226 (
            .O(N__6883),
            .I(N__6874));
    LocalMux I__1225 (
            .O(N__6880),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__1224 (
            .O(N__6877),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__1223 (
            .O(N__6874),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    IoInMux I__1222 (
            .O(N__6867),
            .I(N__6864));
    LocalMux I__1221 (
            .O(N__6864),
            .I(N__6861));
    IoSpan4Mux I__1220 (
            .O(N__6861),
            .I(N__6858));
    Sp12to4 I__1219 (
            .O(N__6858),
            .I(N__6855));
    Span12Mux_s7_v I__1218 (
            .O(N__6855),
            .I(N__6851));
    InMux I__1217 (
            .O(N__6854),
            .I(N__6848));
    Odrv12 I__1216 (
            .O(N__6851),
            .I(DBDIR_c));
    LocalMux I__1215 (
            .O(N__6848),
            .I(DBDIR_c));
    InMux I__1214 (
            .O(N__6843),
            .I(N__6840));
    LocalMux I__1213 (
            .O(N__6840),
            .I(\U712_CHIP_RAM.N_361 ));
    IoInMux I__1212 (
            .O(N__6837),
            .I(N__6834));
    LocalMux I__1211 (
            .O(N__6834),
            .I(N__6831));
    Span4Mux_s3_h I__1210 (
            .O(N__6831),
            .I(N__6828));
    Span4Mux_v I__1209 (
            .O(N__6828),
            .I(N__6825));
    Span4Mux_v I__1208 (
            .O(N__6825),
            .I(N__6822));
    Sp12to4 I__1207 (
            .O(N__6822),
            .I(N__6819));
    Span12Mux_s10_h I__1206 (
            .O(N__6819),
            .I(N__6816));
    Odrv12 I__1205 (
            .O(N__6816),
            .I(CMA_c_5));
    IoInMux I__1204 (
            .O(N__6813),
            .I(N__6810));
    LocalMux I__1203 (
            .O(N__6810),
            .I(N__6807));
    Span4Mux_s0_v I__1202 (
            .O(N__6807),
            .I(N__6804));
    Span4Mux_v I__1201 (
            .O(N__6804),
            .I(N__6801));
    Span4Mux_v I__1200 (
            .O(N__6801),
            .I(N__6798));
    Sp12to4 I__1199 (
            .O(N__6798),
            .I(N__6794));
    InMux I__1198 (
            .O(N__6797),
            .I(N__6791));
    Span12Mux_h I__1197 (
            .O(N__6794),
            .I(N__6788));
    LocalMux I__1196 (
            .O(N__6791),
            .I(N__6785));
    Span12Mux_v I__1195 (
            .O(N__6788),
            .I(N__6780));
    Span12Mux_h I__1194 (
            .O(N__6785),
            .I(N__6780));
    Odrv12 I__1193 (
            .O(N__6780),
            .I(A_c_10));
    InMux I__1192 (
            .O(N__6777),
            .I(N__6774));
    LocalMux I__1191 (
            .O(N__6774),
            .I(N__6771));
    Span4Mux_h I__1190 (
            .O(N__6771),
            .I(N__6768));
    Odrv4 I__1189 (
            .O(N__6768),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__1188 (
            .O(N__6765),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__1187 (
            .O(N__6762),
            .I(N__6759));
    LocalMux I__1186 (
            .O(N__6759),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__1185 (
            .O(N__6756),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__1184 (
            .O(N__6753),
            .I(N__6750));
    LocalMux I__1183 (
            .O(N__6750),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1182 (
            .O(N__6747),
            .I(N__6744));
    LocalMux I__1181 (
            .O(N__6744),
            .I(N__6741));
    Span4Mux_s3_v I__1180 (
            .O(N__6741),
            .I(N__6738));
    Span4Mux_v I__1179 (
            .O(N__6738),
            .I(N__6735));
    Span4Mux_v I__1178 (
            .O(N__6735),
            .I(N__6732));
    Odrv4 I__1177 (
            .O(N__6732),
            .I(CMA_c_1));
    InMux I__1176 (
            .O(N__6729),
            .I(N__6726));
    LocalMux I__1175 (
            .O(N__6726),
            .I(N__6723));
    Odrv4 I__1174 (
            .O(N__6723),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1173 (
            .O(N__6720),
            .I(N__6717));
    LocalMux I__1172 (
            .O(N__6717),
            .I(N__6714));
    Span4Mux_v I__1171 (
            .O(N__6714),
            .I(N__6711));
    Sp12to4 I__1170 (
            .O(N__6711),
            .I(N__6708));
    Span12Mux_h I__1169 (
            .O(N__6708),
            .I(N__6705));
    Odrv12 I__1168 (
            .O(N__6705),
            .I(A_c_13));
    InMux I__1167 (
            .O(N__6702),
            .I(N__6699));
    LocalMux I__1166 (
            .O(N__6699),
            .I(N__6696));
    Span4Mux_h I__1165 (
            .O(N__6696),
            .I(N__6693));
    Sp12to4 I__1164 (
            .O(N__6693),
            .I(N__6690));
    Span12Mux_v I__1163 (
            .O(N__6690),
            .I(N__6687));
    Odrv12 I__1162 (
            .O(N__6687),
            .I(A_c_17));
    CascadeMux I__1161 (
            .O(N__6684),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__1160 (
            .O(N__6681),
            .I(N__6678));
    LocalMux I__1159 (
            .O(N__6678),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    InMux I__1158 (
            .O(N__6675),
            .I(N__6672));
    LocalMux I__1157 (
            .O(N__6672),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1156 (
            .O(N__6669),
            .I(N__6666));
    LocalMux I__1155 (
            .O(N__6666),
            .I(N__6663));
    Span4Mux_s0_h I__1154 (
            .O(N__6663),
            .I(N__6660));
    Sp12to4 I__1153 (
            .O(N__6660),
            .I(N__6657));
    Span12Mux_s9_v I__1152 (
            .O(N__6657),
            .I(N__6654));
    Span12Mux_h I__1151 (
            .O(N__6654),
            .I(N__6651));
    Odrv12 I__1150 (
            .O(N__6651),
            .I(CMA_c_3));
    InMux I__1149 (
            .O(N__6648),
            .I(N__6645));
    LocalMux I__1148 (
            .O(N__6645),
            .I(N__6642));
    Span12Mux_v I__1147 (
            .O(N__6642),
            .I(N__6639));
    Span12Mux_h I__1146 (
            .O(N__6639),
            .I(N__6636));
    Odrv12 I__1145 (
            .O(N__6636),
            .I(A_c_14));
    InMux I__1144 (
            .O(N__6633),
            .I(N__6628));
    CascadeMux I__1143 (
            .O(N__6632),
            .I(N__6623));
    InMux I__1142 (
            .O(N__6631),
            .I(N__6620));
    LocalMux I__1141 (
            .O(N__6628),
            .I(N__6617));
    InMux I__1140 (
            .O(N__6627),
            .I(N__6614));
    InMux I__1139 (
            .O(N__6626),
            .I(N__6609));
    InMux I__1138 (
            .O(N__6623),
            .I(N__6609));
    LocalMux I__1137 (
            .O(N__6620),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1136 (
            .O(N__6617),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1135 (
            .O(N__6614),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1134 (
            .O(N__6609),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    CascadeMux I__1133 (
            .O(N__6600),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    InMux I__1132 (
            .O(N__6597),
            .I(N__6593));
    InMux I__1131 (
            .O(N__6596),
            .I(N__6590));
    LocalMux I__1130 (
            .O(N__6593),
            .I(N__6584));
    LocalMux I__1129 (
            .O(N__6590),
            .I(N__6581));
    InMux I__1128 (
            .O(N__6589),
            .I(N__6574));
    InMux I__1127 (
            .O(N__6588),
            .I(N__6574));
    InMux I__1126 (
            .O(N__6587),
            .I(N__6574));
    Odrv4 I__1125 (
            .O(N__6584),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1124 (
            .O(N__6581),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1123 (
            .O(N__6574),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__1122 (
            .O(N__6567),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ));
    InMux I__1121 (
            .O(N__6564),
            .I(N__6560));
    IoInMux I__1120 (
            .O(N__6563),
            .I(N__6557));
    LocalMux I__1119 (
            .O(N__6560),
            .I(N__6554));
    LocalMux I__1118 (
            .O(N__6557),
            .I(N__6551));
    Span4Mux_v I__1117 (
            .O(N__6554),
            .I(N__6548));
    Span12Mux_s4_v I__1116 (
            .O(N__6551),
            .I(N__6545));
    Span4Mux_v I__1115 (
            .O(N__6548),
            .I(N__6542));
    Span12Mux_v I__1114 (
            .O(N__6545),
            .I(N__6537));
    Sp12to4 I__1113 (
            .O(N__6542),
            .I(N__6537));
    Span12Mux_h I__1112 (
            .O(N__6537),
            .I(N__6534));
    Odrv12 I__1111 (
            .O(N__6534),
            .I(A_c_9));
    InMux I__1110 (
            .O(N__6531),
            .I(N__6528));
    LocalMux I__1109 (
            .O(N__6528),
            .I(N__6525));
    Span4Mux_h I__1108 (
            .O(N__6525),
            .I(N__6522));
    Odrv4 I__1107 (
            .O(N__6522),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    CascadeMux I__1106 (
            .O(N__6519),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    InMux I__1105 (
            .O(N__6516),
            .I(N__6513));
    LocalMux I__1104 (
            .O(N__6513),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1103 (
            .O(N__6510),
            .I(N__6507));
    LocalMux I__1102 (
            .O(N__6507),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__1101 (
            .O(N__6504),
            .I(\U712_CHIP_RAM.N_335_cascade_ ));
    IoInMux I__1100 (
            .O(N__6501),
            .I(N__6498));
    LocalMux I__1099 (
            .O(N__6498),
            .I(N__6495));
    Span12Mux_s7_v I__1098 (
            .O(N__6495),
            .I(N__6492));
    Span12Mux_v I__1097 (
            .O(N__6492),
            .I(N__6489));
    Odrv12 I__1096 (
            .O(N__6489),
            .I(N_202_i));
    InMux I__1095 (
            .O(N__6486),
            .I(N__6483));
    LocalMux I__1094 (
            .O(N__6483),
            .I(N__6479));
    InMux I__1093 (
            .O(N__6482),
            .I(N__6476));
    Span4Mux_h I__1092 (
            .O(N__6479),
            .I(N__6471));
    LocalMux I__1091 (
            .O(N__6476),
            .I(N__6471));
    Span4Mux_v I__1090 (
            .O(N__6471),
            .I(N__6468));
    Sp12to4 I__1089 (
            .O(N__6468),
            .I(N__6465));
    Span12Mux_h I__1088 (
            .O(N__6465),
            .I(N__6462));
    Odrv12 I__1087 (
            .O(N__6462),
            .I(TSn_c));
    InMux I__1086 (
            .O(N__6459),
            .I(N__6456));
    LocalMux I__1085 (
            .O(N__6456),
            .I(N__6453));
    Span4Mux_h I__1084 (
            .O(N__6453),
            .I(N__6450));
    Span4Mux_v I__1083 (
            .O(N__6450),
            .I(N__6447));
    Span4Mux_v I__1082 (
            .O(N__6447),
            .I(N__6444));
    Odrv4 I__1081 (
            .O(N__6444),
            .I(RAMSPACEn_c));
    IoInMux I__1080 (
            .O(N__6441),
            .I(N__6438));
    LocalMux I__1079 (
            .O(N__6438),
            .I(N__6435));
    IoSpan4Mux I__1078 (
            .O(N__6435),
            .I(N__6432));
    Span4Mux_s3_v I__1077 (
            .O(N__6432),
            .I(N__6429));
    Span4Mux_v I__1076 (
            .O(N__6429),
            .I(N__6426));
    Odrv4 I__1075 (
            .O(N__6426),
            .I(N_165_i));
    IoInMux I__1074 (
            .O(N__6423),
            .I(N__6420));
    LocalMux I__1073 (
            .O(N__6420),
            .I(N__6417));
    Span4Mux_s2_h I__1072 (
            .O(N__6417),
            .I(N__6414));
    Span4Mux_v I__1071 (
            .O(N__6414),
            .I(N__6411));
    Span4Mux_h I__1070 (
            .O(N__6411),
            .I(N__6408));
    Sp12to4 I__1069 (
            .O(N__6408),
            .I(N__6405));
    Span12Mux_h I__1068 (
            .O(N__6405),
            .I(N__6402));
    Odrv12 I__1067 (
            .O(N__6402),
            .I(WEn_c));
    IoInMux I__1066 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1065 (
            .O(N__6396),
            .I(N__6393));
    Span4Mux_s0_v I__1064 (
            .O(N__6393),
            .I(N__6390));
    Sp12to4 I__1063 (
            .O(N__6390),
            .I(N__6387));
    Span12Mux_h I__1062 (
            .O(N__6387),
            .I(N__6384));
    Odrv12 I__1061 (
            .O(N__6384),
            .I(RASn_c));
    CascadeMux I__1060 (
            .O(N__6381),
            .I(\U712_CHIP_RAM.N_428_cascade_ ));
    InMux I__1059 (
            .O(N__6378),
            .I(N__6373));
    InMux I__1058 (
            .O(N__6377),
            .I(N__6368));
    InMux I__1057 (
            .O(N__6376),
            .I(N__6368));
    LocalMux I__1056 (
            .O(N__6373),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__1055 (
            .O(N__6368),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    SRMux I__1054 (
            .O(N__6363),
            .I(N__6359));
    SRMux I__1053 (
            .O(N__6362),
            .I(N__6356));
    LocalMux I__1052 (
            .O(N__6359),
            .I(N__6353));
    LocalMux I__1051 (
            .O(N__6356),
            .I(N__6350));
    Odrv4 I__1050 (
            .O(N__6353),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    Odrv4 I__1049 (
            .O(N__6350),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    InMux I__1048 (
            .O(N__6345),
            .I(N__6342));
    LocalMux I__1047 (
            .O(N__6342),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__1046 (
            .O(N__6339),
            .I(N__6333));
    InMux I__1045 (
            .O(N__6338),
            .I(N__6333));
    LocalMux I__1044 (
            .O(N__6333),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__1043 (
            .O(N__6330),
            .I(N__6327));
    LocalMux I__1042 (
            .O(N__6327),
            .I(\U712_CHIP_RAM.N_430 ));
    CascadeMux I__1041 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ));
    InMux I__1040 (
            .O(N__6321),
            .I(N__6318));
    LocalMux I__1039 (
            .O(N__6318),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__1038 (
            .O(N__6315),
            .I(N__6312));
    InMux I__1037 (
            .O(N__6312),
            .I(N__6308));
    CascadeMux I__1036 (
            .O(N__6311),
            .I(N__6304));
    LocalMux I__1035 (
            .O(N__6308),
            .I(N__6301));
    InMux I__1034 (
            .O(N__6307),
            .I(N__6296));
    InMux I__1033 (
            .O(N__6304),
            .I(N__6296));
    Odrv12 I__1032 (
            .O(N__6301),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1031 (
            .O(N__6296),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1030 (
            .O(N__6291),
            .I(N__6288));
    LocalMux I__1029 (
            .O(N__6288),
            .I(N__6283));
    InMux I__1028 (
            .O(N__6287),
            .I(N__6278));
    InMux I__1027 (
            .O(N__6286),
            .I(N__6278));
    Odrv4 I__1026 (
            .O(N__6283),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1025 (
            .O(N__6278),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__1024 (
            .O(N__6273),
            .I(\U712_CHIP_RAM.N_435_cascade_ ));
    CascadeMux I__1023 (
            .O(N__6270),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ));
    CEMux I__1022 (
            .O(N__6267),
            .I(N__6264));
    LocalMux I__1021 (
            .O(N__6264),
            .I(N__6261));
    Odrv12 I__1020 (
            .O(N__6261),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ));
    InMux I__1019 (
            .O(N__6258),
            .I(N__6255));
    LocalMux I__1018 (
            .O(N__6255),
            .I(N__6251));
    InMux I__1017 (
            .O(N__6254),
            .I(N__6248));
    Span4Mux_h I__1016 (
            .O(N__6251),
            .I(N__6245));
    LocalMux I__1015 (
            .O(N__6248),
            .I(\U712_CHIP_RAM.N_325 ));
    Odrv4 I__1014 (
            .O(N__6245),
            .I(\U712_CHIP_RAM.N_325 ));
    InMux I__1013 (
            .O(N__6240),
            .I(N__6236));
    InMux I__1012 (
            .O(N__6239),
            .I(N__6233));
    LocalMux I__1011 (
            .O(N__6236),
            .I(N__6230));
    LocalMux I__1010 (
            .O(N__6233),
            .I(\U712_CHIP_RAM.N_321 ));
    Odrv4 I__1009 (
            .O(N__6230),
            .I(\U712_CHIP_RAM.N_321 ));
    InMux I__1008 (
            .O(N__6225),
            .I(N__6217));
    CascadeMux I__1007 (
            .O(N__6224),
            .I(N__6206));
    CascadeMux I__1006 (
            .O(N__6223),
            .I(N__6203));
    InMux I__1005 (
            .O(N__6222),
            .I(N__6191));
    InMux I__1004 (
            .O(N__6221),
            .I(N__6191));
    InMux I__1003 (
            .O(N__6220),
            .I(N__6188));
    LocalMux I__1002 (
            .O(N__6217),
            .I(N__6185));
    InMux I__1001 (
            .O(N__6216),
            .I(N__6182));
    InMux I__1000 (
            .O(N__6215),
            .I(N__6173));
    InMux I__999 (
            .O(N__6214),
            .I(N__6173));
    InMux I__998 (
            .O(N__6213),
            .I(N__6173));
    InMux I__997 (
            .O(N__6212),
            .I(N__6173));
    InMux I__996 (
            .O(N__6211),
            .I(N__6168));
    InMux I__995 (
            .O(N__6210),
            .I(N__6168));
    InMux I__994 (
            .O(N__6209),
            .I(N__6160));
    InMux I__993 (
            .O(N__6206),
            .I(N__6155));
    InMux I__992 (
            .O(N__6203),
            .I(N__6155));
    InMux I__991 (
            .O(N__6202),
            .I(N__6150));
    InMux I__990 (
            .O(N__6201),
            .I(N__6150));
    InMux I__989 (
            .O(N__6200),
            .I(N__6139));
    InMux I__988 (
            .O(N__6199),
            .I(N__6139));
    InMux I__987 (
            .O(N__6198),
            .I(N__6139));
    InMux I__986 (
            .O(N__6197),
            .I(N__6139));
    InMux I__985 (
            .O(N__6196),
            .I(N__6139));
    LocalMux I__984 (
            .O(N__6191),
            .I(N__6136));
    LocalMux I__983 (
            .O(N__6188),
            .I(N__6125));
    Span4Mux_v I__982 (
            .O(N__6185),
            .I(N__6125));
    LocalMux I__981 (
            .O(N__6182),
            .I(N__6125));
    LocalMux I__980 (
            .O(N__6173),
            .I(N__6125));
    LocalMux I__979 (
            .O(N__6168),
            .I(N__6125));
    InMux I__978 (
            .O(N__6167),
            .I(N__6114));
    InMux I__977 (
            .O(N__6166),
            .I(N__6114));
    InMux I__976 (
            .O(N__6165),
            .I(N__6114));
    InMux I__975 (
            .O(N__6164),
            .I(N__6114));
    InMux I__974 (
            .O(N__6163),
            .I(N__6114));
    LocalMux I__973 (
            .O(N__6160),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__972 (
            .O(N__6155),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__971 (
            .O(N__6150),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__970 (
            .O(N__6139),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__969 (
            .O(N__6136),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__968 (
            .O(N__6125),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__967 (
            .O(N__6114),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__966 (
            .O(N__6099),
            .I(N__6090));
    InMux I__965 (
            .O(N__6098),
            .I(N__6085));
    CascadeMux I__964 (
            .O(N__6097),
            .I(N__6082));
    CascadeMux I__963 (
            .O(N__6096),
            .I(N__6078));
    CascadeMux I__962 (
            .O(N__6095),
            .I(N__6074));
    CascadeMux I__961 (
            .O(N__6094),
            .I(N__6071));
    CascadeMux I__960 (
            .O(N__6093),
            .I(N__6066));
    InMux I__959 (
            .O(N__6090),
            .I(N__6063));
    CascadeMux I__958 (
            .O(N__6089),
            .I(N__6057));
    InMux I__957 (
            .O(N__6088),
            .I(N__6054));
    LocalMux I__956 (
            .O(N__6085),
            .I(N__6051));
    InMux I__955 (
            .O(N__6082),
            .I(N__6040));
    InMux I__954 (
            .O(N__6081),
            .I(N__6040));
    InMux I__953 (
            .O(N__6078),
            .I(N__6040));
    InMux I__952 (
            .O(N__6077),
            .I(N__6040));
    InMux I__951 (
            .O(N__6074),
            .I(N__6031));
    InMux I__950 (
            .O(N__6071),
            .I(N__6031));
    InMux I__949 (
            .O(N__6070),
            .I(N__6031));
    InMux I__948 (
            .O(N__6069),
            .I(N__6031));
    InMux I__947 (
            .O(N__6066),
            .I(N__6018));
    LocalMux I__946 (
            .O(N__6063),
            .I(N__6015));
    InMux I__945 (
            .O(N__6062),
            .I(N__6008));
    InMux I__944 (
            .O(N__6061),
            .I(N__6008));
    InMux I__943 (
            .O(N__6060),
            .I(N__6008));
    InMux I__942 (
            .O(N__6057),
            .I(N__6005));
    LocalMux I__941 (
            .O(N__6054),
            .I(N__6000));
    Span4Mux_h I__940 (
            .O(N__6051),
            .I(N__6000));
    InMux I__939 (
            .O(N__6050),
            .I(N__5995));
    InMux I__938 (
            .O(N__6049),
            .I(N__5995));
    LocalMux I__937 (
            .O(N__6040),
            .I(N__5990));
    LocalMux I__936 (
            .O(N__6031),
            .I(N__5990));
    InMux I__935 (
            .O(N__6030),
            .I(N__5983));
    InMux I__934 (
            .O(N__6029),
            .I(N__5983));
    InMux I__933 (
            .O(N__6028),
            .I(N__5983));
    InMux I__932 (
            .O(N__6027),
            .I(N__5976));
    InMux I__931 (
            .O(N__6026),
            .I(N__5976));
    InMux I__930 (
            .O(N__6025),
            .I(N__5976));
    InMux I__929 (
            .O(N__6024),
            .I(N__5967));
    InMux I__928 (
            .O(N__6023),
            .I(N__5967));
    InMux I__927 (
            .O(N__6022),
            .I(N__5967));
    InMux I__926 (
            .O(N__6021),
            .I(N__5967));
    LocalMux I__925 (
            .O(N__6018),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__924 (
            .O(N__6015),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__923 (
            .O(N__6008),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__922 (
            .O(N__6005),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__921 (
            .O(N__6000),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__920 (
            .O(N__5995),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__919 (
            .O(N__5990),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__918 (
            .O(N__5983),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__917 (
            .O(N__5976),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__916 (
            .O(N__5967),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__915 (
            .O(N__5946),
            .I(N__5942));
    InMux I__914 (
            .O(N__5945),
            .I(N__5938));
    LocalMux I__913 (
            .O(N__5942),
            .I(N__5935));
    InMux I__912 (
            .O(N__5941),
            .I(N__5932));
    LocalMux I__911 (
            .O(N__5938),
            .I(\U712_CHIP_RAM.N_551 ));
    Odrv4 I__910 (
            .O(N__5935),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__909 (
            .O(N__5932),
            .I(\U712_CHIP_RAM.N_551 ));
    CascadeMux I__908 (
            .O(N__5925),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ));
    InMux I__907 (
            .O(N__5922),
            .I(N__5919));
    LocalMux I__906 (
            .O(N__5919),
            .I(N__5916));
    Span4Mux_h I__905 (
            .O(N__5916),
            .I(N__5913));
    Odrv4 I__904 (
            .O(N__5913),
            .I(\U712_CHIP_RAM.LATCH_CLK_6 ));
    IoInMux I__903 (
            .O(N__5910),
            .I(N__5906));
    IoInMux I__902 (
            .O(N__5909),
            .I(N__5903));
    LocalMux I__901 (
            .O(N__5906),
            .I(N__5898));
    LocalMux I__900 (
            .O(N__5903),
            .I(N__5898));
    IoSpan4Mux I__899 (
            .O(N__5898),
            .I(N__5895));
    IoSpan4Mux I__898 (
            .O(N__5895),
            .I(N__5892));
    Sp12to4 I__897 (
            .O(N__5892),
            .I(N__5889));
    Span12Mux_s6_v I__896 (
            .O(N__5889),
            .I(N__5885));
    InMux I__895 (
            .O(N__5888),
            .I(N__5882));
    Odrv12 I__894 (
            .O(N__5885),
            .I(RAMENn_c));
    LocalMux I__893 (
            .O(N__5882),
            .I(RAMENn_c));
    InMux I__892 (
            .O(N__5877),
            .I(N__5873));
    CascadeMux I__891 (
            .O(N__5876),
            .I(N__5868));
    LocalMux I__890 (
            .O(N__5873),
            .I(N__5865));
    CascadeMux I__889 (
            .O(N__5872),
            .I(N__5861));
    InMux I__888 (
            .O(N__5871),
            .I(N__5854));
    InMux I__887 (
            .O(N__5868),
            .I(N__5851));
    Span4Mux_v I__886 (
            .O(N__5865),
            .I(N__5848));
    InMux I__885 (
            .O(N__5864),
            .I(N__5843));
    InMux I__884 (
            .O(N__5861),
            .I(N__5843));
    InMux I__883 (
            .O(N__5860),
            .I(N__5836));
    InMux I__882 (
            .O(N__5859),
            .I(N__5836));
    InMux I__881 (
            .O(N__5858),
            .I(N__5836));
    InMux I__880 (
            .O(N__5857),
            .I(N__5833));
    LocalMux I__879 (
            .O(N__5854),
            .I(N__5830));
    LocalMux I__878 (
            .O(N__5851),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__877 (
            .O(N__5848),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__876 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__875 (
            .O(N__5836),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__874 (
            .O(N__5833),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__873 (
            .O(N__5830),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__872 (
            .O(N__5817),
            .I(N__5813));
    InMux I__871 (
            .O(N__5816),
            .I(N__5810));
    LocalMux I__870 (
            .O(N__5813),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    LocalMux I__869 (
            .O(N__5810),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    IoInMux I__868 (
            .O(N__5805),
            .I(N__5802));
    LocalMux I__867 (
            .O(N__5802),
            .I(N__5799));
    IoSpan4Mux I__866 (
            .O(N__5799),
            .I(N__5796));
    Span4Mux_s0_v I__865 (
            .O(N__5796),
            .I(N__5793));
    Sp12to4 I__864 (
            .O(N__5793),
            .I(N__5789));
    InMux I__863 (
            .O(N__5792),
            .I(N__5786));
    Span12Mux_s8_v I__862 (
            .O(N__5789),
            .I(N__5783));
    LocalMux I__861 (
            .O(N__5786),
            .I(N__5780));
    Span12Mux_v I__860 (
            .O(N__5783),
            .I(N__5777));
    Span4Mux_v I__859 (
            .O(N__5780),
            .I(N__5774));
    Span12Mux_h I__858 (
            .O(N__5777),
            .I(N__5769));
    Sp12to4 I__857 (
            .O(N__5774),
            .I(N__5769));
    Odrv12 I__856 (
            .O(N__5769),
            .I(A_c_11));
    InMux I__855 (
            .O(N__5766),
            .I(N__5763));
    LocalMux I__854 (
            .O(N__5763),
            .I(N__5760));
    Odrv4 I__853 (
            .O(N__5760),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__852 (
            .O(N__5757),
            .I(N__5753));
    InMux I__851 (
            .O(N__5756),
            .I(N__5750));
    LocalMux I__850 (
            .O(N__5753),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    LocalMux I__849 (
            .O(N__5750),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    InMux I__848 (
            .O(N__5745),
            .I(N__5742));
    LocalMux I__847 (
            .O(N__5742),
            .I(\U712_CHIP_RAM.m93_i_a2_5 ));
    CascadeMux I__846 (
            .O(N__5739),
            .I(N__5736));
    InMux I__845 (
            .O(N__5736),
            .I(N__5733));
    LocalMux I__844 (
            .O(N__5733),
            .I(N__5727));
    CascadeMux I__843 (
            .O(N__5732),
            .I(N__5724));
    InMux I__842 (
            .O(N__5731),
            .I(N__5719));
    InMux I__841 (
            .O(N__5730),
            .I(N__5719));
    Span4Mux_h I__840 (
            .O(N__5727),
            .I(N__5716));
    InMux I__839 (
            .O(N__5724),
            .I(N__5713));
    LocalMux I__838 (
            .O(N__5719),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    Odrv4 I__837 (
            .O(N__5716),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    LocalMux I__836 (
            .O(N__5713),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    InMux I__835 (
            .O(N__5706),
            .I(N__5703));
    LocalMux I__834 (
            .O(N__5703),
            .I(\U712_CHIP_RAM.m93_i_a2_4 ));
    IoInMux I__833 (
            .O(N__5700),
            .I(N__5697));
    LocalMux I__832 (
            .O(N__5697),
            .I(N__5694));
    Span12Mux_s7_h I__831 (
            .O(N__5694),
            .I(N__5691));
    Span12Mux_h I__830 (
            .O(N__5691),
            .I(N__5688));
    Odrv12 I__829 (
            .O(N__5688),
            .I(CMA_c_8));
    InMux I__828 (
            .O(N__5685),
            .I(N__5682));
    LocalMux I__827 (
            .O(N__5682),
            .I(N__5679));
    Odrv4 I__826 (
            .O(N__5679),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__825 (
            .O(N__5676),
            .I(N__5673));
    LocalMux I__824 (
            .O(N__5673),
            .I(N__5670));
    Span4Mux_v I__823 (
            .O(N__5670),
            .I(N__5667));
    Span4Mux_v I__822 (
            .O(N__5667),
            .I(N__5664));
    Span4Mux_v I__821 (
            .O(N__5664),
            .I(N__5661));
    Sp12to4 I__820 (
            .O(N__5661),
            .I(N__5658));
    Odrv12 I__819 (
            .O(N__5658),
            .I(A_c_19));
    IoInMux I__818 (
            .O(N__5655),
            .I(N__5652));
    LocalMux I__817 (
            .O(N__5652),
            .I(N__5649));
    Span12Mux_s7_h I__816 (
            .O(N__5649),
            .I(N__5646));
    Span12Mux_h I__815 (
            .O(N__5646),
            .I(N__5643));
    Odrv12 I__814 (
            .O(N__5643),
            .I(CMA_c_9));
    InMux I__813 (
            .O(N__5640),
            .I(N__5637));
    LocalMux I__812 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.m123_i_2 ));
    CascadeMux I__811 (
            .O(N__5634),
            .I(N__5630));
    InMux I__810 (
            .O(N__5633),
            .I(N__5626));
    InMux I__809 (
            .O(N__5630),
            .I(N__5623));
    InMux I__808 (
            .O(N__5629),
            .I(N__5620));
    LocalMux I__807 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__806 (
            .O(N__5623),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__805 (
            .O(N__5620),
            .I(\U712_CHIP_RAM.N_305 ));
    InMux I__804 (
            .O(N__5613),
            .I(N__5610));
    LocalMux I__803 (
            .O(N__5610),
            .I(\U712_CHIP_RAM.N_190 ));
    InMux I__802 (
            .O(N__5607),
            .I(N__5604));
    LocalMux I__801 (
            .O(N__5604),
            .I(N__5600));
    InMux I__800 (
            .O(N__5603),
            .I(N__5597));
    Odrv4 I__799 (
            .O(N__5600),
            .I(\U712_CHIP_RAM.N_476 ));
    LocalMux I__798 (
            .O(N__5597),
            .I(\U712_CHIP_RAM.N_476 ));
    InMux I__797 (
            .O(N__5592),
            .I(N__5589));
    LocalMux I__796 (
            .O(N__5589),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ));
    InMux I__795 (
            .O(N__5586),
            .I(N__5583));
    LocalMux I__794 (
            .O(N__5583),
            .I(\U712_CHIP_RAM.N_344 ));
    CascadeMux I__793 (
            .O(N__5580),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ));
    InMux I__792 (
            .O(N__5577),
            .I(N__5573));
    InMux I__791 (
            .O(N__5576),
            .I(N__5568));
    LocalMux I__790 (
            .O(N__5573),
            .I(N__5565));
    InMux I__789 (
            .O(N__5572),
            .I(N__5562));
    InMux I__788 (
            .O(N__5571),
            .I(N__5559));
    LocalMux I__787 (
            .O(N__5568),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__786 (
            .O(N__5565),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__785 (
            .O(N__5562),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__784 (
            .O(N__5559),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__783 (
            .O(N__5550),
            .I(N__5539));
    CascadeMux I__782 (
            .O(N__5549),
            .I(N__5536));
    InMux I__781 (
            .O(N__5548),
            .I(N__5533));
    InMux I__780 (
            .O(N__5547),
            .I(N__5528));
    InMux I__779 (
            .O(N__5546),
            .I(N__5528));
    InMux I__778 (
            .O(N__5545),
            .I(N__5525));
    CascadeMux I__777 (
            .O(N__5544),
            .I(N__5520));
    InMux I__776 (
            .O(N__5543),
            .I(N__5517));
    InMux I__775 (
            .O(N__5542),
            .I(N__5510));
    InMux I__774 (
            .O(N__5539),
            .I(N__5510));
    InMux I__773 (
            .O(N__5536),
            .I(N__5510));
    LocalMux I__772 (
            .O(N__5533),
            .I(N__5507));
    LocalMux I__771 (
            .O(N__5528),
            .I(N__5504));
    LocalMux I__770 (
            .O(N__5525),
            .I(N__5498));
    InMux I__769 (
            .O(N__5524),
            .I(N__5495));
    InMux I__768 (
            .O(N__5523),
            .I(N__5492));
    InMux I__767 (
            .O(N__5520),
            .I(N__5489));
    LocalMux I__766 (
            .O(N__5517),
            .I(N__5484));
    LocalMux I__765 (
            .O(N__5510),
            .I(N__5484));
    Span4Mux_v I__764 (
            .O(N__5507),
            .I(N__5479));
    Span4Mux_v I__763 (
            .O(N__5504),
            .I(N__5479));
    InMux I__762 (
            .O(N__5503),
            .I(N__5474));
    InMux I__761 (
            .O(N__5502),
            .I(N__5474));
    InMux I__760 (
            .O(N__5501),
            .I(N__5471));
    Span4Mux_h I__759 (
            .O(N__5498),
            .I(N__5468));
    LocalMux I__758 (
            .O(N__5495),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__757 (
            .O(N__5492),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__756 (
            .O(N__5489),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__755 (
            .O(N__5484),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__754 (
            .O(N__5479),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__753 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__752 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__751 (
            .O(N__5468),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__750 (
            .O(N__5451),
            .I(N__5447));
    InMux I__749 (
            .O(N__5450),
            .I(N__5437));
    LocalMux I__748 (
            .O(N__5447),
            .I(N__5434));
    CascadeMux I__747 (
            .O(N__5446),
            .I(N__5429));
    InMux I__746 (
            .O(N__5445),
            .I(N__5425));
    InMux I__745 (
            .O(N__5444),
            .I(N__5422));
    InMux I__744 (
            .O(N__5443),
            .I(N__5410));
    InMux I__743 (
            .O(N__5442),
            .I(N__5410));
    InMux I__742 (
            .O(N__5441),
            .I(N__5410));
    InMux I__741 (
            .O(N__5440),
            .I(N__5410));
    LocalMux I__740 (
            .O(N__5437),
            .I(N__5407));
    Span4Mux_v I__739 (
            .O(N__5434),
            .I(N__5404));
    InMux I__738 (
            .O(N__5433),
            .I(N__5401));
    InMux I__737 (
            .O(N__5432),
            .I(N__5398));
    InMux I__736 (
            .O(N__5429),
            .I(N__5395));
    InMux I__735 (
            .O(N__5428),
            .I(N__5392));
    LocalMux I__734 (
            .O(N__5425),
            .I(N__5387));
    LocalMux I__733 (
            .O(N__5422),
            .I(N__5387));
    InMux I__732 (
            .O(N__5421),
            .I(N__5382));
    InMux I__731 (
            .O(N__5420),
            .I(N__5382));
    InMux I__730 (
            .O(N__5419),
            .I(N__5379));
    LocalMux I__729 (
            .O(N__5410),
            .I(N__5374));
    Span4Mux_h I__728 (
            .O(N__5407),
            .I(N__5374));
    Odrv4 I__727 (
            .O(N__5404),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__726 (
            .O(N__5401),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__725 (
            .O(N__5398),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__724 (
            .O(N__5395),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__723 (
            .O(N__5392),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__722 (
            .O(N__5387),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__721 (
            .O(N__5382),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__720 (
            .O(N__5379),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__719 (
            .O(N__5374),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__718 (
            .O(N__5355),
            .I(N__5349));
    InMux I__717 (
            .O(N__5354),
            .I(N__5343));
    InMux I__716 (
            .O(N__5353),
            .I(N__5343));
    InMux I__715 (
            .O(N__5352),
            .I(N__5340));
    LocalMux I__714 (
            .O(N__5349),
            .I(N__5336));
    InMux I__713 (
            .O(N__5348),
            .I(N__5333));
    LocalMux I__712 (
            .O(N__5343),
            .I(N__5328));
    LocalMux I__711 (
            .O(N__5340),
            .I(N__5328));
    InMux I__710 (
            .O(N__5339),
            .I(N__5325));
    Odrv4 I__709 (
            .O(N__5336),
            .I(\U712_CHIP_RAM.N_307 ));
    LocalMux I__708 (
            .O(N__5333),
            .I(\U712_CHIP_RAM.N_307 ));
    Odrv4 I__707 (
            .O(N__5328),
            .I(\U712_CHIP_RAM.N_307 ));
    LocalMux I__706 (
            .O(N__5325),
            .I(\U712_CHIP_RAM.N_307 ));
    CascadeMux I__705 (
            .O(N__5316),
            .I(\U712_CHIP_RAM.N_551_cascade_ ));
    CascadeMux I__704 (
            .O(N__5313),
            .I(N__5310));
    InMux I__703 (
            .O(N__5310),
            .I(N__5307));
    LocalMux I__702 (
            .O(N__5307),
            .I(N__5302));
    InMux I__701 (
            .O(N__5306),
            .I(N__5299));
    InMux I__700 (
            .O(N__5305),
            .I(N__5296));
    Odrv4 I__699 (
            .O(N__5302),
            .I(\U712_CHIP_RAM.N_304 ));
    LocalMux I__698 (
            .O(N__5299),
            .I(\U712_CHIP_RAM.N_304 ));
    LocalMux I__697 (
            .O(N__5296),
            .I(\U712_CHIP_RAM.N_304 ));
    CascadeMux I__696 (
            .O(N__5289),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ));
    InMux I__695 (
            .O(N__5286),
            .I(N__5283));
    LocalMux I__694 (
            .O(N__5283),
            .I(\U712_CHIP_RAM.N_378 ));
    InMux I__693 (
            .O(N__5280),
            .I(N__5271));
    InMux I__692 (
            .O(N__5279),
            .I(N__5271));
    InMux I__691 (
            .O(N__5278),
            .I(N__5271));
    LocalMux I__690 (
            .O(N__5271),
            .I(N__5267));
    InMux I__689 (
            .O(N__5270),
            .I(N__5263));
    Span4Mux_h I__688 (
            .O(N__5267),
            .I(N__5260));
    InMux I__687 (
            .O(N__5266),
            .I(N__5257));
    LocalMux I__686 (
            .O(N__5263),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__685 (
            .O(N__5260),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__684 (
            .O(N__5257),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__683 (
            .O(N__5250),
            .I(N__5247));
    InMux I__682 (
            .O(N__5247),
            .I(N__5242));
    InMux I__681 (
            .O(N__5246),
            .I(N__5237));
    InMux I__680 (
            .O(N__5245),
            .I(N__5237));
    LocalMux I__679 (
            .O(N__5242),
            .I(N__5231));
    LocalMux I__678 (
            .O(N__5237),
            .I(N__5231));
    InMux I__677 (
            .O(N__5236),
            .I(N__5227));
    Span4Mux_h I__676 (
            .O(N__5231),
            .I(N__5224));
    InMux I__675 (
            .O(N__5230),
            .I(N__5221));
    LocalMux I__674 (
            .O(N__5227),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv4 I__673 (
            .O(N__5224),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__672 (
            .O(N__5221),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__671 (
            .O(N__5214),
            .I(N__5205));
    InMux I__670 (
            .O(N__5213),
            .I(N__5205));
    InMux I__669 (
            .O(N__5212),
            .I(N__5205));
    LocalMux I__668 (
            .O(N__5205),
            .I(\U712_CHIP_RAM.SDRAM_CMDs_0_4 ));
    CascadeMux I__667 (
            .O(N__5202),
            .I(\U712_CHIP_RAM.N_396_cascade_ ));
    InMux I__666 (
            .O(N__5199),
            .I(N__5196));
    LocalMux I__665 (
            .O(N__5196),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_0_2 ));
    InMux I__664 (
            .O(N__5193),
            .I(N__5190));
    LocalMux I__663 (
            .O(N__5190),
            .I(\U712_CHIP_RAM.N_397 ));
    InMux I__662 (
            .O(N__5187),
            .I(N__5184));
    LocalMux I__661 (
            .O(N__5184),
            .I(N__5181));
    Span4Mux_h I__660 (
            .O(N__5181),
            .I(N__5178));
    Odrv4 I__659 (
            .O(N__5178),
            .I(\U712_CHIP_RAM.N_555 ));
    InMux I__658 (
            .O(N__5175),
            .I(N__5172));
    LocalMux I__657 (
            .O(N__5172),
            .I(N__5169));
    Span4Mux_h I__656 (
            .O(N__5169),
            .I(N__5166));
    Odrv4 I__655 (
            .O(N__5166),
            .I(\U712_CHIP_RAM.N_449 ));
    CascadeMux I__654 (
            .O(N__5163),
            .I(N__5160));
    InMux I__653 (
            .O(N__5160),
            .I(N__5154));
    InMux I__652 (
            .O(N__5159),
            .I(N__5154));
    LocalMux I__651 (
            .O(N__5154),
            .I(N__5151));
    Span4Mux_h I__650 (
            .O(N__5151),
            .I(N__5148));
    Odrv4 I__649 (
            .O(N__5148),
            .I(\U712_CHIP_RAM.SDRAM_CMDs_0_1 ));
    InMux I__648 (
            .O(N__5145),
            .I(N__5142));
    LocalMux I__647 (
            .O(N__5142),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_3 ));
    CEMux I__646 (
            .O(N__5139),
            .I(N__5136));
    LocalMux I__645 (
            .O(N__5136),
            .I(N__5133));
    Span4Mux_v I__644 (
            .O(N__5133),
            .I(N__5130));
    Odrv4 I__643 (
            .O(N__5130),
            .I(\U712_CHIP_RAM.N_194_0 ));
    InMux I__642 (
            .O(N__5127),
            .I(N__5124));
    LocalMux I__641 (
            .O(N__5124),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa ));
    CascadeMux I__640 (
            .O(N__5121),
            .I(N__5117));
    InMux I__639 (
            .O(N__5120),
            .I(N__5105));
    InMux I__638 (
            .O(N__5117),
            .I(N__5105));
    InMux I__637 (
            .O(N__5116),
            .I(N__5099));
    InMux I__636 (
            .O(N__5115),
            .I(N__5099));
    InMux I__635 (
            .O(N__5114),
            .I(N__5094));
    InMux I__634 (
            .O(N__5113),
            .I(N__5094));
    InMux I__633 (
            .O(N__5112),
            .I(N__5091));
    InMux I__632 (
            .O(N__5111),
            .I(N__5080));
    InMux I__631 (
            .O(N__5110),
            .I(N__5080));
    LocalMux I__630 (
            .O(N__5105),
            .I(N__5077));
    InMux I__629 (
            .O(N__5104),
            .I(N__5074));
    LocalMux I__628 (
            .O(N__5099),
            .I(N__5069));
    LocalMux I__627 (
            .O(N__5094),
            .I(N__5069));
    LocalMux I__626 (
            .O(N__5091),
            .I(N__5066));
    InMux I__625 (
            .O(N__5090),
            .I(N__5061));
    InMux I__624 (
            .O(N__5089),
            .I(N__5061));
    InMux I__623 (
            .O(N__5088),
            .I(N__5054));
    InMux I__622 (
            .O(N__5087),
            .I(N__5054));
    InMux I__621 (
            .O(N__5086),
            .I(N__5054));
    InMux I__620 (
            .O(N__5085),
            .I(N__5051));
    LocalMux I__619 (
            .O(N__5080),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__618 (
            .O(N__5077),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__617 (
            .O(N__5074),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__616 (
            .O(N__5069),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__615 (
            .O(N__5066),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__614 (
            .O(N__5061),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__613 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__612 (
            .O(N__5051),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__611 (
            .O(N__5034),
            .I(N__5031));
    LocalMux I__610 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    IoInMux I__609 (
            .O(N__5028),
            .I(N__5025));
    LocalMux I__608 (
            .O(N__5025),
            .I(N__5022));
    IoSpan4Mux I__607 (
            .O(N__5022),
            .I(N__5019));
    Sp12to4 I__606 (
            .O(N__5019),
            .I(N__5016));
    Span12Mux_s7_h I__605 (
            .O(N__5016),
            .I(N__5013));
    Span12Mux_h I__604 (
            .O(N__5013),
            .I(N__5010));
    Odrv12 I__603 (
            .O(N__5010),
            .I(CMA_c_6));
    InMux I__602 (
            .O(N__5007),
            .I(N__5004));
    LocalMux I__601 (
            .O(N__5004),
            .I(N__5001));
    Sp12to4 I__600 (
            .O(N__5001),
            .I(N__4998));
    Span12Mux_v I__599 (
            .O(N__4998),
            .I(N__4995));
    Span12Mux_h I__598 (
            .O(N__4995),
            .I(N__4992));
    Odrv12 I__597 (
            .O(N__4992),
            .I(A_c_12));
    InMux I__596 (
            .O(N__4989),
            .I(N__4986));
    LocalMux I__595 (
            .O(N__4986),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    CascadeMux I__594 (
            .O(N__4983),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__593 (
            .O(N__4980),
            .I(N__4977));
    LocalMux I__592 (
            .O(N__4977),
            .I(N__4974));
    Sp12to4 I__591 (
            .O(N__4974),
            .I(N__4971));
    Span12Mux_v I__590 (
            .O(N__4971),
            .I(N__4968));
    Span12Mux_h I__589 (
            .O(N__4968),
            .I(N__4965));
    Odrv12 I__588 (
            .O(N__4965),
            .I(A_c_16));
    InMux I__587 (
            .O(N__4962),
            .I(N__4959));
    LocalMux I__586 (
            .O(N__4959),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    IoInMux I__585 (
            .O(N__4956),
            .I(N__4953));
    LocalMux I__584 (
            .O(N__4953),
            .I(N__4950));
    Span4Mux_s1_v I__583 (
            .O(N__4950),
            .I(N__4947));
    Span4Mux_v I__582 (
            .O(N__4947),
            .I(N__4944));
    Span4Mux_v I__581 (
            .O(N__4944),
            .I(N__4941));
    Odrv4 I__580 (
            .O(N__4941),
            .I(VBENn_c));
    InMux I__579 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__578 (
            .O(N__4935),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_6 ));
    InMux I__577 (
            .O(N__4932),
            .I(N__4928));
    InMux I__576 (
            .O(N__4931),
            .I(N__4925));
    LocalMux I__575 (
            .O(N__4928),
            .I(\U712_CHIP_RAM.N_194 ));
    LocalMux I__574 (
            .O(N__4925),
            .I(\U712_CHIP_RAM.N_194 ));
    CascadeMux I__573 (
            .O(N__4920),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ));
    InMux I__572 (
            .O(N__4917),
            .I(N__4914));
    LocalMux I__571 (
            .O(N__4914),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1 ));
    InMux I__570 (
            .O(N__4911),
            .I(N__4908));
    LocalMux I__569 (
            .O(N__4908),
            .I(N__4903));
    CascadeMux I__568 (
            .O(N__4907),
            .I(N__4900));
    InMux I__567 (
            .O(N__4906),
            .I(N__4897));
    Span4Mux_h I__566 (
            .O(N__4903),
            .I(N__4894));
    InMux I__565 (
            .O(N__4900),
            .I(N__4891));
    LocalMux I__564 (
            .O(N__4897),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    Odrv4 I__563 (
            .O(N__4894),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__562 (
            .O(N__4891),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__561 (
            .O(N__4884),
            .I(N__4881));
    LocalMux I__560 (
            .O(N__4881),
            .I(N__4877));
    InMux I__559 (
            .O(N__4880),
            .I(N__4873));
    Span4Mux_h I__558 (
            .O(N__4877),
            .I(N__4870));
    InMux I__557 (
            .O(N__4876),
            .I(N__4867));
    LocalMux I__556 (
            .O(N__4873),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__555 (
            .O(N__4870),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__554 (
            .O(N__4867),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__553 (
            .O(N__4860),
            .I(N__4855));
    InMux I__552 (
            .O(N__4859),
            .I(N__4852));
    InMux I__551 (
            .O(N__4858),
            .I(N__4849));
    InMux I__550 (
            .O(N__4855),
            .I(N__4846));
    LocalMux I__549 (
            .O(N__4852),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    LocalMux I__548 (
            .O(N__4849),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    LocalMux I__547 (
            .O(N__4846),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    InMux I__546 (
            .O(N__4839),
            .I(N__4835));
    InMux I__545 (
            .O(N__4838),
            .I(N__4832));
    LocalMux I__544 (
            .O(N__4835),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    LocalMux I__543 (
            .O(N__4832),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    InMux I__542 (
            .O(N__4827),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ));
    InMux I__541 (
            .O(N__4824),
            .I(N__4820));
    InMux I__540 (
            .O(N__4823),
            .I(N__4817));
    LocalMux I__539 (
            .O(N__4820),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    LocalMux I__538 (
            .O(N__4817),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    InMux I__537 (
            .O(N__4812),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ));
    InMux I__536 (
            .O(N__4809),
            .I(N__4805));
    InMux I__535 (
            .O(N__4808),
            .I(N__4802));
    LocalMux I__534 (
            .O(N__4805),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    LocalMux I__533 (
            .O(N__4802),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    InMux I__532 (
            .O(N__4797),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ));
    InMux I__531 (
            .O(N__4794),
            .I(N__4790));
    InMux I__530 (
            .O(N__4793),
            .I(N__4787));
    LocalMux I__529 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    LocalMux I__528 (
            .O(N__4787),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    InMux I__527 (
            .O(N__4782),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ));
    InMux I__526 (
            .O(N__4779),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ));
    InMux I__525 (
            .O(N__4776),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ));
    InMux I__524 (
            .O(N__4773),
            .I(N__4769));
    InMux I__523 (
            .O(N__4772),
            .I(N__4766));
    LocalMux I__522 (
            .O(N__4769),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    LocalMux I__521 (
            .O(N__4766),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    InMux I__520 (
            .O(N__4761),
            .I(N__4757));
    InMux I__519 (
            .O(N__4760),
            .I(N__4754));
    LocalMux I__518 (
            .O(N__4757),
            .I(N__4751));
    LocalMux I__517 (
            .O(N__4754),
            .I(N__4748));
    Span4Mux_v I__516 (
            .O(N__4751),
            .I(N__4745));
    Span4Mux_v I__515 (
            .O(N__4748),
            .I(N__4742));
    Sp12to4 I__514 (
            .O(N__4745),
            .I(N__4737));
    Sp12to4 I__513 (
            .O(N__4742),
            .I(N__4737));
    Span12Mux_h I__512 (
            .O(N__4737),
            .I(N__4734));
    Span12Mux_v I__511 (
            .O(N__4734),
            .I(N__4731));
    Odrv12 I__510 (
            .O(N__4731),
            .I(DBRn_c));
    CascadeMux I__509 (
            .O(N__4728),
            .I(\U712_CHIP_RAM.N_307_cascade_ ));
    CascadeMux I__508 (
            .O(N__4725),
            .I(\U712_CHIP_RAM.N_467_cascade_ ));
    CascadeMux I__507 (
            .O(N__4722),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__506 (
            .O(N__4719),
            .I(N__4716));
    LocalMux I__505 (
            .O(N__4716),
            .I(N__4713));
    Span4Mux_h I__504 (
            .O(N__4713),
            .I(N__4710));
    Odrv4 I__503 (
            .O(N__4710),
            .I(\U712_CHIP_RAM.N_440 ));
    CascadeMux I__502 (
            .O(N__4707),
            .I(\U712_CHIP_RAM.N_304_cascade_ ));
    CascadeMux I__501 (
            .O(N__4704),
            .I(\U712_CHIP_RAM.N_312_cascade_ ));
    CascadeMux I__500 (
            .O(N__4701),
            .I(N__4698));
    InMux I__499 (
            .O(N__4698),
            .I(N__4695));
    LocalMux I__498 (
            .O(N__4695),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__497 (
            .O(N__4692),
            .I(N__4679));
    InMux I__496 (
            .O(N__4691),
            .I(N__4679));
    InMux I__495 (
            .O(N__4690),
            .I(N__4679));
    InMux I__494 (
            .O(N__4689),
            .I(N__4676));
    InMux I__493 (
            .O(N__4688),
            .I(N__4669));
    InMux I__492 (
            .O(N__4687),
            .I(N__4669));
    InMux I__491 (
            .O(N__4686),
            .I(N__4669));
    LocalMux I__490 (
            .O(N__4679),
            .I(\U712_CHIP_RAM.N_39 ));
    LocalMux I__489 (
            .O(N__4676),
            .I(\U712_CHIP_RAM.N_39 ));
    LocalMux I__488 (
            .O(N__4669),
            .I(\U712_CHIP_RAM.N_39 ));
    InMux I__487 (
            .O(N__4662),
            .I(N__4659));
    LocalMux I__486 (
            .O(N__4659),
            .I(N__4655));
    InMux I__485 (
            .O(N__4658),
            .I(N__4652));
    Sp12to4 I__484 (
            .O(N__4655),
            .I(N__4649));
    LocalMux I__483 (
            .O(N__4652),
            .I(\U712_CHIP_RAM.N_326 ));
    Odrv12 I__482 (
            .O(N__4649),
            .I(\U712_CHIP_RAM.N_326 ));
    CascadeMux I__481 (
            .O(N__4644),
            .I(\U712_CHIP_RAM.N_39_cascade_ ));
    CEMux I__480 (
            .O(N__4641),
            .I(N__4638));
    LocalMux I__479 (
            .O(N__4638),
            .I(N__4634));
    CEMux I__478 (
            .O(N__4637),
            .I(N__4631));
    Sp12to4 I__477 (
            .O(N__4634),
            .I(N__4626));
    LocalMux I__476 (
            .O(N__4631),
            .I(N__4626));
    Odrv12 I__475 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__474 (
            .O(N__4623),
            .I(N__4620));
    InMux I__473 (
            .O(N__4620),
            .I(N__4616));
    InMux I__472 (
            .O(N__4619),
            .I(N__4613));
    LocalMux I__471 (
            .O(N__4616),
            .I(\U712_CHIP_RAM.N_20_0 ));
    LocalMux I__470 (
            .O(N__4613),
            .I(\U712_CHIP_RAM.N_20_0 ));
    InMux I__469 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__468 (
            .O(N__4605),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ));
    InMux I__467 (
            .O(N__4602),
            .I(N__4599));
    LocalMux I__466 (
            .O(N__4599),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    InMux I__465 (
            .O(N__4596),
            .I(N__4593));
    LocalMux I__464 (
            .O(N__4593),
            .I(\U712_CHIP_RAM.m101_i_1 ));
    CascadeMux I__463 (
            .O(N__4590),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    InMux I__462 (
            .O(N__4587),
            .I(N__4584));
    LocalMux I__461 (
            .O(N__4584),
            .I(\U712_CHIP_RAM.N_376 ));
    CascadeMux I__460 (
            .O(N__4581),
            .I(\U712_CHIP_RAM.m101_i_0_cascade_ ));
    InMux I__459 (
            .O(N__4578),
            .I(N__4575));
    LocalMux I__458 (
            .O(N__4575),
            .I(\U712_CHIP_RAM.m101_i_2 ));
    InMux I__457 (
            .O(N__4572),
            .I(N__4569));
    LocalMux I__456 (
            .O(N__4569),
            .I(N__4566));
    Span12Mux_v I__455 (
            .O(N__4566),
            .I(N__4563));
    Odrv12 I__454 (
            .O(N__4563),
            .I(A_c_5));
    InMux I__453 (
            .O(N__4560),
            .I(N__4557));
    LocalMux I__452 (
            .O(N__4557),
            .I(N__4554));
    Span4Mux_h I__451 (
            .O(N__4554),
            .I(N__4551));
    Sp12to4 I__450 (
            .O(N__4551),
            .I(N__4548));
    Span12Mux_v I__449 (
            .O(N__4548),
            .I(N__4545));
    Odrv12 I__448 (
            .O(N__4545),
            .I(A_c_18));
    CascadeMux I__447 (
            .O(N__4542),
            .I(\U712_CHIP_RAM.N_436_cascade_ ));
    CascadeMux I__446 (
            .O(N__4539),
            .I(\U712_CHIP_RAM.N_194_cascade_ ));
    InMux I__445 (
            .O(N__4536),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__444 (
            .O(N__4533),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__443 (
            .O(N__4530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__442 (
            .O(N__4527),
            .I(N__4524));
    LocalMux I__441 (
            .O(N__4524),
            .I(N__4521));
    Span4Mux_v I__440 (
            .O(N__4521),
            .I(N__4518));
    Sp12to4 I__439 (
            .O(N__4518),
            .I(N__4515));
    Odrv12 I__438 (
            .O(N__4515),
            .I(A_c_8));
    InMux I__437 (
            .O(N__4512),
            .I(N__4509));
    LocalMux I__436 (
            .O(N__4509),
            .I(N__4506));
    Span12Mux_h I__435 (
            .O(N__4506),
            .I(N__4503));
    Span12Mux_v I__434 (
            .O(N__4503),
            .I(N__4500));
    Odrv12 I__433 (
            .O(N__4500),
            .I(A_c_2));
    InMux I__432 (
            .O(N__4497),
            .I(N__4494));
    LocalMux I__431 (
            .O(N__4494),
            .I(N__4491));
    Span4Mux_h I__430 (
            .O(N__4491),
            .I(N__4488));
    Sp12to4 I__429 (
            .O(N__4488),
            .I(N__4485));
    Span12Mux_v I__428 (
            .O(N__4485),
            .I(N__4482));
    Odrv12 I__427 (
            .O(N__4482),
            .I(A_c_3));
    InMux I__426 (
            .O(N__4479),
            .I(N__4476));
    LocalMux I__425 (
            .O(N__4476),
            .I(N__4473));
    Span4Mux_v I__424 (
            .O(N__4473),
            .I(N__4470));
    Span4Mux_v I__423 (
            .O(N__4470),
            .I(N__4467));
    Sp12to4 I__422 (
            .O(N__4467),
            .I(N__4464));
    Odrv12 I__421 (
            .O(N__4464),
            .I(A_c_4));
    InMux I__420 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__419 (
            .O(N__4458),
            .I(N__4455));
    Span4Mux_v I__418 (
            .O(N__4455),
            .I(N__4452));
    Sp12to4 I__417 (
            .O(N__4452),
            .I(N__4449));
    Odrv12 I__416 (
            .O(N__4449),
            .I(A_c_7));
    IoInMux I__415 (
            .O(N__4446),
            .I(N__4443));
    LocalMux I__414 (
            .O(N__4443),
            .I(N__4440));
    IoSpan4Mux I__413 (
            .O(N__4440),
            .I(N__4437));
    Sp12to4 I__412 (
            .O(N__4437),
            .I(N__4434));
    Span12Mux_s9_h I__411 (
            .O(N__4434),
            .I(N__4431));
    Span12Mux_h I__410 (
            .O(N__4431),
            .I(N__4427));
    InMux I__409 (
            .O(N__4430),
            .I(N__4424));
    Odrv12 I__408 (
            .O(N__4427),
            .I(CLK_EN_c));
    LocalMux I__407 (
            .O(N__4424),
            .I(CLK_EN_c));
    CascadeMux I__406 (
            .O(N__4419),
            .I(\U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ));
    InMux I__405 (
            .O(N__4416),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__404 (
            .O(N__4413),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__403 (
            .O(N__4410),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__402 (
            .O(N__4407),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    IoInMux I__401 (
            .O(N__4404),
            .I(N__4401));
    LocalMux I__400 (
            .O(N__4401),
            .I(N__4398));
    Span4Mux_s3_v I__399 (
            .O(N__4398),
            .I(N__4395));
    Span4Mux_h I__398 (
            .O(N__4395),
            .I(N__4392));
    Odrv4 I__397 (
            .O(N__4392),
            .I(CLK80_PLL_i_i));
    InMux I__396 (
            .O(N__4389),
            .I(N__4386));
    LocalMux I__395 (
            .O(N__4386),
            .I(N__4383));
    Span12Mux_h I__394 (
            .O(N__4383),
            .I(N__4380));
    Span12Mux_v I__393 (
            .O(N__4380),
            .I(N__4377));
    Odrv12 I__392 (
            .O(N__4377),
            .I(REGSPACEn_c));
    CascadeMux I__391 (
            .O(N__4374),
            .I(\U712_CHIP_RAM.N_555_cascade_ ));
    CascadeMux I__390 (
            .O(N__4371),
            .I(\U712_CHIP_RAM.N_390_cascade_ ));
    InMux I__389 (
            .O(N__4368),
            .I(N__4365));
    LocalMux I__388 (
            .O(N__4365),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_0 ));
    CascadeMux I__387 (
            .O(N__4362),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_ ));
    InMux I__386 (
            .O(N__4359),
            .I(N__4356));
    LocalMux I__385 (
            .O(N__4356),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_2 ));
    IoInMux I__384 (
            .O(N__4353),
            .I(N__4350));
    LocalMux I__383 (
            .O(N__4350),
            .I(N__4347));
    Odrv12 I__382 (
            .O(N__4347),
            .I(DBRn_c_i_0));
    IoInMux I__381 (
            .O(N__4344),
            .I(N__4341));
    LocalMux I__380 (
            .O(N__4341),
            .I(N__4338));
    Span4Mux_s0_v I__379 (
            .O(N__4338),
            .I(N__4335));
    Span4Mux_v I__378 (
            .O(N__4335),
            .I(N__4332));
    Sp12to4 I__377 (
            .O(N__4332),
            .I(N__4329));
    Span12Mux_h I__376 (
            .O(N__4329),
            .I(N__4326));
    Span12Mux_v I__375 (
            .O(N__4326),
            .I(N__4323));
    Odrv12 I__374 (
            .O(N__4323),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__7492));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__7491));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__7486));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__7489));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__7493));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__7487));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__7490));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__7494));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__8468),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9195),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4353),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__8169),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_4  (
            .in0(N__9828),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8615),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_0 (
            .in0(N__9993),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__6486),
            .in2(_gnd_net_),
            .in3(N__4389),
            .lcout(\U712_REG_SM.N_402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_7_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_7_5_0 .LUT_INIT=16'b1111000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_7_5_0  (
            .in0(N__5114),
            .in1(N__6199),
            .in2(N__5550),
            .in3(N__6081),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_7_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_7_5_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_7_5_1  (
            .in0(N__6196),
            .in1(N__5441),
            .in2(_gnd_net_),
            .in3(N__5113),
            .lcout(\U712_CHIP_RAM.N_555 ),
            .ltout(\U712_CHIP_RAM.N_555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_7_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_7_5_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_7_5_2  (
            .in0(N__5542),
            .in1(_gnd_net_),
            .in2(N__4374),
            .in3(N__5633),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_7_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_7_5_3 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_7_5_3  (
            .in0(N__5355),
            .in1(_gnd_net_),
            .in2(N__4371),
            .in3(N__4368),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_5_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_5_4 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_7_5_4  (
            .in0(N__4359),
            .in1(N__4932),
            .in2(N__4362),
            .in3(N__7904),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9953),
            .ce(),
            .sr(N__9799));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_5_5 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_5_5  (
            .in0(N__6200),
            .in1(_gnd_net_),
            .in2(N__6097),
            .in3(N__5443),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_6  (
            .in0(N__5440),
            .in1(N__6197),
            .in2(N__5549),
            .in3(N__6077),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDs_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_7_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_7_5_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_7_5_7  (
            .in0(N__6198),
            .in1(_gnd_net_),
            .in2(N__6096),
            .in3(N__5442),
            .lcout(\U712_CHIP_RAM.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_7_6_1 .LUT_INIT=16'b1011111100000100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_7_6_1  (
            .in0(N__5354),
            .in1(N__4608),
            .in2(N__4623),
            .in3(N__4430),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9959),
            .ce(),
            .sr(N__9794));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_6_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_6_4  (
            .in0(N__6240),
            .in1(N__5433),
            .in2(N__6089),
            .in3(N__10946),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_6_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_6_5  (
            .in0(N__5353),
            .in1(N__4619),
            .in2(N__4419),
            .in3(N__5523),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_7_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_7_0  (
            .in0(N__7440),
            .in1(N__5104),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_6 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_7_1  (
            .in0(N__4690),
            .in1(N__5432),
            .in2(_gnd_net_),
            .in3(N__4416),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__6088),
            .in2(_gnd_net_),
            .in3(N__4413),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_7_3  (
            .in0(N__4691),
            .in1(N__5524),
            .in2(_gnd_net_),
            .in3(N__4410),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_7_4  (
            .in0(N__4686),
            .in1(N__5270),
            .in2(_gnd_net_),
            .in3(N__4407),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_7_5  (
            .in0(N__4692),
            .in1(N__4880),
            .in2(_gnd_net_),
            .in3(N__4536),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_7_6  (
            .in0(N__4687),
            .in1(N__5236),
            .in2(_gnd_net_),
            .in3(N__4533),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_7_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_7_7  (
            .in0(N__4906),
            .in1(N__4688),
            .in2(_gnd_net_),
            .in3(N__4530),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(N__4641),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4527),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9972),
            .ce(N__7551),
            .sr(N__9784));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_9_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_9_0  (
            .in0(N__4512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9977),
            .ce(N__7559),
            .sr(N__9774));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4497),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9977),
            .ce(N__7559),
            .sr(N__9774));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4479),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9977),
            .ce(N__7559),
            .sr(N__9774));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_9_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_9_3  (
            .in0(N__4461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9977),
            .ce(N__7559),
            .sr(N__9774));
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_7_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_1_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__5730),
            .in2(_gnd_net_),
            .in3(N__4859),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9982),
            .ce(),
            .sr(N__6363));
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_7_10_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_0_LC_7_10_2  (
            .in0(N__5731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9982),
            .ce(),
            .sr(N__6363));
    defparam DBRn_ibuf_RNIBAB_LC_7_11_1.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_7_11_1 (
            .in0(N__4761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_8_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_8_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_8_4_1  (
            .in0(N__4572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9943),
            .ce(N__7558),
            .sr(N__9800));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4560),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9943),
            .ce(N__7558),
            .sr(N__9800));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_8_5_0 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_8_5_0  (
            .in0(N__6596),
            .in1(N__8334),
            .in2(_gnd_net_),
            .in3(N__6627),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_5_1 .LUT_INIT=16'b0111111101111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_5_1  (
            .in0(N__6201),
            .in1(N__5445),
            .in2(N__6094),
            .in3(N__5115),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_8_5_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9183),
            .in3(N__6070),
            .lcout(\U712_CHIP_RAM.DBENn_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_5_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_5_3  (
            .in0(N__6069),
            .in1(N__6258),
            .in2(_gnd_net_),
            .in3(N__5629),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_5_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_5_4  (
            .in0(N__4578),
            .in1(N__4587),
            .in2(N__4542),
            .in3(N__4596),
            .lcout(\U712_CHIP_RAM.N_194 ),
            .ltout(\U712_CHIP_RAM.N_194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_8_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_8_5_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4539),
            .in3(N__9827),
            .lcout(\U712_CHIP_RAM.N_194_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_8_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_8_5_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_8_5_6  (
            .in0(N__5577),
            .in1(N__10944),
            .in2(_gnd_net_),
            .in3(N__5444),
            .lcout(\U712_CHIP_RAM.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_5_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_5_7  (
            .in0(N__6202),
            .in1(N__5543),
            .in2(N__6095),
            .in3(N__5116),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_6_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_6_0  (
            .in0(N__10409),
            .in1(N__4602),
            .in2(N__8712),
            .in3(N__5613),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9954),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_1  (
            .in0(N__6167),
            .in1(N__10410),
            .in2(_gnd_net_),
            .in3(N__5127),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9954),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_8_6_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_8_6_2  (
            .in0(N__5421),
            .in1(N__6165),
            .in2(_gnd_net_),
            .in3(N__5352),
            .lcout(\U712_CHIP_RAM.m101_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__5420),
            .in2(_gnd_net_),
            .in3(N__5086),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_6_4 .LUT_INIT=16'b1111000000001011;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_6_4  (
            .in0(N__6022),
            .in1(N__5871),
            .in2(N__4590),
            .in3(N__5503),
            .lcout(\U712_CHIP_RAM.N_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_6_5 .LUT_INIT=16'b1100100111001101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_6_5  (
            .in0(N__6166),
            .in1(N__5088),
            .in2(N__5446),
            .in3(N__6024),
            .lcout(\U712_CHIP_RAM.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_6_6 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_6_6  (
            .in0(N__6021),
            .in1(N__6163),
            .in2(N__10418),
            .in3(N__5502),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m101_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_6_7 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_6_7  (
            .in0(N__6164),
            .in1(N__6023),
            .in2(N__4581),
            .in3(N__5087),
            .lcout(\U712_CHIP_RAM.m101_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_7_0 .LUT_INIT=16'b1111010110001111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_7_0  (
            .in0(N__5428),
            .in1(N__5306),
            .in2(N__5544),
            .in3(N__6026),
            .lcout(\U712_CHIP_RAM.m123_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__5571),
            .in2(_gnd_net_),
            .in3(N__5089),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(\U712_CHIP_RAM.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_8_7_2 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_8_7_2  (
            .in0(N__5090),
            .in1(N__6221),
            .in2(N__4707),
            .in3(N__6025),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_8_7_3 .LUT_INIT=16'b1010000011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_8_7_3  (
            .in0(N__5941),
            .in1(_gnd_net_),
            .in2(N__4704),
            .in3(N__10408),
            .lcout(\U712_CHIP_RAM.N_326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_7_4  (
            .in0(N__10407),
            .in1(N__5592),
            .in2(N__4701),
            .in3(N__4689),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9960),
            .ce(N__4637),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_8_7_6 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_8_7_6  (
            .in0(N__4662),
            .in1(N__6222),
            .in2(N__6995),
            .in3(N__6027),
            .lcout(\U712_CHIP_RAM.N_39 ),
            .ltout(\U712_CHIP_RAM.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_7_7  (
            .in0(N__4658),
            .in1(N__5034),
            .in2(N__4644),
            .in3(N__4719),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9960),
            .ce(N__4637),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_8_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_8_0  (
            .in0(N__6254),
            .in1(N__10393),
            .in2(N__5872),
            .in3(N__5603),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_8_1  (
            .in0(N__5230),
            .in1(N__4876),
            .in2(N__4907),
            .in3(N__5266),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(\U712_CHIP_RAM.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_8_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_8_8_2  (
            .in0(N__5501),
            .in1(N__5419),
            .in2(N__4728),
            .in3(N__5085),
            .lcout(\U712_CHIP_RAM.N_467 ),
            .ltout(\U712_CHIP_RAM.N_467_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_3  (
            .in0(N__6212),
            .in1(_gnd_net_),
            .in2(N__4725),
            .in3(N__6028),
            .lcout(\U712_CHIP_RAM.N_476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_8_8_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_8_8_4  (
            .in0(N__6029),
            .in1(N__5816),
            .in2(N__6987),
            .in3(N__6213),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_8_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4722),
            .in3(N__9825),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_8_6  (
            .in0(N__6030),
            .in1(N__6214),
            .in2(N__6988),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_8_7  (
            .in0(N__6215),
            .in1(N__5864),
            .in2(N__6093),
            .in3(N__6979),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9967),
            .ce(N__6267),
            .sr(N__9775));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_8_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_8_9_0  (
            .in0(N__4838),
            .in1(N__4772),
            .in2(N__4860),
            .in3(N__4823),
            .lcout(\U712_CHIP_RAM.m93_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_9_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_9_2  (
            .in0(N__4793),
            .in1(N__4808),
            .in2(_gnd_net_),
            .in3(N__6378),
            .lcout(\U712_CHIP_RAM.m93_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_9_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__5572),
            .in2(_gnd_net_),
            .in3(N__5112),
            .lcout(\U712_CHIP_RAM.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_5 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_9_5  (
            .in0(N__7441),
            .in1(N__6330),
            .in2(N__5876),
            .in3(N__10384),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9973),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_8_10_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_8_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__4858),
            .in2(N__5732),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_10_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_2_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__4839),
            .in2(_gnd_net_),
            .in3(N__4827),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_10_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_3_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__4824),
            .in2(_gnd_net_),
            .in3(N__4812),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_10_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_4_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__4809),
            .in2(_gnd_net_),
            .in3(N__4797),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_10_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_5_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__4794),
            .in2(_gnd_net_),
            .in3(N__4782),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_10_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_6_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__5757),
            .in2(_gnd_net_),
            .in3(N__4779),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_7_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__4773),
            .in2(_gnd_net_),
            .in3(N__4776),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9978),
            .ce(),
            .sr(N__6362));
    defparam DBR_SYNC_0_LC_8_12_7.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_8_12_7.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_8_12_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_8_12_7 (
            .in0(N__4760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9987),
            .ce(),
            .sr(N__9755));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_4_2  (
            .in0(N__5007),
            .in1(N__4989),
            .in2(_gnd_net_),
            .in3(N__8332),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_4_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_9_4_3  (
            .in0(N__8333),
            .in1(N__10947),
            .in2(N__4983),
            .in3(N__9123),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_4_4  (
            .in0(N__4980),
            .in1(N__4962),
            .in2(_gnd_net_),
            .in3(N__8331),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_9_4_6  (
            .in0(N__10948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11897),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_5_0 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_5_0  (
            .in0(N__4917),
            .in1(N__5213),
            .in2(N__5313),
            .in3(N__6220),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_5_1 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_5_1  (
            .in0(N__4938),
            .in1(N__4931),
            .in2(N__4920),
            .in3(N__6631),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9944),
            .ce(),
            .sr(N__9791));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_5_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_5_2  (
            .in0(N__5546),
            .in1(N__5245),
            .in2(_gnd_net_),
            .in3(N__5278),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_9_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__4911),
            .in2(_gnd_net_),
            .in3(N__4884),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDs_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_9_5_4 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_9_5_4  (
            .in0(N__6098),
            .in1(N__5246),
            .in2(N__5121),
            .in3(N__5279),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_9_5_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_9_5_5  (
            .in0(N__5212),
            .in1(N__5547),
            .in2(N__5289),
            .in3(N__5120),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_9_5_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_9_5_6  (
            .in0(N__5286),
            .in1(N__5280),
            .in2(N__5250),
            .in3(N__5214),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_9_6_0 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_9_6_0  (
            .in0(N__6062),
            .in1(N__6209),
            .in2(N__6315),
            .in3(N__5451),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_9_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_9_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_9_6_1  (
            .in0(N__5159),
            .in1(N__5193),
            .in2(N__5202),
            .in3(N__5199),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9947),
            .ce(N__5139),
            .sr(N__9785));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_9_6_2 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_9_6_2  (
            .in0(N__6060),
            .in1(N__5548),
            .in2(N__6223),
            .in3(N__5877),
            .lcout(\U712_CHIP_RAM.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_9_6_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_9_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_9_6_3  (
            .in0(N__5187),
            .in1(N__5175),
            .in2(N__5163),
            .in3(N__5145),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9947),
            .ce(N__5139),
            .sr(N__9785));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_6_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_6_4  (
            .in0(N__6061),
            .in1(N__5946),
            .in2(N__6224),
            .in3(N__5111),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__7364),
            .in2(_gnd_net_),
            .in3(N__5110),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_9_7_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_9_7_2  (
            .in0(N__7787),
            .in1(N__9099),
            .in2(N__7757),
            .in3(N__7053),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(N__7654),
            .sr(N__9776));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_4 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_9_7_4  (
            .in0(N__7788),
            .in1(N__9090),
            .in2(N__7758),
            .in3(N__6681),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(N__7654),
            .sr(N__9776));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_9_7_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_9_7_5  (
            .in0(N__5685),
            .in1(N__5676),
            .in2(N__10945),
            .in3(N__9234),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(N__7654),
            .sr(N__9776));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_7_6 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_7_6  (
            .in0(N__5640),
            .in1(N__6216),
            .in2(N__5634),
            .in3(N__5348),
            .lcout(\U712_CHIP_RAM.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_8_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_8_0  (
            .in0(N__5859),
            .in1(N__6932),
            .in2(_gnd_net_),
            .in3(N__11258),
            .lcout(\U712_CHIP_RAM.N_344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1  (
            .in0(N__5607),
            .in1(N__5817),
            .in2(_gnd_net_),
            .in3(N__5860),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_2  (
            .in0(N__10385),
            .in1(N__5586),
            .in2(N__5580),
            .in3(N__5576),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9961),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_8_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_8_3  (
            .in0(N__5545),
            .in1(N__5450),
            .in2(_gnd_net_),
            .in3(N__5339),
            .lcout(\U712_CHIP_RAM.N_551 ),
            .ltout(\U712_CHIP_RAM.N_551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_8_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_9_8_4  (
            .in0(N__6050),
            .in1(N__6211),
            .in2(N__5316),
            .in3(N__5305),
            .lcout(\U712_CHIP_RAM.N_435 ),
            .ltout(\U712_CHIP_RAM.N_435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_9_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6273),
            .in3(N__6883),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_8_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_8_6  (
            .in0(N__9824),
            .in1(_gnd_net_),
            .in2(N__6270),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_8_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_9_8_7  (
            .in0(N__6210),
            .in1(N__5858),
            .in2(N__6986),
            .in3(N__6049),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1  (
            .in0(N__7192),
            .in1(_gnd_net_),
            .in2(N__6311),
            .in3(N__6376),
            .lcout(\U712_CHIP_RAM.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_2  (
            .in0(N__6239),
            .in1(N__6225),
            .in2(N__6099),
            .in3(N__5945),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_9_9_3  (
            .in0(N__10404),
            .in1(N__5888),
            .in2(N__5925),
            .in3(N__5922),
            .lcout(RAMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9968),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_4  (
            .in0(N__6377),
            .in1(N__6307),
            .in2(N__7200),
            .in3(N__5857),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_5  (
            .in0(N__5792),
            .in1(N__5766),
            .in2(_gnd_net_),
            .in3(N__8358),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_9_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_9_6  (
            .in0(N__5756),
            .in1(N__5745),
            .in2(N__5739),
            .in3(N__5706),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_9_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_9_7  (
            .in0(N__10405),
            .in1(N__8997),
            .in2(N__6381),
            .in3(N__6291),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9968),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__10381),
            .in2(_gnd_net_),
            .in3(N__9021),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9974),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_2  (
            .in0(N__10380),
            .in1(N__8996),
            .in2(_gnd_net_),
            .in3(N__6287),
            .lcout(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3  (
            .in0(N__6339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10382),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9974),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_4  (
            .in0(N__6345),
            .in1(N__6338),
            .in2(_gnd_net_),
            .in3(N__6286),
            .lcout(\U712_CHIP_RAM.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_5  (
            .in0(N__7136),
            .in1(N__7151),
            .in2(N__7122),
            .in3(N__7166),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__7523),
            .in2(_gnd_net_),
            .in3(N__7103),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_10_7 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_10_7  (
            .in0(N__10383),
            .in1(N__7505),
            .in2(N__6324),
            .in3(N__6321),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9974),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_0  (
            .in0(N__10253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6516),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9979),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_4  (
            .in0(N__7415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7448),
            .lcout(\U712_CHIP_RAM.m50_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_11_7 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_9_11_7  (
            .in0(N__11122),
            .in1(N__10252),
            .in2(_gnd_net_),
            .in3(N__11055),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9979),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_1_LC_9_12_1.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_12_1.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_9_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6510),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9983),
            .ce(),
            .sr(N__9754));
    defparam \U712_CHIP_RAM.m37_i_o2_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m37_i_o2_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m37_i_o2_LC_9_14_4 .LUT_INIT=16'b1110110010111011;
    LogicCell40 \U712_CHIP_RAM.m37_i_o2_LC_9_14_4  (
            .in0(N__11688),
            .in1(N__11497),
            .in2(N__11601),
            .in3(N__11358),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_9_14_5 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_9_14_5  (
            .in0(N__11051),
            .in1(N__11747),
            .in2(N__6504),
            .in3(N__10952),
            .lcout(N_202_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__6482),
            .in2(_gnd_net_),
            .in3(N__6459),
            .lcout(\U712_CHIP_RAM.N_419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_165_i_LC_9_19_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_165_i_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_165_i_LC_9_19_0 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.N_165_i_LC_9_19_0  (
            .in0(N__11127),
            .in1(N__11044),
            .in2(_gnd_net_),
            .in3(N__11174),
            .lcout(N_165_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_10_2_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_10_2_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_10_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_10_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6633),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9937),
            .ce(),
            .sr(N__9801));
    defparam \U712_CHIP_RAM.RASn_LC_10_3_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_10_3_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_10_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_10_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6597),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9938),
            .ce(),
            .sr(N__9795));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_10_4_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_10_4_2  (
            .in0(N__7798),
            .in1(N__7830),
            .in2(N__7754),
            .in3(N__6675),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9940),
            .ce(N__7650),
            .sr(N__9792));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_5_0 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_5_0  (
            .in0(N__10949),
            .in1(N__7719),
            .in2(N__8330),
            .in3(N__8202),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_1  (
            .in0(N__6648),
            .in1(N__10950),
            .in2(_gnd_net_),
            .in3(N__9111),
            .lcout(\U712_CHIP_RAM.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_10_5_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__6626),
            .in2(_gnd_net_),
            .in3(N__6589),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_10_5_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_10_5_3  (
            .in0(N__6587),
            .in1(N__8284),
            .in2(N__6632),
            .in3(N__7905),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_5_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_5_4  (
            .in0(N__8285),
            .in1(N__7906),
            .in2(N__6600),
            .in3(N__6588),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_10_5_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6567),
            .in3(N__9826),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_5_6  (
            .in0(N__8286),
            .in1(N__6564),
            .in2(_gnd_net_),
            .in3(N__6531),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_5_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_5_7  (
            .in0(N__8211),
            .in1(N__10951),
            .in2(N__6519),
            .in3(N__8290),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_6_0 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_10_6_0  (
            .in0(N__7721),
            .in1(N__6843),
            .in2(N__8368),
            .in3(N__7221),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(N__7656),
            .sr(N__9777));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_6_4 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_6_4  (
            .in0(N__7720),
            .in1(N__10909),
            .in2(N__8367),
            .in3(N__8198),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_5  (
            .in0(N__6797),
            .in1(N__6777),
            .in2(_gnd_net_),
            .in3(N__8353),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_6_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_6_6  (
            .in0(N__8354),
            .in1(N__10910),
            .in2(N__6765),
            .in3(N__8748),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_6_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__6762),
            .in2(N__6756),
            .in3(N__6753),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(N__7656),
            .sr(N__9777));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_0  (
            .in0(N__10888),
            .in1(N__6729),
            .in2(N__8338),
            .in3(N__9447),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_1  (
            .in0(N__6720),
            .in1(N__7569),
            .in2(_gnd_net_),
            .in3(N__8304),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_7_2  (
            .in0(N__7031),
            .in1(N__8313),
            .in2(_gnd_net_),
            .in3(N__6702),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_7_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_7_3  (
            .in0(N__8315),
            .in1(N__10889),
            .in2(N__6684),
            .in3(N__8595),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_7_4 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_10_7_4  (
            .in0(N__6925),
            .in1(N__11155),
            .in2(N__10406),
            .in3(N__6885),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9948),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_5  (
            .in0(N__7089),
            .in1(N__7068),
            .in2(_gnd_net_),
            .in3(N__8306),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_6  (
            .in0(N__10887),
            .in1(N__8314),
            .in2(N__7056),
            .in3(N__8736),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_10_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__10886),
            .in2(_gnd_net_),
            .in3(N__8305),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_8_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_8_0  (
            .in0(N__7020),
            .in1(N__7047),
            .in2(N__10743),
            .in3(N__7032),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(N__9762));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_10_8_1  (
            .in0(N__10896),
            .in1(N__7019),
            .in2(_gnd_net_),
            .in3(N__7008),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(N__9762));
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_8_2 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_8_2  (
            .in0(N__7002),
            .in1(N__7404),
            .in2(N__6996),
            .in3(N__6945),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(N__9762));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_8_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_8_6  (
            .in0(N__6854),
            .in1(N__6933),
            .in2(_gnd_net_),
            .in3(N__6884),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(N__9762));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7  (
            .in0(N__8648),
            .in1(N__7245),
            .in2(N__7965),
            .in3(N__8574),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(N__9762));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_3  (
            .in0(N__7230),
            .in1(N__10891),
            .in2(_gnd_net_),
            .in3(N__9030),
            .lcout(\U712_CHIP_RAM.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_5 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_5  (
            .in0(N__7212),
            .in1(N__10892),
            .in2(N__10417),
            .in3(N__7196),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9962),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_10_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__7176),
            .in2(_gnd_net_),
            .in3(N__7170),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_10_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__7167),
            .in2(_gnd_net_),
            .in3(N__7155),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_10_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__7152),
            .in2(_gnd_net_),
            .in3(N__7140),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_10_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__7137),
            .in2(_gnd_net_),
            .in3(N__7125),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_10_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__7121),
            .in2(_gnd_net_),
            .in3(N__7107),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_10_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__7104),
            .in2(_gnd_net_),
            .in3(N__7092),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_10_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__7524),
            .in2(_gnd_net_),
            .in3(N__7512),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__7506),
            .in2(_gnd_net_),
            .in3(N__7509),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7488),
            .ce(),
            .sr(N__7461));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_11_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_11_2  (
            .in0(N__7452),
            .in1(N__7414),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.START_RST_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_10_12_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_10_12_1  (
            .in0(N__7376),
            .in1(N__8086),
            .in2(_gnd_net_),
            .in3(N__8785),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9980),
            .ce(),
            .sr(N__9750));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_10_13_5 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_10_13_5  (
            .in0(N__7386),
            .in1(N__7377),
            .in2(N__10419),
            .in3(N__8109),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9984),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_1_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_1_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_1_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_11_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_11_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_11_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7913),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9939),
            .ce(),
            .sr(N__9786));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2  (
            .in0(N__7799),
            .in1(N__9297),
            .in2(N__7753),
            .in3(N__7314),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__7643),
            .sr(N__9778));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_5_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_11_5_3  (
            .in0(N__7914),
            .in1(N__8365),
            .in2(_gnd_net_),
            .in3(N__7736),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__7643),
            .sr(N__9778));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_6  (
            .in0(N__10932),
            .in1(N__7857),
            .in2(N__8370),
            .in3(N__8178),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_5_7  (
            .in0(N__7740),
            .in1(N__7800),
            .in2(N__7845),
            .in3(N__9504),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__7643),
            .sr(N__9778));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_0  (
            .in0(N__9163),
            .in1(N__10741),
            .in2(_gnd_net_),
            .in3(N__9603),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9222),
            .ce(N__10494),
            .sr(N__9766));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_11_7_3  (
            .in0(N__7786),
            .in1(N__8184),
            .in2(N__7755),
            .in3(N__7596),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9946),
            .ce(N__7655),
            .sr(N__9763));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_11_7_4 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_11_7_4  (
            .in0(N__7789),
            .in1(N__9081),
            .in2(N__7756),
            .in3(N__7677),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9946),
            .ce(N__7655),
            .sr(N__9763));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_3  (
            .in0(N__10890),
            .in1(N__7602),
            .in2(N__8369),
            .in3(N__10515),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_11_8_7  (
            .in0(N__7590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9949),
            .ce(N__7563),
            .sr(N__9759));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_0 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_0  (
            .in0(N__7985),
            .in1(N__8641),
            .in2(N__7932),
            .in3(N__8727),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__9756));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_9_3 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_11_9_3  (
            .in0(N__7989),
            .in1(N__8004),
            .in2(_gnd_net_),
            .in3(N__8721),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__9756));
    defparam \U712_REG_SM.REG_TACK_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_9_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_9_5  (
            .in0(N__8066),
            .in1(N__8688),
            .in2(N__7923),
            .in3(N__7971),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__9756));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_10_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_10_0  (
            .in0(N__10396),
            .in1(_gnd_net_),
            .in2(N__7961),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9963),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_11_10_1 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_11_10_1  (
            .in0(N__8883),
            .in1(N__8836),
            .in2(_gnd_net_),
            .in3(N__10097),
            .lcout(\U712_REG_SM.N_373 ),
            .ltout(\U712_REG_SM.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_10_2 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__8132),
            .in2(N__7974),
            .in3(N__8912),
            .lcout(\U712_REG_SM.N_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__10395),
            .in2(_gnd_net_),
            .in3(N__7941),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9963),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_10_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_10_4  (
            .in0(N__10394),
            .in1(N__8573),
            .in2(_gnd_net_),
            .in3(N__8649),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9963),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__7954),
            .in2(_gnd_net_),
            .in3(N__7940),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_10_7 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_11_10_7  (
            .in0(N__8913),
            .in1(N__8837),
            .in2(_gnd_net_),
            .in3(N__10098),
            .lcout(\U712_REG_SM.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8153),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9969),
            .ce(),
            .sr(N__9751));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_11_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_11_11_3  (
            .in0(N__11234),
            .in1(N__8133),
            .in2(_gnd_net_),
            .in3(N__8088),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9969),
            .ce(),
            .sr(N__9751));
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_11_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8121),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9969),
            .ce(),
            .sr(N__9751));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_11_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__8949),
            .in2(_gnd_net_),
            .in3(N__8777),
            .lcout(\U712_REG_SM.N_328 ),
            .ltout(\U712_REG_SM.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_12_1  (
            .in0(N__8108),
            .in1(N__8914),
            .in2(N__8115),
            .in3(N__8882),
            .lcout(\U712_REG_SM.N_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__8844),
            .in2(_gnd_net_),
            .in3(N__10101),
            .lcout(),
            .ltout(\U712_REG_SM.N_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_12_7 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_11_12_7  (
            .in0(N__8778),
            .in1(N__10400),
            .in2(N__8112),
            .in3(N__8087),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9975),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_11_13_0 .LUT_INIT=16'b0100000001100010;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_11_13_0  (
            .in0(N__8846),
            .in1(N__8393),
            .in2(N__8786),
            .in3(N__8107),
            .lcout(\U712_REG_SM.REGENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_11_13_4  (
            .in0(N__8847),
            .in1(N__8106),
            .in2(N__10104),
            .in3(N__8414),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_7 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_13_7  (
            .in0(N__8928),
            .in1(N__8922),
            .in2(N__8067),
            .in3(N__8475),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9981),
            .ce(),
            .sr(N__9745));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_14_0  (
            .in0(N__8469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9985),
            .ce(),
            .sr(N__9744));
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8433),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9985),
            .ce(),
            .sr(N__9744));
    defparam \U712_REG_SM.REGENn_LC_11_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_11_15_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_11_15_3 .LUT_INIT=16'b1100011011000100;
    LogicCell40 \U712_REG_SM.REGENn_LC_11_15_3  (
            .in0(N__8427),
            .in1(N__8389),
            .in2(N__10113),
            .in3(N__8418),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9988),
            .ce(),
            .sr(N__9743));
    defparam \U712_CHIP_RAM.CASn_LC_12_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_12_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_12_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8366),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9936),
            .ce(),
            .sr(N__9773));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_5_0  (
            .in0(N__9544),
            .in1(N__10733),
            .in2(_gnd_net_),
            .in3(N__9350),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10499),
            .sr(N__9765));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_1  (
            .in0(N__9552),
            .in1(N__10729),
            .in2(_gnd_net_),
            .in3(N__9351),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9221),
            .ce(N__10497),
            .sr(N__9761));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_6_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_6_4  (
            .in0(N__9171),
            .in1(_gnd_net_),
            .in2(N__10742),
            .in3(N__10797),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9221),
            .ce(N__10497),
            .sr(N__9761));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_7_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_7_1  (
            .in0(N__9602),
            .in1(N__10721),
            .in2(_gnd_net_),
            .in3(N__9154),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10495),
            .sr(N__9758));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_7_4  (
            .in0(N__9551),
            .in1(N__10720),
            .in2(_gnd_net_),
            .in3(N__9601),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10495),
            .sr(N__9758));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_7_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_7_7  (
            .in0(N__9069),
            .in1(N__10722),
            .in2(_gnd_net_),
            .in3(N__9495),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10495),
            .sr(N__9758));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_0  (
            .in0(N__8685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8713),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_8_3 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_12_8_3  (
            .in0(N__8714),
            .in1(N__8686),
            .in2(_gnd_net_),
            .in3(N__8665),
            .lcout(\U712_CYCLE_TERM.N_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_8_5 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_8_5  (
            .in0(N__8715),
            .in1(N__8687),
            .in2(N__8670),
            .in3(N__8640),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_8_6 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_12_8_6  (
            .in0(N__8666),
            .in1(N__10318),
            .in2(N__8652),
            .in3(N__8568),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9942),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_12_9_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_12_9_7  (
            .in0(N__8619),
            .in1(N__10736),
            .in2(N__8594),
            .in3(N__9282),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__9753));
    defparam pll_RNI8MQ3_LC_12_10_2.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8569),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_11_0 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_12_11_0  (
            .in0(N__9003),
            .in1(N__10232),
            .in2(N__8853),
            .in3(N__10103),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9958),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_12_11_3 .LUT_INIT=16'b1111100011011000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_12_11_3  (
            .in0(N__10231),
            .in1(N__8961),
            .in2(N__11884),
            .in3(N__9012),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9958),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_12_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__8993),
            .in2(_gnd_net_),
            .in3(N__8843),
            .lcout(),
            .ltout(\U712_REG_SM.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_12_12_1 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_12_12_1  (
            .in0(N__10325),
            .in1(N__8934),
            .in2(N__9006),
            .in3(N__10102),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9965),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_12_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_12_4  (
            .in0(N__8911),
            .in1(N__8841),
            .in2(N__8955),
            .in3(N__8994),
            .lcout(\U712_REG_SM.N_413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_5  (
            .in0(N__10100),
            .in1(N__8995),
            .in2(N__8852),
            .in3(N__8953),
            .lcout(\U712_REG_SM.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_12_6 .LUT_INIT=16'b0101010101000101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_12_6  (
            .in0(N__8954),
            .in1(N__8842),
            .in2(N__8787),
            .in3(N__10099),
            .lcout(\U712_REG_SM.STATE_COUNTc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_12_13_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_12_13_0  (
            .in0(N__8881),
            .in1(N__10065),
            .in2(_gnd_net_),
            .in3(N__8848),
            .lcout(\U712_REG_SM.N_308 ),
            .ltout(\U712_REG_SM.N_308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_13_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_12_13_1  (
            .in0(N__8877),
            .in1(N__8921),
            .in2(N__8886),
            .in3(N__10326),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9971),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_13_7 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_12_13_7  (
            .in0(N__8876),
            .in1(N__8845),
            .in2(N__10096),
            .in3(N__8776),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_15_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10327),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_5_1  (
            .in0(N__9349),
            .in1(N__10735),
            .in2(_gnd_net_),
            .in3(N__9396),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10503),
            .sr(N__9779));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_6_6  (
            .in0(N__9170),
            .in1(N__10734),
            .in2(_gnd_net_),
            .in3(N__10796),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10500),
            .sr(N__9767));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_7_0  (
            .in0(N__10557),
            .in1(N__10715),
            .in2(_gnd_net_),
            .in3(N__10795),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9218),
            .ce(N__10498),
            .sr(N__9764));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_4  (
            .in0(N__10558),
            .in1(N__10716),
            .in2(_gnd_net_),
            .in3(N__9068),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9218),
            .ce(N__10498),
            .sr(N__9764));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_5  (
            .in0(N__9494),
            .in1(_gnd_net_),
            .in2(N__10737),
            .in3(N__9288),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9218),
            .ce(N__10498),
            .sr(N__9764));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_8_1  (
            .in0(N__9493),
            .in1(N__10702),
            .in2(_gnd_net_),
            .in3(N__9067),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9217),
            .ce(N__10496),
            .sr(N__9760));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_4  (
            .in0(N__10560),
            .in1(N__10701),
            .in2(_gnd_net_),
            .in3(N__9066),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10493),
            .sr(N__9757));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__10317),
            .in2(_gnd_net_),
            .in3(N__10179),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9964),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_13_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__9823),
            .in2(_gnd_net_),
            .in3(N__10127),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_5_2  (
            .in0(N__9589),
            .in1(N__10714),
            .in2(_gnd_net_),
            .in3(N__9543),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9220),
            .ce(N__10505),
            .sr(N__9787));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_7_4  (
            .in0(N__9287),
            .in1(N__10642),
            .in2(_gnd_net_),
            .in3(N__9483),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10501),
            .sr(N__9768));
    defparam \U712_REG_SM.ASn_ess_LC_14_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_14_13_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_14_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10116),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9986),
            .ce(N__9414),
            .sr(N__9749));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_5 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_14_14_5  (
            .in0(N__11467),
            .in1(N__11602),
            .in2(N__11400),
            .in3(N__11250),
            .lcout(\U712_REG_SM.N_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_2 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \U712_CHIP_RAM.N_336_i_LC_14_20_2  (
            .in0(N__11689),
            .in1(N__11466),
            .in2(N__11617),
            .in3(N__11343),
            .lcout(N_336_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_5_2  (
            .in0(N__9392),
            .in1(N__9339),
            .in2(_gnd_net_),
            .in3(N__10713),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9219),
            .ce(N__10506),
            .sr(N__9793));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_15_7_1  (
            .in0(N__10665),
            .in1(N__10445),
            .in2(_gnd_net_),
            .in3(N__9286),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9216),
            .ce(N__10504),
            .sr(N__9780));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_2  (
            .in0(N__10785),
            .in1(N__10712),
            .in2(_gnd_net_),
            .in3(N__10559),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10502),
            .sr(N__9769));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_15_9_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_15_9_6  (
            .in0(N__10350),
            .in1(N__10458),
            .in2(_gnd_net_),
            .in3(N__10446),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9970),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_15_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__10300),
            .in2(_gnd_net_),
            .in3(N__10185),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9976),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_LC_15_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_15_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_15_13_6 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \U712_REG_SM.LDSn_LC_15_13_6  (
            .in0(N__10114),
            .in1(N__9636),
            .in2(N__10137),
            .in3(N__10154),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9989),
            .ce(),
            .sr(N__9752));
    defparam \U712_REG_SM.UDSn_LC_15_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_15_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_15_13_7 .LUT_INIT=16'b1111001111100010;
    LogicCell40 \U712_REG_SM.UDSn_LC_15_13_7  (
            .in0(N__10143),
            .in1(N__10136),
            .in2(N__10010),
            .in3(N__10115),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9989),
            .ce(),
            .sr(N__9752));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_15_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_15_14_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_15_14_5  (
            .in0(N__11603),
            .in1(N__11515),
            .in2(N__11259),
            .in3(N__11397),
            .lcout(\U712_REG_SM.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_335_i_LC_15_20_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_335_i_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_335_i_LC_15_20_0 .LUT_INIT=16'b0000010101110000;
    LogicCell40 \U712_CHIP_RAM.N_335_i_LC_15_20_0  (
            .in0(N__11690),
            .in1(N__11607),
            .in2(N__11380),
            .in3(N__11498),
            .lcout(N_335_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_337_i_LC_15_20_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_337_i_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_337_i_LC_15_20_4 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_CHIP_RAM.N_337_i_LC_15_20_4  (
            .in0(N__11691),
            .in1(N__11608),
            .in2(N__11381),
            .in3(N__11499),
            .lcout(N_337_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_177_i_LC_17_11_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_177_i_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_177_i_LC_17_11_1 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_177_i_LC_17_11_1  (
            .in0(N__11804),
            .in1(N__11043),
            .in2(N__11820),
            .in3(N__10965),
            .lcout(N_177_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m40_i_o2_LC_17_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m40_i_o2_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m40_i_o2_LC_17_14_0 .LUT_INIT=16'b1111010101001111;
    LogicCell40 \U712_CHIP_RAM.m40_i_o2_LC_17_14_0  (
            .in0(N__11705),
            .in1(N__11612),
            .in2(N__11379),
            .in3(N__11517),
            .lcout(N_334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_175_i_LC_18_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_175_i_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_175_i_LC_18_11_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_175_i_LC_18_11_0  (
            .in0(N__11123),
            .in1(N__11808),
            .in2(N__11766),
            .in3(N__10966),
            .lcout(N_175_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m58_i_o2_LC_18_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m58_i_o2_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m58_i_o2_LC_18_14_5 .LUT_INIT=16'b1100110100110111;
    LogicCell40 \U712_CHIP_RAM.m58_i_o2_LC_18_14_5  (
            .in0(N__11616),
            .in1(N__11399),
            .in2(N__11706),
            .in3(N__11482),
            .lcout(N_336),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m34_i_o2_LC_18_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m34_i_o2_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m34_i_o2_LC_18_14_6 .LUT_INIT=16'b1010111001011101;
    LogicCell40 \U712_CHIP_RAM.m34_i_o2_LC_18_14_6  (
            .in0(N__11481),
            .in1(N__11701),
            .in2(N__11619),
            .in3(N__11398),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_18_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_18_14_7 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_18_14_7  (
            .in0(N__10973),
            .in1(N__11754),
            .in2(N__11730),
            .in3(N__11110),
            .lcout(N_200_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_334_i_LC_18_20_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_334_i_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_334_i_LC_18_20_1 .LUT_INIT=16'b0000101110100000;
    LogicCell40 \U712_CHIP_RAM.N_334_i_LC_18_20_1  (
            .in0(N__11692),
            .in1(N__11618),
            .in2(N__11516),
            .in3(N__11368),
            .lcout(N_334_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_2 .LUT_INIT=16'b0010000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_2  (
            .in0(N__11120),
            .in1(N__11257),
            .in2(N__11020),
            .in3(N__11175),
            .lcout(N_379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_167_i_LC_24_19_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_167_i_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_167_i_LC_24_19_6 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_BUFFERS.N_167_i_LC_24_19_6  (
            .in0(N__11121),
            .in1(N__11013),
            .in2(N__10977),
            .in3(N__11898),
            .lcout(N_167_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP
